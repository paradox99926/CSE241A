/*
###############################################################
#  Design:            dynamic_node_top
###############################################################
*/
module dynamic_node_top (
	clk, 
	reset_in, 
	dataIn_N_63_, 
	dataIn_N_62_, 
	dataIn_N_61_, 
	dataIn_N_60_, 
	dataIn_N_59_, 
	dataIn_N_58_, 
	dataIn_N_57_, 
	dataIn_N_56_, 
	dataIn_N_55_, 
	dataIn_N_54_, 
	dataIn_N_53_, 
	dataIn_N_52_, 
	dataIn_N_51_, 
	dataIn_N_50_, 
	dataIn_N_49_, 
	dataIn_N_48_, 
	dataIn_N_47_, 
	dataIn_N_46_, 
	dataIn_N_45_, 
	dataIn_N_44_, 
	dataIn_N_43_, 
	dataIn_N_42_, 
	dataIn_N_41_, 
	dataIn_N_40_, 
	dataIn_N_39_, 
	dataIn_N_38_, 
	dataIn_N_37_, 
	dataIn_N_36_, 
	dataIn_N_35_, 
	dataIn_N_34_, 
	dataIn_N_33_, 
	dataIn_N_32_, 
	dataIn_N_31_, 
	dataIn_N_30_, 
	dataIn_N_29_, 
	dataIn_N_28_, 
	dataIn_N_27_, 
	dataIn_N_26_, 
	dataIn_N_25_, 
	dataIn_N_24_, 
	dataIn_N_23_, 
	dataIn_N_22_, 
	dataIn_N_21_, 
	dataIn_N_20_, 
	dataIn_N_19_, 
	dataIn_N_18_, 
	dataIn_N_17_, 
	dataIn_N_16_, 
	dataIn_N_15_, 
	dataIn_N_14_, 
	dataIn_N_13_, 
	dataIn_N_12_, 
	dataIn_N_11_, 
	dataIn_N_10_, 
	dataIn_N_9_, 
	dataIn_N_8_, 
	dataIn_N_7_, 
	dataIn_N_6_, 
	dataIn_N_5_, 
	dataIn_N_4_, 
	dataIn_N_3_, 
	dataIn_N_2_, 
	dataIn_N_1_, 
	dataIn_N_0_, 
	dataIn_E_63_, 
	dataIn_E_62_, 
	dataIn_E_61_, 
	dataIn_E_60_, 
	dataIn_E_59_, 
	dataIn_E_58_, 
	dataIn_E_57_, 
	dataIn_E_56_, 
	dataIn_E_55_, 
	dataIn_E_54_, 
	dataIn_E_53_, 
	dataIn_E_52_, 
	dataIn_E_51_, 
	dataIn_E_50_, 
	dataIn_E_49_, 
	dataIn_E_48_, 
	dataIn_E_47_, 
	dataIn_E_46_, 
	dataIn_E_45_, 
	dataIn_E_44_, 
	dataIn_E_43_, 
	dataIn_E_42_, 
	dataIn_E_41_, 
	dataIn_E_40_, 
	dataIn_E_39_, 
	dataIn_E_38_, 
	dataIn_E_37_, 
	dataIn_E_36_, 
	dataIn_E_35_, 
	dataIn_E_34_, 
	dataIn_E_33_, 
	dataIn_E_32_, 
	dataIn_E_31_, 
	dataIn_E_30_, 
	dataIn_E_29_, 
	dataIn_E_28_, 
	dataIn_E_27_, 
	dataIn_E_26_, 
	dataIn_E_25_, 
	dataIn_E_24_, 
	dataIn_E_23_, 
	dataIn_E_22_, 
	dataIn_E_21_, 
	dataIn_E_20_, 
	dataIn_E_19_, 
	dataIn_E_18_, 
	dataIn_E_17_, 
	dataIn_E_16_, 
	dataIn_E_15_, 
	dataIn_E_14_, 
	dataIn_E_13_, 
	dataIn_E_12_, 
	dataIn_E_11_, 
	dataIn_E_10_, 
	dataIn_E_9_, 
	dataIn_E_8_, 
	dataIn_E_7_, 
	dataIn_E_6_, 
	dataIn_E_5_, 
	dataIn_E_4_, 
	dataIn_E_3_, 
	dataIn_E_2_, 
	dataIn_E_1_, 
	dataIn_E_0_, 
	dataIn_S_63_, 
	dataIn_S_62_, 
	dataIn_S_61_, 
	dataIn_S_60_, 
	dataIn_S_59_, 
	dataIn_S_58_, 
	dataIn_S_57_, 
	dataIn_S_56_, 
	dataIn_S_55_, 
	dataIn_S_54_, 
	dataIn_S_53_, 
	dataIn_S_52_, 
	dataIn_S_51_, 
	dataIn_S_50_, 
	dataIn_S_49_, 
	dataIn_S_48_, 
	dataIn_S_47_, 
	dataIn_S_46_, 
	dataIn_S_45_, 
	dataIn_S_44_, 
	dataIn_S_43_, 
	dataIn_S_42_, 
	dataIn_S_41_, 
	dataIn_S_40_, 
	dataIn_S_39_, 
	dataIn_S_38_, 
	dataIn_S_37_, 
	dataIn_S_36_, 
	dataIn_S_35_, 
	dataIn_S_34_, 
	dataIn_S_33_, 
	dataIn_S_32_, 
	dataIn_S_31_, 
	dataIn_S_30_, 
	dataIn_S_29_, 
	dataIn_S_28_, 
	dataIn_S_27_, 
	dataIn_S_26_, 
	dataIn_S_25_, 
	dataIn_S_24_, 
	dataIn_S_23_, 
	dataIn_S_22_, 
	dataIn_S_21_, 
	dataIn_S_20_, 
	dataIn_S_19_, 
	dataIn_S_18_, 
	dataIn_S_17_, 
	dataIn_S_16_, 
	dataIn_S_15_, 
	dataIn_S_14_, 
	dataIn_S_13_, 
	dataIn_S_12_, 
	dataIn_S_11_, 
	dataIn_S_10_, 
	dataIn_S_9_, 
	dataIn_S_8_, 
	dataIn_S_7_, 
	dataIn_S_6_, 
	dataIn_S_5_, 
	dataIn_S_4_, 
	dataIn_S_3_, 
	dataIn_S_2_, 
	dataIn_S_1_, 
	dataIn_S_0_, 
	dataIn_W_63_, 
	dataIn_W_62_, 
	dataIn_W_61_, 
	dataIn_W_60_, 
	dataIn_W_59_, 
	dataIn_W_58_, 
	dataIn_W_57_, 
	dataIn_W_56_, 
	dataIn_W_55_, 
	dataIn_W_54_, 
	dataIn_W_53_, 
	dataIn_W_52_, 
	dataIn_W_51_, 
	dataIn_W_50_, 
	dataIn_W_49_, 
	dataIn_W_48_, 
	dataIn_W_47_, 
	dataIn_W_46_, 
	dataIn_W_45_, 
	dataIn_W_44_, 
	dataIn_W_43_, 
	dataIn_W_42_, 
	dataIn_W_41_, 
	dataIn_W_40_, 
	dataIn_W_39_, 
	dataIn_W_38_, 
	dataIn_W_37_, 
	dataIn_W_36_, 
	dataIn_W_35_, 
	dataIn_W_34_, 
	dataIn_W_33_, 
	dataIn_W_32_, 
	dataIn_W_31_, 
	dataIn_W_30_, 
	dataIn_W_29_, 
	dataIn_W_28_, 
	dataIn_W_27_, 
	dataIn_W_26_, 
	dataIn_W_25_, 
	dataIn_W_24_, 
	dataIn_W_23_, 
	dataIn_W_22_, 
	dataIn_W_21_, 
	dataIn_W_20_, 
	dataIn_W_19_, 
	dataIn_W_18_, 
	dataIn_W_17_, 
	dataIn_W_16_, 
	dataIn_W_15_, 
	dataIn_W_14_, 
	dataIn_W_13_, 
	dataIn_W_12_, 
	dataIn_W_11_, 
	dataIn_W_10_, 
	dataIn_W_9_, 
	dataIn_W_8_, 
	dataIn_W_7_, 
	dataIn_W_6_, 
	dataIn_W_5_, 
	dataIn_W_4_, 
	dataIn_W_3_, 
	dataIn_W_2_, 
	dataIn_W_1_, 
	dataIn_W_0_, 
	dataIn_P_63_, 
	dataIn_P_62_, 
	dataIn_P_61_, 
	dataIn_P_60_, 
	dataIn_P_59_, 
	dataIn_P_58_, 
	dataIn_P_57_, 
	dataIn_P_56_, 
	dataIn_P_55_, 
	dataIn_P_54_, 
	dataIn_P_53_, 
	dataIn_P_52_, 
	dataIn_P_51_, 
	dataIn_P_50_, 
	dataIn_P_49_, 
	dataIn_P_48_, 
	dataIn_P_47_, 
	dataIn_P_46_, 
	dataIn_P_45_, 
	dataIn_P_44_, 
	dataIn_P_43_, 
	dataIn_P_42_, 
	dataIn_P_41_, 
	dataIn_P_40_, 
	dataIn_P_39_, 
	dataIn_P_38_, 
	dataIn_P_37_, 
	dataIn_P_36_, 
	dataIn_P_35_, 
	dataIn_P_34_, 
	dataIn_P_33_, 
	dataIn_P_32_, 
	dataIn_P_31_, 
	dataIn_P_30_, 
	dataIn_P_29_, 
	dataIn_P_28_, 
	dataIn_P_27_, 
	dataIn_P_26_, 
	dataIn_P_25_, 
	dataIn_P_24_, 
	dataIn_P_23_, 
	dataIn_P_22_, 
	dataIn_P_21_, 
	dataIn_P_20_, 
	dataIn_P_19_, 
	dataIn_P_18_, 
	dataIn_P_17_, 
	dataIn_P_16_, 
	dataIn_P_15_, 
	dataIn_P_14_, 
	dataIn_P_13_, 
	dataIn_P_12_, 
	dataIn_P_11_, 
	dataIn_P_10_, 
	dataIn_P_9_, 
	dataIn_P_8_, 
	dataIn_P_7_, 
	dataIn_P_6_, 
	dataIn_P_5_, 
	dataIn_P_4_, 
	dataIn_P_3_, 
	dataIn_P_2_, 
	dataIn_P_1_, 
	dataIn_P_0_, 
	validIn_N, 
	validIn_E, 
	validIn_S, 
	validIn_W, 
	validIn_P, 
	yummyIn_N, 
	yummyIn_E, 
	yummyIn_S, 
	yummyIn_W, 
	yummyIn_P, 
	myLocX_7_, 
	myLocX_6_, 
	myLocX_5_, 
	myLocX_4_, 
	myLocX_3_, 
	myLocX_2_, 
	myLocX_1_, 
	myLocX_0_, 
	myLocY_7_, 
	myLocY_6_, 
	myLocY_5_, 
	myLocY_4_, 
	myLocY_3_, 
	myLocY_2_, 
	myLocY_1_, 
	myLocY_0_, 
	myChipID_13_, 
	myChipID_12_, 
	myChipID_11_, 
	myChipID_10_, 
	myChipID_9_, 
	myChipID_8_, 
	myChipID_7_, 
	myChipID_6_, 
	myChipID_5_, 
	myChipID_4_, 
	myChipID_3_, 
	myChipID_2_, 
	myChipID_1_, 
	myChipID_0_, 
	store_meter_partner_address_X_4_, 
	store_meter_partner_address_X_3_, 
	store_meter_partner_address_X_2_, 
	store_meter_partner_address_X_1_, 
	store_meter_partner_address_X_0_, 
	store_meter_partner_address_Y_4_, 
	store_meter_partner_address_Y_3_, 
	store_meter_partner_address_Y_2_, 
	store_meter_partner_address_Y_1_, 
	store_meter_partner_address_Y_0_, 
	ec_cfg_14_, 
	ec_cfg_13_, 
	ec_cfg_12_, 
	ec_cfg_11_, 
	ec_cfg_10_, 
	ec_cfg_9_, 
	ec_cfg_8_, 
	ec_cfg_7_, 
	ec_cfg_6_, 
	ec_cfg_5_, 
	ec_cfg_4_, 
	ec_cfg_3_, 
	ec_cfg_2_, 
	ec_cfg_1_, 
	ec_cfg_0_, 
	dataOut_N_63_, 
	dataOut_N_62_, 
	dataOut_N_61_, 
	dataOut_N_60_, 
	dataOut_N_59_, 
	dataOut_N_58_, 
	dataOut_N_57_, 
	dataOut_N_56_, 
	dataOut_N_55_, 
	dataOut_N_54_, 
	dataOut_N_53_, 
	dataOut_N_52_, 
	dataOut_N_51_, 
	dataOut_N_50_, 
	dataOut_N_49_, 
	dataOut_N_48_, 
	dataOut_N_47_, 
	dataOut_N_46_, 
	dataOut_N_45_, 
	dataOut_N_44_, 
	dataOut_N_43_, 
	dataOut_N_42_, 
	dataOut_N_41_, 
	dataOut_N_40_, 
	dataOut_N_39_, 
	dataOut_N_38_, 
	dataOut_N_37_, 
	dataOut_N_36_, 
	dataOut_N_35_, 
	dataOut_N_34_, 
	dataOut_N_33_, 
	dataOut_N_32_, 
	dataOut_N_31_, 
	dataOut_N_30_, 
	dataOut_N_29_, 
	dataOut_N_28_, 
	dataOut_N_27_, 
	dataOut_N_26_, 
	dataOut_N_25_, 
	dataOut_N_24_, 
	dataOut_N_23_, 
	dataOut_N_22_, 
	dataOut_N_21_, 
	dataOut_N_20_, 
	dataOut_N_19_, 
	dataOut_N_18_, 
	dataOut_N_17_, 
	dataOut_N_16_, 
	dataOut_N_15_, 
	dataOut_N_14_, 
	dataOut_N_13_, 
	dataOut_N_12_, 
	dataOut_N_11_, 
	dataOut_N_10_, 
	dataOut_N_9_, 
	dataOut_N_8_, 
	dataOut_N_7_, 
	dataOut_N_6_, 
	dataOut_N_5_, 
	dataOut_N_4_, 
	dataOut_N_3_, 
	dataOut_N_2_, 
	dataOut_N_1_, 
	dataOut_N_0_, 
	dataOut_E_63_, 
	dataOut_E_62_, 
	dataOut_E_61_, 
	dataOut_E_60_, 
	dataOut_E_59_, 
	dataOut_E_58_, 
	dataOut_E_57_, 
	dataOut_E_56_, 
	dataOut_E_55_, 
	dataOut_E_54_, 
	dataOut_E_53_, 
	dataOut_E_52_, 
	dataOut_E_51_, 
	dataOut_E_50_, 
	dataOut_E_49_, 
	dataOut_E_48_, 
	dataOut_E_47_, 
	dataOut_E_46_, 
	dataOut_E_45_, 
	dataOut_E_44_, 
	dataOut_E_43_, 
	dataOut_E_42_, 
	dataOut_E_41_, 
	dataOut_E_40_, 
	dataOut_E_39_, 
	dataOut_E_38_, 
	dataOut_E_37_, 
	dataOut_E_36_, 
	dataOut_E_35_, 
	dataOut_E_34_, 
	dataOut_E_33_, 
	dataOut_E_32_, 
	dataOut_E_31_, 
	dataOut_E_30_, 
	dataOut_E_29_, 
	dataOut_E_28_, 
	dataOut_E_27_, 
	dataOut_E_26_, 
	dataOut_E_25_, 
	dataOut_E_24_, 
	dataOut_E_23_, 
	dataOut_E_22_, 
	dataOut_E_21_, 
	dataOut_E_20_, 
	dataOut_E_19_, 
	dataOut_E_18_, 
	dataOut_E_17_, 
	dataOut_E_16_, 
	dataOut_E_15_, 
	dataOut_E_14_, 
	dataOut_E_13_, 
	dataOut_E_12_, 
	dataOut_E_11_, 
	dataOut_E_10_, 
	dataOut_E_9_, 
	dataOut_E_8_, 
	dataOut_E_7_, 
	dataOut_E_6_, 
	dataOut_E_5_, 
	dataOut_E_4_, 
	dataOut_E_3_, 
	dataOut_E_2_, 
	dataOut_E_1_, 
	dataOut_E_0_, 
	dataOut_S_63_, 
	dataOut_S_62_, 
	dataOut_S_61_, 
	dataOut_S_60_, 
	dataOut_S_59_, 
	dataOut_S_58_, 
	dataOut_S_57_, 
	dataOut_S_56_, 
	dataOut_S_55_, 
	dataOut_S_54_, 
	dataOut_S_53_, 
	dataOut_S_52_, 
	dataOut_S_51_, 
	dataOut_S_50_, 
	dataOut_S_49_, 
	dataOut_S_48_, 
	dataOut_S_47_, 
	dataOut_S_46_, 
	dataOut_S_45_, 
	dataOut_S_44_, 
	dataOut_S_43_, 
	dataOut_S_42_, 
	dataOut_S_41_, 
	dataOut_S_40_, 
	dataOut_S_39_, 
	dataOut_S_38_, 
	dataOut_S_37_, 
	dataOut_S_36_, 
	dataOut_S_35_, 
	dataOut_S_34_, 
	dataOut_S_33_, 
	dataOut_S_32_, 
	dataOut_S_31_, 
	dataOut_S_30_, 
	dataOut_S_29_, 
	dataOut_S_28_, 
	dataOut_S_27_, 
	dataOut_S_26_, 
	dataOut_S_25_, 
	dataOut_S_24_, 
	dataOut_S_23_, 
	dataOut_S_22_, 
	dataOut_S_21_, 
	dataOut_S_20_, 
	dataOut_S_19_, 
	dataOut_S_18_, 
	dataOut_S_17_, 
	dataOut_S_16_, 
	dataOut_S_15_, 
	dataOut_S_14_, 
	dataOut_S_13_, 
	dataOut_S_12_, 
	dataOut_S_11_, 
	dataOut_S_10_, 
	dataOut_S_9_, 
	dataOut_S_8_, 
	dataOut_S_7_, 
	dataOut_S_6_, 
	dataOut_S_5_, 
	dataOut_S_4_, 
	dataOut_S_3_, 
	dataOut_S_2_, 
	dataOut_S_1_, 
	dataOut_S_0_, 
	dataOut_W_63_, 
	dataOut_W_62_, 
	dataOut_W_61_, 
	dataOut_W_60_, 
	dataOut_W_59_, 
	dataOut_W_58_, 
	dataOut_W_57_, 
	dataOut_W_56_, 
	dataOut_W_55_, 
	dataOut_W_54_, 
	dataOut_W_53_, 
	dataOut_W_52_, 
	dataOut_W_51_, 
	dataOut_W_50_, 
	dataOut_W_49_, 
	dataOut_W_48_, 
	dataOut_W_47_, 
	dataOut_W_46_, 
	dataOut_W_45_, 
	dataOut_W_44_, 
	dataOut_W_43_, 
	dataOut_W_42_, 
	dataOut_W_41_, 
	dataOut_W_40_, 
	dataOut_W_39_, 
	dataOut_W_38_, 
	dataOut_W_37_, 
	dataOut_W_36_, 
	dataOut_W_35_, 
	dataOut_W_34_, 
	dataOut_W_33_, 
	dataOut_W_32_, 
	dataOut_W_31_, 
	dataOut_W_30_, 
	dataOut_W_29_, 
	dataOut_W_28_, 
	dataOut_W_27_, 
	dataOut_W_26_, 
	dataOut_W_25_, 
	dataOut_W_24_, 
	dataOut_W_23_, 
	dataOut_W_22_, 
	dataOut_W_21_, 
	dataOut_W_20_, 
	dataOut_W_19_, 
	dataOut_W_18_, 
	dataOut_W_17_, 
	dataOut_W_16_, 
	dataOut_W_15_, 
	dataOut_W_14_, 
	dataOut_W_13_, 
	dataOut_W_12_, 
	dataOut_W_11_, 
	dataOut_W_10_, 
	dataOut_W_9_, 
	dataOut_W_8_, 
	dataOut_W_7_, 
	dataOut_W_6_, 
	dataOut_W_5_, 
	dataOut_W_4_, 
	dataOut_W_3_, 
	dataOut_W_2_, 
	dataOut_W_1_, 
	dataOut_W_0_, 
	dataOut_P_63_, 
	dataOut_P_62_, 
	dataOut_P_61_, 
	dataOut_P_60_, 
	dataOut_P_59_, 
	dataOut_P_58_, 
	dataOut_P_57_, 
	dataOut_P_56_, 
	dataOut_P_55_, 
	dataOut_P_54_, 
	dataOut_P_53_, 
	dataOut_P_52_, 
	dataOut_P_51_, 
	dataOut_P_50_, 
	dataOut_P_49_, 
	dataOut_P_48_, 
	dataOut_P_47_, 
	dataOut_P_46_, 
	dataOut_P_45_, 
	dataOut_P_44_, 
	dataOut_P_43_, 
	dataOut_P_42_, 
	dataOut_P_41_, 
	dataOut_P_40_, 
	dataOut_P_39_, 
	dataOut_P_38_, 
	dataOut_P_37_, 
	dataOut_P_36_, 
	dataOut_P_35_, 
	dataOut_P_34_, 
	dataOut_P_33_, 
	dataOut_P_32_, 
	dataOut_P_31_, 
	dataOut_P_30_, 
	dataOut_P_29_, 
	dataOut_P_28_, 
	dataOut_P_27_, 
	dataOut_P_26_, 
	dataOut_P_25_, 
	dataOut_P_24_, 
	dataOut_P_23_, 
	dataOut_P_22_, 
	dataOut_P_21_, 
	dataOut_P_20_, 
	dataOut_P_19_, 
	dataOut_P_18_, 
	dataOut_P_17_, 
	dataOut_P_16_, 
	dataOut_P_15_, 
	dataOut_P_14_, 
	dataOut_P_13_, 
	dataOut_P_12_, 
	dataOut_P_11_, 
	dataOut_P_10_, 
	dataOut_P_9_, 
	dataOut_P_8_, 
	dataOut_P_7_, 
	dataOut_P_6_, 
	dataOut_P_5_, 
	dataOut_P_4_, 
	dataOut_P_3_, 
	dataOut_P_2_, 
	dataOut_P_1_, 
	dataOut_P_0_, 
	validOut_N, 
	validOut_E, 
	validOut_S, 
	validOut_W, 
	validOut_P, 
	yummyOut_N, 
	yummyOut_E, 
	yummyOut_S, 
	yummyOut_W, 
	yummyOut_P, 
	thanksIn_P, 
	external_interrupt, 
	store_meter_ack_partner, 
	store_meter_ack_non_partner, 
	ec_out_4_, 
	ec_out_3_, 
	ec_out_2_, 
	ec_out_1_, 
	ec_out_0_);
   input clk;
   input reset_in;
   input dataIn_N_63_;
   input dataIn_N_62_;
   input dataIn_N_61_;
   input dataIn_N_60_;
   input dataIn_N_59_;
   input dataIn_N_58_;
   input dataIn_N_57_;
   input dataIn_N_56_;
   input dataIn_N_55_;
   input dataIn_N_54_;
   input dataIn_N_53_;
   input dataIn_N_52_;
   input dataIn_N_51_;
   input dataIn_N_50_;
   input dataIn_N_49_;
   input dataIn_N_48_;
   input dataIn_N_47_;
   input dataIn_N_46_;
   input dataIn_N_45_;
   input dataIn_N_44_;
   input dataIn_N_43_;
   input dataIn_N_42_;
   input dataIn_N_41_;
   input dataIn_N_40_;
   input dataIn_N_39_;
   input dataIn_N_38_;
   input dataIn_N_37_;
   input dataIn_N_36_;
   input dataIn_N_35_;
   input dataIn_N_34_;
   input dataIn_N_33_;
   input dataIn_N_32_;
   input dataIn_N_31_;
   input dataIn_N_30_;
   input dataIn_N_29_;
   input dataIn_N_28_;
   input dataIn_N_27_;
   input dataIn_N_26_;
   input dataIn_N_25_;
   input dataIn_N_24_;
   input dataIn_N_23_;
   input dataIn_N_22_;
   input dataIn_N_21_;
   input dataIn_N_20_;
   input dataIn_N_19_;
   input dataIn_N_18_;
   input dataIn_N_17_;
   input dataIn_N_16_;
   input dataIn_N_15_;
   input dataIn_N_14_;
   input dataIn_N_13_;
   input dataIn_N_12_;
   input dataIn_N_11_;
   input dataIn_N_10_;
   input dataIn_N_9_;
   input dataIn_N_8_;
   input dataIn_N_7_;
   input dataIn_N_6_;
   input dataIn_N_5_;
   input dataIn_N_4_;
   input dataIn_N_3_;
   input dataIn_N_2_;
   input dataIn_N_1_;
   input dataIn_N_0_;
   input dataIn_E_63_;
   input dataIn_E_62_;
   input dataIn_E_61_;
   input dataIn_E_60_;
   input dataIn_E_59_;
   input dataIn_E_58_;
   input dataIn_E_57_;
   input dataIn_E_56_;
   input dataIn_E_55_;
   input dataIn_E_54_;
   input dataIn_E_53_;
   input dataIn_E_52_;
   input dataIn_E_51_;
   input dataIn_E_50_;
   input dataIn_E_49_;
   input dataIn_E_48_;
   input dataIn_E_47_;
   input dataIn_E_46_;
   input dataIn_E_45_;
   input dataIn_E_44_;
   input dataIn_E_43_;
   input dataIn_E_42_;
   input dataIn_E_41_;
   input dataIn_E_40_;
   input dataIn_E_39_;
   input dataIn_E_38_;
   input dataIn_E_37_;
   input dataIn_E_36_;
   input dataIn_E_35_;
   input dataIn_E_34_;
   input dataIn_E_33_;
   input dataIn_E_32_;
   input dataIn_E_31_;
   input dataIn_E_30_;
   input dataIn_E_29_;
   input dataIn_E_28_;
   input dataIn_E_27_;
   input dataIn_E_26_;
   input dataIn_E_25_;
   input dataIn_E_24_;
   input dataIn_E_23_;
   input dataIn_E_22_;
   input dataIn_E_21_;
   input dataIn_E_20_;
   input dataIn_E_19_;
   input dataIn_E_18_;
   input dataIn_E_17_;
   input dataIn_E_16_;
   input dataIn_E_15_;
   input dataIn_E_14_;
   input dataIn_E_13_;
   input dataIn_E_12_;
   input dataIn_E_11_;
   input dataIn_E_10_;
   input dataIn_E_9_;
   input dataIn_E_8_;
   input dataIn_E_7_;
   input dataIn_E_6_;
   input dataIn_E_5_;
   input dataIn_E_4_;
   input dataIn_E_3_;
   input dataIn_E_2_;
   input dataIn_E_1_;
   input dataIn_E_0_;
   input dataIn_S_63_;
   input dataIn_S_62_;
   input dataIn_S_61_;
   input dataIn_S_60_;
   input dataIn_S_59_;
   input dataIn_S_58_;
   input dataIn_S_57_;
   input dataIn_S_56_;
   input dataIn_S_55_;
   input dataIn_S_54_;
   input dataIn_S_53_;
   input dataIn_S_52_;
   input dataIn_S_51_;
   input dataIn_S_50_;
   input dataIn_S_49_;
   input dataIn_S_48_;
   input dataIn_S_47_;
   input dataIn_S_46_;
   input dataIn_S_45_;
   input dataIn_S_44_;
   input dataIn_S_43_;
   input dataIn_S_42_;
   input dataIn_S_41_;
   input dataIn_S_40_;
   input dataIn_S_39_;
   input dataIn_S_38_;
   input dataIn_S_37_;
   input dataIn_S_36_;
   input dataIn_S_35_;
   input dataIn_S_34_;
   input dataIn_S_33_;
   input dataIn_S_32_;
   input dataIn_S_31_;
   input dataIn_S_30_;
   input dataIn_S_29_;
   input dataIn_S_28_;
   input dataIn_S_27_;
   input dataIn_S_26_;
   input dataIn_S_25_;
   input dataIn_S_24_;
   input dataIn_S_23_;
   input dataIn_S_22_;
   input dataIn_S_21_;
   input dataIn_S_20_;
   input dataIn_S_19_;
   input dataIn_S_18_;
   input dataIn_S_17_;
   input dataIn_S_16_;
   input dataIn_S_15_;
   input dataIn_S_14_;
   input dataIn_S_13_;
   input dataIn_S_12_;
   input dataIn_S_11_;
   input dataIn_S_10_;
   input dataIn_S_9_;
   input dataIn_S_8_;
   input dataIn_S_7_;
   input dataIn_S_6_;
   input dataIn_S_5_;
   input dataIn_S_4_;
   input dataIn_S_3_;
   input dataIn_S_2_;
   input dataIn_S_1_;
   input dataIn_S_0_;
   input dataIn_W_63_;
   input dataIn_W_62_;
   input dataIn_W_61_;
   input dataIn_W_60_;
   input dataIn_W_59_;
   input dataIn_W_58_;
   input dataIn_W_57_;
   input dataIn_W_56_;
   input dataIn_W_55_;
   input dataIn_W_54_;
   input dataIn_W_53_;
   input dataIn_W_52_;
   input dataIn_W_51_;
   input dataIn_W_50_;
   input dataIn_W_49_;
   input dataIn_W_48_;
   input dataIn_W_47_;
   input dataIn_W_46_;
   input dataIn_W_45_;
   input dataIn_W_44_;
   input dataIn_W_43_;
   input dataIn_W_42_;
   input dataIn_W_41_;
   input dataIn_W_40_;
   input dataIn_W_39_;
   input dataIn_W_38_;
   input dataIn_W_37_;
   input dataIn_W_36_;
   input dataIn_W_35_;
   input dataIn_W_34_;
   input dataIn_W_33_;
   input dataIn_W_32_;
   input dataIn_W_31_;
   input dataIn_W_30_;
   input dataIn_W_29_;
   input dataIn_W_28_;
   input dataIn_W_27_;
   input dataIn_W_26_;
   input dataIn_W_25_;
   input dataIn_W_24_;
   input dataIn_W_23_;
   input dataIn_W_22_;
   input dataIn_W_21_;
   input dataIn_W_20_;
   input dataIn_W_19_;
   input dataIn_W_18_;
   input dataIn_W_17_;
   input dataIn_W_16_;
   input dataIn_W_15_;
   input dataIn_W_14_;
   input dataIn_W_13_;
   input dataIn_W_12_;
   input dataIn_W_11_;
   input dataIn_W_10_;
   input dataIn_W_9_;
   input dataIn_W_8_;
   input dataIn_W_7_;
   input dataIn_W_6_;
   input dataIn_W_5_;
   input dataIn_W_4_;
   input dataIn_W_3_;
   input dataIn_W_2_;
   input dataIn_W_1_;
   input dataIn_W_0_;
   input dataIn_P_63_;
   input dataIn_P_62_;
   input dataIn_P_61_;
   input dataIn_P_60_;
   input dataIn_P_59_;
   input dataIn_P_58_;
   input dataIn_P_57_;
   input dataIn_P_56_;
   input dataIn_P_55_;
   input dataIn_P_54_;
   input dataIn_P_53_;
   input dataIn_P_52_;
   input dataIn_P_51_;
   input dataIn_P_50_;
   input dataIn_P_49_;
   input dataIn_P_48_;
   input dataIn_P_47_;
   input dataIn_P_46_;
   input dataIn_P_45_;
   input dataIn_P_44_;
   input dataIn_P_43_;
   input dataIn_P_42_;
   input dataIn_P_41_;
   input dataIn_P_40_;
   input dataIn_P_39_;
   input dataIn_P_38_;
   input dataIn_P_37_;
   input dataIn_P_36_;
   input dataIn_P_35_;
   input dataIn_P_34_;
   input dataIn_P_33_;
   input dataIn_P_32_;
   input dataIn_P_31_;
   input dataIn_P_30_;
   input dataIn_P_29_;
   input dataIn_P_28_;
   input dataIn_P_27_;
   input dataIn_P_26_;
   input dataIn_P_25_;
   input dataIn_P_24_;
   input dataIn_P_23_;
   input dataIn_P_22_;
   input dataIn_P_21_;
   input dataIn_P_20_;
   input dataIn_P_19_;
   input dataIn_P_18_;
   input dataIn_P_17_;
   input dataIn_P_16_;
   input dataIn_P_15_;
   input dataIn_P_14_;
   input dataIn_P_13_;
   input dataIn_P_12_;
   input dataIn_P_11_;
   input dataIn_P_10_;
   input dataIn_P_9_;
   input dataIn_P_8_;
   input dataIn_P_7_;
   input dataIn_P_6_;
   input dataIn_P_5_;
   input dataIn_P_4_;
   input dataIn_P_3_;
   input dataIn_P_2_;
   input dataIn_P_1_;
   input dataIn_P_0_;
   input validIn_N;
   input validIn_E;
   input validIn_S;
   input validIn_W;
   input validIn_P;
   input yummyIn_N;
   input yummyIn_E;
   input yummyIn_S;
   input yummyIn_W;
   input yummyIn_P;
   input myLocX_7_;
   input myLocX_6_;
   input myLocX_5_;
   input myLocX_4_;
   input myLocX_3_;
   input myLocX_2_;
   input myLocX_1_;
   input myLocX_0_;
   input myLocY_7_;
   input myLocY_6_;
   input myLocY_5_;
   input myLocY_4_;
   input myLocY_3_;
   input myLocY_2_;
   input myLocY_1_;
   input myLocY_0_;
   input myChipID_13_;
   input myChipID_12_;
   input myChipID_11_;
   input myChipID_10_;
   input myChipID_9_;
   input myChipID_8_;
   input myChipID_7_;
   input myChipID_6_;
   input myChipID_5_;
   input myChipID_4_;
   input myChipID_3_;
   input myChipID_2_;
   input myChipID_1_;
   input myChipID_0_;
   input store_meter_partner_address_X_4_;
   input store_meter_partner_address_X_3_;
   input store_meter_partner_address_X_2_;
   input store_meter_partner_address_X_1_;
   input store_meter_partner_address_X_0_;
   input store_meter_partner_address_Y_4_;
   input store_meter_partner_address_Y_3_;
   input store_meter_partner_address_Y_2_;
   input store_meter_partner_address_Y_1_;
   input store_meter_partner_address_Y_0_;
   input ec_cfg_14_;
   input ec_cfg_13_;
   input ec_cfg_12_;
   input ec_cfg_11_;
   input ec_cfg_10_;
   input ec_cfg_9_;
   input ec_cfg_8_;
   input ec_cfg_7_;
   input ec_cfg_6_;
   input ec_cfg_5_;
   input ec_cfg_4_;
   input ec_cfg_3_;
   input ec_cfg_2_;
   input ec_cfg_1_;
   input ec_cfg_0_;
   output dataOut_N_63_;
   output dataOut_N_62_;
   output dataOut_N_61_;
   output dataOut_N_60_;
   output dataOut_N_59_;
   output dataOut_N_58_;
   output dataOut_N_57_;
   output dataOut_N_56_;
   output dataOut_N_55_;
   output dataOut_N_54_;
   output dataOut_N_53_;
   output dataOut_N_52_;
   output dataOut_N_51_;
   output dataOut_N_50_;
   output dataOut_N_49_;
   output dataOut_N_48_;
   output dataOut_N_47_;
   output dataOut_N_46_;
   output dataOut_N_45_;
   output dataOut_N_44_;
   output dataOut_N_43_;
   output dataOut_N_42_;
   output dataOut_N_41_;
   output dataOut_N_40_;
   output dataOut_N_39_;
   output dataOut_N_38_;
   output dataOut_N_37_;
   output dataOut_N_36_;
   output dataOut_N_35_;
   output dataOut_N_34_;
   output dataOut_N_33_;
   output dataOut_N_32_;
   output dataOut_N_31_;
   output dataOut_N_30_;
   output dataOut_N_29_;
   output dataOut_N_28_;
   output dataOut_N_27_;
   output dataOut_N_26_;
   output dataOut_N_25_;
   output dataOut_N_24_;
   output dataOut_N_23_;
   output dataOut_N_22_;
   output dataOut_N_21_;
   output dataOut_N_20_;
   output dataOut_N_19_;
   output dataOut_N_18_;
   output dataOut_N_17_;
   output dataOut_N_16_;
   output dataOut_N_15_;
   output dataOut_N_14_;
   output dataOut_N_13_;
   output dataOut_N_12_;
   output dataOut_N_11_;
   output dataOut_N_10_;
   output dataOut_N_9_;
   output dataOut_N_8_;
   output dataOut_N_7_;
   output dataOut_N_6_;
   output dataOut_N_5_;
   output dataOut_N_4_;
   output dataOut_N_3_;
   output dataOut_N_2_;
   output dataOut_N_1_;
   output dataOut_N_0_;
   output dataOut_E_63_;
   output dataOut_E_62_;
   output dataOut_E_61_;
   output dataOut_E_60_;
   output dataOut_E_59_;
   output dataOut_E_58_;
   output dataOut_E_57_;
   output dataOut_E_56_;
   output dataOut_E_55_;
   output dataOut_E_54_;
   output dataOut_E_53_;
   output dataOut_E_52_;
   output dataOut_E_51_;
   output dataOut_E_50_;
   output dataOut_E_49_;
   output dataOut_E_48_;
   output dataOut_E_47_;
   output dataOut_E_46_;
   output dataOut_E_45_;
   output dataOut_E_44_;
   output dataOut_E_43_;
   output dataOut_E_42_;
   output dataOut_E_41_;
   output dataOut_E_40_;
   output dataOut_E_39_;
   output dataOut_E_38_;
   output dataOut_E_37_;
   output dataOut_E_36_;
   output dataOut_E_35_;
   output dataOut_E_34_;
   output dataOut_E_33_;
   output dataOut_E_32_;
   output dataOut_E_31_;
   output dataOut_E_30_;
   output dataOut_E_29_;
   output dataOut_E_28_;
   output dataOut_E_27_;
   output dataOut_E_26_;
   output dataOut_E_25_;
   output dataOut_E_24_;
   output dataOut_E_23_;
   output dataOut_E_22_;
   output dataOut_E_21_;
   output dataOut_E_20_;
   output dataOut_E_19_;
   output dataOut_E_18_;
   output dataOut_E_17_;
   output dataOut_E_16_;
   output dataOut_E_15_;
   output dataOut_E_14_;
   output dataOut_E_13_;
   output dataOut_E_12_;
   output dataOut_E_11_;
   output dataOut_E_10_;
   output dataOut_E_9_;
   output dataOut_E_8_;
   output dataOut_E_7_;
   output dataOut_E_6_;
   output dataOut_E_5_;
   output dataOut_E_4_;
   output dataOut_E_3_;
   output dataOut_E_2_;
   output dataOut_E_1_;
   output dataOut_E_0_;
   output dataOut_S_63_;
   output dataOut_S_62_;
   output dataOut_S_61_;
   output dataOut_S_60_;
   output dataOut_S_59_;
   output dataOut_S_58_;
   output dataOut_S_57_;
   output dataOut_S_56_;
   output dataOut_S_55_;
   output dataOut_S_54_;
   output dataOut_S_53_;
   output dataOut_S_52_;
   output dataOut_S_51_;
   output dataOut_S_50_;
   output dataOut_S_49_;
   output dataOut_S_48_;
   output dataOut_S_47_;
   output dataOut_S_46_;
   output dataOut_S_45_;
   output dataOut_S_44_;
   output dataOut_S_43_;
   output dataOut_S_42_;
   output dataOut_S_41_;
   output dataOut_S_40_;
   output dataOut_S_39_;
   output dataOut_S_38_;
   output dataOut_S_37_;
   output dataOut_S_36_;
   output dataOut_S_35_;
   output dataOut_S_34_;
   output dataOut_S_33_;
   output dataOut_S_32_;
   output dataOut_S_31_;
   output dataOut_S_30_;
   output dataOut_S_29_;
   output dataOut_S_28_;
   output dataOut_S_27_;
   output dataOut_S_26_;
   output dataOut_S_25_;
   output dataOut_S_24_;
   output dataOut_S_23_;
   output dataOut_S_22_;
   output dataOut_S_21_;
   output dataOut_S_20_;
   output dataOut_S_19_;
   output dataOut_S_18_;
   output dataOut_S_17_;
   output dataOut_S_16_;
   output dataOut_S_15_;
   output dataOut_S_14_;
   output dataOut_S_13_;
   output dataOut_S_12_;
   output dataOut_S_11_;
   output dataOut_S_10_;
   output dataOut_S_9_;
   output dataOut_S_8_;
   output dataOut_S_7_;
   output dataOut_S_6_;
   output dataOut_S_5_;
   output dataOut_S_4_;
   output dataOut_S_3_;
   output dataOut_S_2_;
   output dataOut_S_1_;
   output dataOut_S_0_;
   output dataOut_W_63_;
   output dataOut_W_62_;
   output dataOut_W_61_;
   output dataOut_W_60_;
   output dataOut_W_59_;
   output dataOut_W_58_;
   output dataOut_W_57_;
   output dataOut_W_56_;
   output dataOut_W_55_;
   output dataOut_W_54_;
   output dataOut_W_53_;
   output dataOut_W_52_;
   output dataOut_W_51_;
   output dataOut_W_50_;
   output dataOut_W_49_;
   output dataOut_W_48_;
   output dataOut_W_47_;
   output dataOut_W_46_;
   output dataOut_W_45_;
   output dataOut_W_44_;
   output dataOut_W_43_;
   output dataOut_W_42_;
   output dataOut_W_41_;
   output dataOut_W_40_;
   output dataOut_W_39_;
   output dataOut_W_38_;
   output dataOut_W_37_;
   output dataOut_W_36_;
   output dataOut_W_35_;
   output dataOut_W_34_;
   output dataOut_W_33_;
   output dataOut_W_32_;
   output dataOut_W_31_;
   output dataOut_W_30_;
   output dataOut_W_29_;
   output dataOut_W_28_;
   output dataOut_W_27_;
   output dataOut_W_26_;
   output dataOut_W_25_;
   output dataOut_W_24_;
   output dataOut_W_23_;
   output dataOut_W_22_;
   output dataOut_W_21_;
   output dataOut_W_20_;
   output dataOut_W_19_;
   output dataOut_W_18_;
   output dataOut_W_17_;
   output dataOut_W_16_;
   output dataOut_W_15_;
   output dataOut_W_14_;
   output dataOut_W_13_;
   output dataOut_W_12_;
   output dataOut_W_11_;
   output dataOut_W_10_;
   output dataOut_W_9_;
   output dataOut_W_8_;
   output dataOut_W_7_;
   output dataOut_W_6_;
   output dataOut_W_5_;
   output dataOut_W_4_;
   output dataOut_W_3_;
   output dataOut_W_2_;
   output dataOut_W_1_;
   output dataOut_W_0_;
   output dataOut_P_63_;
   output dataOut_P_62_;
   output dataOut_P_61_;
   output dataOut_P_60_;
   output dataOut_P_59_;
   output dataOut_P_58_;
   output dataOut_P_57_;
   output dataOut_P_56_;
   output dataOut_P_55_;
   output dataOut_P_54_;
   output dataOut_P_53_;
   output dataOut_P_52_;
   output dataOut_P_51_;
   output dataOut_P_50_;
   output dataOut_P_49_;
   output dataOut_P_48_;
   output dataOut_P_47_;
   output dataOut_P_46_;
   output dataOut_P_45_;
   output dataOut_P_44_;
   output dataOut_P_43_;
   output dataOut_P_42_;
   output dataOut_P_41_;
   output dataOut_P_40_;
   output dataOut_P_39_;
   output dataOut_P_38_;
   output dataOut_P_37_;
   output dataOut_P_36_;
   output dataOut_P_35_;
   output dataOut_P_34_;
   output dataOut_P_33_;
   output dataOut_P_32_;
   output dataOut_P_31_;
   output dataOut_P_30_;
   output dataOut_P_29_;
   output dataOut_P_28_;
   output dataOut_P_27_;
   output dataOut_P_26_;
   output dataOut_P_25_;
   output dataOut_P_24_;
   output dataOut_P_23_;
   output dataOut_P_22_;
   output dataOut_P_21_;
   output dataOut_P_20_;
   output dataOut_P_19_;
   output dataOut_P_18_;
   output dataOut_P_17_;
   output dataOut_P_16_;
   output dataOut_P_15_;
   output dataOut_P_14_;
   output dataOut_P_13_;
   output dataOut_P_12_;
   output dataOut_P_11_;
   output dataOut_P_10_;
   output dataOut_P_9_;
   output dataOut_P_8_;
   output dataOut_P_7_;
   output dataOut_P_6_;
   output dataOut_P_5_;
   output dataOut_P_4_;
   output dataOut_P_3_;
   output dataOut_P_2_;
   output dataOut_P_1_;
   output dataOut_P_0_;
   output validOut_N;
   output validOut_E;
   output validOut_S;
   output validOut_W;
   output validOut_P;
   output yummyOut_N;
   output yummyOut_E;
   output yummyOut_S;
   output yummyOut_W;
   output yummyOut_P;
   output thanksIn_P;
   output external_interrupt;
   output store_meter_ack_partner;
   output store_meter_ack_non_partner;
   output ec_out_4_;
   output ec_out_3_;
   output ec_out_2_;
   output ec_out_1_;
   output ec_out_0_;

   // Internal wires
   wire FE_OFN25981_n21666;
   wire FE_OFN25980_n21666;
   wire FE_OFN25979_n21666;
   wire FE_OFN25978_n21666;
   wire FE_OFN25977_n21666;
   wire FE_OFN25976_n21666;
   wire FE_OFN25975_n21666;
   wire FE_OFN25974_n21666;
   wire FE_OFN25973_n21666;
   wire FE_OFN25972_n20135;
   wire FE_OFN25971_n20135;
   wire FE_RN_69;
   wire FE_OCPN25970_n24342;
   wire FE_RN_57_0;
   wire FE_RN_56_0;
   wire FE_RN_55_0;
   wire FE_RN_54_0;
   wire FE_RN_53_0;
   wire FE_RN_52_0;
   wire FE_RN_51_0;
   wire FE_RN_68;
   wire FE_RN_67;
   wire FE_RN_66;
   wire FE_RN_65;
   wire FE_RN_64;
   wire FE_RN_50_0;
   wire FE_RN_48_0;
   wire FE_RN_47_0;
   wire FE_RN_46_0;
   wire FE_RN_45_0;
   wire FE_RN_63;
   wire FE_RN_62;
   wire FE_RN_44_0;
   wire FE_RN_43_0;
   wire FE_RN_42_0;
   wire FE_RN_61;
   wire FE_RN_60;
   wire FE_RN_44;
   wire FE_RN_41_0;
   wire FE_RN_40_0;
   wire FE_RN_39_0;
   wire FE_OCPN25969_n19500;
   wire FE_OCPN25968_n19500;
   wire FE_OCPN25967_n19500;
   wire FE_RN_59;
   wire FE_OCPN25966_proc_input_NIB_head_ptr_f_2;
   wire FE_OCPN25965_proc_input_NIB_head_ptr_f_2;
   wire FE_RN_58;
   wire FE_RN_57;
   wire FE_RN_56;
   wire FE_RN_55;
   wire FE_RN_38_0;
   wire FE_RN_37_0;
   wire FE_RN_36_0;
   wire FE_RN_10;
   wire FE_OCPN25964_n18039;
   wire FE_OCPN25963_n18039;
   wire FE_OCPN25962_n18039;
   wire FE_OCPN25961_n18039;
   wire FE_OCPN25960_n18039;
   wire FE_OCPN25959_n18039;
   wire FE_OCPN25958_n18039;
   wire FE_OCPN25957_n18039;
   wire FE_OCPN25956_n18039;
   wire FE_OCPN25955_n18039;
   wire FE_OCPN25954_n18039;
   wire FE_OCPN25953_n18039;
   wire FE_OCPN25952_n18039;
   wire FE_OCPN25951_n18039;
   wire FE_OCPN25950_n18039;
   wire FE_OCPN25949_n18039;
   wire FE_RN_54;
   wire FE_RN_53;
   wire FE_RN_35_0;
   wire FE_RN_34_0;
   wire FE_RN_33_0;
   wire FE_OCPN25948_n19595;
   wire FE_OCPN25947_n19595;
   wire FE_RN_52;
   wire FE_RN_51;
   wire FE_RN_50;
   wire FE_RN_49;
   wire FE_RN_48;
   wire FE_RN_32_0;
   wire FE_RN_31_0;
   wire FE_RN_30_0;
   wire FE_RN_47;
   wire FE_RN_46;
   wire FE_RN_45;
   wire FE_RN_43;
   wire FE_RN_42;
   wire FE_RN_41;
   wire FE_RN_40;
   wire FE_RN_39;
   wire FE_RN_38;
   wire FE_RN_37;
   wire FE_RN_36;
   wire FE_RN_35;
   wire FE_RN_34;
   wire FE_OCPN25946_n19501;
   wire FE_RN_33;
   wire FE_RN_29_0;
   wire FE_RN_28_0;
   wire FE_RN_27_0;
   wire FE_RN_26_0;
   wire FE_RN_25_0;
   wire FE_RN_24_0;
   wire FE_RN_32;
   wire FE_OCPN25945_n24965;
   wire FE_OCPN25944_n24965;
   wire FE_OCPN25943_n24965;
   wire FE_OCPN25942_n24965;
   wire FE_OCPN25941_n24965;
   wire FE_OCPN25940_n24965;
   wire FE_OCPN25939_n24965;
   wire FE_OCPN25938_n24965;
   wire FE_OCPN25937_n24965;
   wire FE_OCPN25936_n24965;
   wire FE_OCPN25935_n24965;
   wire FE_RN_25;
   wire FE_RN_31;
   wire FE_RN_30;
   wire FE_OCPN25934_n24342;
   wire FE_OCPN25933_n24342;
   wire FE_OCPN25932_n19501;
   wire FE_OCPN25931_n19501;
   wire FE_OCPN25929_n18828;
   wire FE_OCPN25927_n18828;
   wire FE_OCPN25926_n18828;
   wire FE_OCPN25925_n18828;
   wire FE_RN_29;
   wire FE_RN_28;
   wire FE_RN_27;
   wire FE_RN_26;
   wire FE_RN_24;
   wire FE_RN_23;
   wire FE_RN_16;
   wire FE_OCPN25924_n19547;
   wire FE_OCPN25923_n19547;
   wire FE_OCPN25922_n19547;
   wire FE_OCPN25921_n19547;
   wire FE_OCPN25920_n19547;
   wire FE_OCPN25919_n19547;
   wire FE_OCPN25918_n19547;
   wire FE_OCPN25917_n19547;
   wire FE_OCPN25916_n19547;
   wire FE_OCPN25915_n19547;
   wire FE_OCPN25914_n19547;
   wire FE_OCPN25913_n19547;
   wire FE_OCPN25912_n19547;
   wire FE_OCPN25911_n19547;
   wire FE_OCPN25910_n19547;
   wire FE_OCPN25909_n19547;
   wire FE_OCPN25908_n19547;
   wire FE_RN_22;
   wire FE_RN_21;
   wire FE_RN_20;
   wire FE_RN_19;
   wire FE_RN_18;
   wire FE_RN_17;
   wire FE_RN_15;
   wire FE_RN_14;
   wire FE_RN_13;
   wire FE_RN_12;
   wire FE_RN_11;
   wire FE_RN_9;
   wire FE_RN_2;
   wire FE_OCPN25907_n19306;
   wire FE_OCPN25906_n19306;
   wire FE_OCPN25905_n19306;
   wire FE_RN_8;
   wire FE_RN_7;
   wire FE_RN_6;
   wire FE_RN_5;
   wire FE_RN_23_0;
   wire FE_RN_22_0;
   wire FE_RN_4;
   wire FE_OCPN25904_n18927;
   wire FE_RN_3;
   wire FE_RN_1;
   wire FE_RN_20_0;
   wire FE_RN_19_0;
   wire FE_RN_18_0;
   wire FE_OCPN25903_west_input_NIB_head_ptr_f_0;
   wire FE_OCPN25902_west_input_NIB_head_ptr_f_0;
   wire FE_OCPN25901_west_input_NIB_head_ptr_f_0;
   wire FE_OCPN25900_west_input_NIB_head_ptr_f_0;
   wire FE_OCPN25899_west_input_NIB_head_ptr_f_0;
   wire FE_OFN25895_n25395;
   wire FE_OFN25892_n25395;
   wire FE_OFN25891_n25395;
   wire FE_OFN25889_n25395;
   wire FE_OFN25888_n25395;
   wire FE_OFN25887_dataOut_S_48;
   wire FE_OFN25886_dataOut_S_48;
   wire FE_OFN25885_dataOut_N_48;
   wire FE_OFN25884_dataOut_N_48;
   wire FE_OFN25883_n19446;
   wire FE_OFN25882_n19446;
   wire FE_OFN25881_n19446;
   wire FE_OFN25880_n19446;
   wire FE_OFN25879_n19446;
   wire FE_OFN25878_n19446;
   wire FE_OFN25877_n19446;
   wire FE_OFN25876_n25842;
   wire FE_OFN25875_n25842;
   wire FE_OFN25874_n25842;
   wire FE_OFN25872_FE_OFN42_n19022;
   wire FE_OFN25871_FE_OFN42_n19022;
   wire FE_OFN25869_n21666;
   wire FE_OFN25868_n21666;
   wire FE_OFN25866_FE_OFN24766_n21069;
   wire FE_OFN25865_FE_OFN24766_n21069;
   wire FE_OFN25862_FE_OFN24766_n21069;
   wire FE_OFN25861_FE_OFN24766_n21069;
   wire FE_OFN25860_FE_OFN24766_n21069;
   wire FE_OFN25857_FE_OFN899_n17770;
   wire FE_OFN25855_FE_OFN899_n17770;
   wire FE_OFN25854_FE_OFN899_n17770;
   wire FE_OFN25853_FE_OFN899_n17770;
   wire FE_OFN25850_FE_OFN899_n17770;
   wire FE_OFN25849_FE_OFN899_n17770;
   wire FE_OFN25847_FE_OFN899_n17770;
   wire FE_OFN25846_FE_OFN899_n17770;
   wire FE_OFN25845_n20699;
   wire FE_OFN25843_n25972;
   wire FE_RN_17_0;
   wire FE_RN_16_0;
   wire FE_RN_15_0;
   wire FE_RN_14_0;
   wire FE_RN_13_0;
   wire FE_RN_12_0;
   wire FE_RN_11_0;
   wire FE_RN_10_0;
   wire FE_RN_9_0;
   wire FE_OCPN25841_n24342;
   wire FE_OCPN25840_n24342;
   wire FE_OCPN25839_n24342;
   wire FE_OCPN25838_n24342;
   wire FE_OCPN25837_n24342;
   wire FE_OCPN25836_n24342;
   wire FE_OCPN25835_n24342;
   wire FE_OCPN25834_n;
   wire FE_OCPN25832_n19500;
   wire FE_RN_8_0;
   wire FE_RN_6_0;
   wire FE_OCPN25831_n20535;
   wire FE_RN_5_0;
   wire FE_RN_4_0;
   wire FE_RN_3_0;
   wire FE_OCPN25830_n;
   wire FE_OCPN25829_n21745;
   wire FE_OCPN25828_n21745;
   wire FE_OCPN25827_n21745;
   wire FE_OCPN25826_n21745;
   wire FE_OCPN25825_n21745;
   wire FE_OCPN25824_n21745;
   wire FE_OCPN25823_n21745;
   wire FE_OCPN25822_n21745;
   wire FE_OCPN25821_n19632;
   wire FE_OCPN25820_west_input_NIB_head_ptr_f_1;
   wire FE_OCPN25819_n24342;
   wire FE_OCPN25816_n20147;
   wire FE_OCPN25814_FE_OFN186_n24453;
   wire FE_OCPN25813_FE_OFN24735_n19306;
   wire FE_OCPN25811_n18959;
   wire FE_OCPN25810_n18959;
   wire FE_OCPN25809_n18959;
   wire FE_OCPN25807_n18959;
   wire FE_RN_2_0;
   wire FE_RN_1_0;
   wire FE_RN_0_0;
   wire FE_OFN25806_n23051;
   wire FE_OFN25802_n23051;
   wire FE_OFN25801_n23051;
   wire FE_OFN25798_n23051;
   wire FE_OFN25797_n23051;
   wire FE_OFN25796_n23051;
   wire FE_OFN25795_n23051;
   wire FE_OFN25794_n21053;
   wire FE_OFN25792_n21053;
   wire FE_OFN25791_n21053;
   wire FE_OFN25790_n21053;
   wire FE_OFN25789_n21053;
   wire FE_OFN25788_n21053;
   wire FE_OFN25787_n17770;
   wire FE_OFN25785_n17770;
   wire FE_OFN25783_n17770;
   wire FE_OFN25782_FE_OFN448_n23236;
   wire FE_OFN25781_FE_OFN448_n23236;
   wire FE_OFN25780_FE_OFN448_n23236;
   wire FE_OFN25779_FE_OFN448_n23236;
   wire FE_OFN25778_FE_OFN582_n25619;
   wire FE_OFN25777_FE_OFN582_n25619;
   wire FE_OFN25776_FE_OFN582_n25619;
   wire FE_OFN25775_FE_OFN582_n25619;
   wire FE_OFN25774_FE_OFN582_n25619;
   wire FE_OFN25773_FE_OFN582_n25619;
   wire FE_OFN25772_FE_OFN582_n25619;
   wire FE_OFN25771_FE_OFN582_n25619;
   wire FE_OFN25770_FE_OFN582_n25619;
   wire FE_OFN25769_FE_OFN582_n25619;
   wire FE_OFN25768_FE_OFN1077_n17766;
   wire FE_OFN25767_FE_OFN1077_n17766;
   wire FE_OFN25766_FE_OFN1077_n17766;
   wire FE_OFN25765_FE_OFN1077_n17766;
   wire FE_OFN25763_FE_OFN1077_n17766;
   wire FE_OFN25762_FE_OFN1077_n17766;
   wire FE_OFN25761_FE_OFN1077_n17766;
   wire FE_OFN25760_FE_OFN1077_n17766;
   wire FE_OFN25759_FE_OFN1077_n17766;
   wire FE_OFN25758_FE_OFN1077_n17766;
   wire FE_OFN25757_FE_OFN1077_n17766;
   wire FE_OFN25756_FE_OFN1077_n17766;
   wire FE_OFN25755_FE_OFN1077_n17766;
   wire FE_OFN25754_FE_OFN1077_n17766;
   wire FE_OFN25753_FE_OFN24796_n20854;
   wire FE_OFN25751_FE_OFN24796_n20854;
   wire FE_OFN25750_FE_OFN24796_n20854;
   wire FE_OFN25749_FE_OFN24796_n20854;
   wire FE_OFN25748_FE_OFN24796_n20854;
   wire FE_OFN25747_FE_OFN24796_n20854;
   wire FE_OFN25745_FE_OFN24796_n20854;
   wire FE_OFN25744_FE_OFN24796_n20854;
   wire FE_OFN25743_FE_OFN24796_n20854;
   wire FE_OFN25742_FE_OFN25605_n21944;
   wire FE_OFN25741_FE_OFN25605_n21944;
   wire FE_OFN25740_FE_OFN25605_n21944;
   wire FE_OFN25739_FE_OFN25605_n21944;
   wire FE_OFN25738_FE_OFN25605_n21944;
   wire FE_OFN25737_FE_OFN25605_n21944;
   wire FE_OFN25736_FE_OFN25605_n21944;
   wire FE_OFN25735_FE_OFN25605_n21944;
   wire FE_OFN25734_dataOut_E_8;
   wire FE_OFN25733_dataOut_E_8;
   wire FE_OFN25732_dataOut_P_9;
   wire FE_OFN25731_dataOut_P_9;
   wire FE_OFN25730_dataOut_W_9;
   wire FE_OFN25729_dataOut_W_9;
   wire FE_OFN25728_dataOut_P_31;
   wire FE_OFN25727_dataOut_P_31;
   wire FE_OFN25726_dataOut_E_37;
   wire FE_OFN25725_dataOut_E_37;
   wire FE_OFN25724_dataOut_W_31;
   wire FE_OFN25723_dataOut_W_31;
   wire FE_OFN25722_dataOut_N_31;
   wire FE_OFN25721_dataOut_N_31;
   wire FE_OFN25720_dataOut_E_22;
   wire FE_OFN25719_dataOut_E_22;
   wire FE_OFN25718_dataOut_P_37;
   wire FE_OFN25717_dataOut_P_37;
   wire FE_OFN25716_dataOut_W_37;
   wire FE_OFN25715_dataOut_W_37;
   wire FE_OFN25714_dataOut_W_48;
   wire FE_OFN25713_dataOut_W_48;
   wire FE_OFN25712_dataOut_P_49;
   wire FE_OFN25711_dataOut_P_49;
   wire FE_OFN25710_dataOut_W_49;
   wire FE_OFN25709_dataOut_W_49;
   wire FE_OFN25708_dataOut_P_35;
   wire FE_OFN25707_dataOut_P_35;
   wire FE_OFN25706_dataOut_N_35;
   wire FE_OFN25705_dataOut_N_35;
   wire FE_OFN25704_dataOut_N_37;
   wire FE_OFN25703_dataOut_N_37;
   wire FE_OFN25702_dataOut_W_35;
   wire FE_OFN25701_dataOut_W_35;
   wire FE_OFN25700_dataOut_P_48;
   wire FE_OFN25699_dataOut_P_48;
   wire FE_OFN25698_dataOut_E_39;
   wire FE_OFN25697_dataOut_E_39;
   wire FE_OFN25696_n19372;
   wire FE_OFN25693_n19503;
   wire FE_OFN25692_n19503;
   wire FE_OFN25691_n19503;
   wire FE_OFN25690_n19503;
   wire FE_OFN25689_n19503;
   wire FE_OFN25688_n19500;
   wire FE_OFN25687_n19500;
   wire FE_OFN25686_n19500;
   wire FE_OFN25685_n19500;
   wire FE_OFN25684_n25474;
   wire FE_OFN25682_n17814;
   wire FE_OFN25681_n17814;
   wire FE_OFN25680_n17814;
   wire FE_OFN25679_n17814;
   wire FE_OFN25678_n17814;
   wire FE_OFN25677_n17814;
   wire FE_OFN25676_n20422;
   wire FE_OFN25675_n17777;
   wire FE_OFN25674_n18033;
   wire FE_OFN25673_n18033;
   wire FE_OFN25672_n22773;
   wire FE_OFN25671_n19655;
   wire FE_OFN25668_n18038;
   wire FE_OFN25667_n18959;
   wire FE_OFN25664_n19914;
   wire FE_OFN25663_n19914;
   wire FE_OFN25662_n19914;
   wire FE_OFN25661_n19914;
   wire FE_OFN25659_n19914;
   wire FE_OFN25652_n25499;
   wire FE_OFN25651_n25499;
   wire FE_OFN25648_n18762;
   wire FE_OFN25647_reset;
   wire FE_OFN25646_reset;
   wire FE_OFN25645_n21748;
   wire FE_OFN25644_n19504;
   wire FE_OFN25643_n19504;
   wire FE_OFN25642_n25062;
   wire FE_OFN25640_n19498;
   wire FE_OFN25638_n19230;
   wire FE_OFN25637_n19595;
   wire FE_OFN25636_n19595;
   wire FE_OFN25635_n19595;
   wire FE_OFN25634_n19595;
   wire FE_OFN25633_n19595;
   wire FE_OFN25632_n19595;
   wire FE_OFN25630_n19165;
   wire FE_OFN25629_n21910;
   wire FE_OFN25628_n21910;
   wire FE_OFN25627_n21910;
   wire FE_OFN25626_n21910;
   wire FE_OFN25624_n19003;
   wire FE_OFN25623_n19123;
   wire FE_OFN25622_n23789;
   wire FE_OFN25621_n23789;
   wire FE_OFN25620_n23789;
   wire FE_OFN25619_n23789;
   wire FE_OFN25618_n23789;
   wire FE_OFN25617_north_input_NIB_head_ptr_f_1;
   wire FE_OFN25616_n19007;
   wire FE_OFN25615_n19007;
   wire FE_OFN25614_n19237;
   wire FE_OFN25613_n17934;
   wire FE_OFN25610_n19071;
   wire FE_OFN25609_n18377;
   wire FE_OFN25607_n18151;
   wire FE_OFN25606_n19508;
   wire FE_OFN25605_n21944;
   wire FE_OFN25604_n19530;
   wire FE_OFN25602_n19530;
   wire FE_OFN25601_reset;
   wire FE_OFN25600_reset;
   wire FE_OFN25599_reset;
   wire FE_OFN25598_reset;
   wire FE_OFN25597_reset;
   wire FE_OFN25596_reset;
   wire FE_OFN24862_n22945;
   wire FE_OFN24861_n22945;
   wire FE_OFN24860_n22945;
   wire FE_OFN24859_n22945;
   wire FE_OFN24858_n22945;
   wire FE_OFN24857_n22945;
   wire FE_OFN24856_n22945;
   wire FE_OFN24855_n22945;
   wire FE_OFN24854_n22945;
   wire FE_OFN24853_n22945;
   wire FE_OFN24852_n22945;
   wire FE_OFN24851_n22945;
   wire FE_OFN24850_n22945;
   wire FE_OFN24849_n22945;
   wire FE_OFN24848_n22945;
   wire FE_OFN24847_n22945;
   wire FE_OFN24846_n22945;
   wire FE_OFN24845_n22945;
   wire FE_OFN24844_n22945;
   wire FE_OFN24843_n22945;
   wire FE_OFN24842_n22945;
   wire FE_OFN24841_n22945;
   wire FE_OFN24840_n22945;
   wire FE_OFN24839_n22945;
   wire FE_OFN24838_n22945;
   wire FE_OFN24837_n22945;
   wire FE_OFN24836_n22517;
   wire FE_OFN24835_n22517;
   wire FE_OFN24834_n22517;
   wire FE_OFN24833_n25232;
   wire FE_OFN24832_n25232;
   wire FE_OFN24831_n25232;
   wire FE_OFN24830_n25499;
   wire FE_OFN24829_n25499;
   wire FE_OFN24828_n25499;
   wire FE_OFN24827_n25499;
   wire FE_OFN24826_n25499;
   wire FE_OFN24825_n25499;
   wire FE_OFN24824_n24921;
   wire FE_OFN24823_n24921;
   wire FE_OFN24822_n24921;
   wire FE_OFN24821_n24921;
   wire FE_OFN24820_n24921;
   wire FE_OFN24819_n24921;
   wire FE_OFN24818_n24921;
   wire FE_OFN24817_n24921;
   wire FE_OFN24816_n24921;
   wire FE_OFN24815_n22958;
   wire FE_OFN24814_n22958;
   wire FE_OFN24813_n22958;
   wire FE_OFN24812_n22958;
   wire FE_OFN24811_n22958;
   wire FE_OFN24810_n22958;
   wire FE_OFN24809_n22958;
   wire FE_OFN24808_n22958;
   wire FE_OFN24807_n22958;
   wire FE_OFN24806_n19655;
   wire FE_OFN24803_n19500;
   wire FE_OFN24800_n20506;
   wire FE_OFN24799_n20506;
   wire FE_OFN24798_n19503;
   wire FE_OFN24796_n20854;
   wire FE_OFN24795_n20854;
   wire FE_OFN24794_n20854;
   wire FE_OFN24793_n17934;
   wire FE_OFN24792_n17934;
   wire FE_OFN24791_n24965;
   wire FE_OFN24788_n24965;
   wire FE_OFN24787_n19932;
   wire FE_OFN24780_n19932;
   wire FE_OFN24779_n19932;
   wire FE_OFN24778_n19932;
   wire FE_OFN24777_n19932;
   wire FE_OFN24776_n19073;
   wire FE_OFN24774_n19073;
   wire FE_OFN24773_n19075;
   wire FE_OFN24772_n19075;
   wire FE_OFN24771_n19075;
   wire FE_OFN24770_n19075;
   wire FE_OFN24769_n19075;
   wire FE_OFN24768_n19075;
   wire FE_OFN24767_n21069;
   wire FE_OFN24766_n21069;
   wire FE_OFN24764_n18960;
   wire FE_OFN24763_n18960;
   wire FE_OFN24762_n18960;
   wire FE_OFN24761_west_input_NIB_head_ptr_f_0;
   wire FE_OFN24748_n18828;
   wire FE_OFN24745_n18648;
   wire FE_OFN24744_n18648;
   wire FE_OFN24743_n19499;
   wire FE_OFN24742_n18683;
   wire FE_OFN24741_n18683;
   wire FE_OFN24737_n19306;
   wire FE_OFN24736_n19306;
   wire FE_OFN24735_n19306;
   wire FE_OFN24733_n19306;
   wire FE_OFN24732_n19306;
   wire FE_OFN24731_n18131;
   wire FE_OFN24730_n;
   wire FE_OFN24729_n;
   wire FE_OFN1102_n25965;
   wire FE_OFN1101_n25965;
   wire FE_OFN1100_n25937;
   wire FE_OFN1099_n25937;
   wire FE_OFN1098_n25937;
   wire FE_OFN1092_n20934;
   wire FE_OFN1090_n20855;
   wire FE_OFN1089_n20855;
   wire FE_OFN1087_n20656;
   wire FE_OFN1086_n22923;
   wire FE_OFN1085_n22923;
   wire FE_OFN1084_n20854;
   wire FE_OFN1083_n20854;
   wire FE_OFN1081_n17767;
   wire FE_OFN1080_n17767;
   wire FE_OFN1077_n17766;
   wire FE_OFN1076_n17766;
   wire FE_OFN1075_n17766;
   wire FE_OFN1074_n17766;
   wire FE_OFN1073_dataOut_P_2;
   wire FE_OFN1072_dataOut_P_2;
   wire FE_OFN1071_dataOut_P_3;
   wire FE_OFN1070_dataOut_P_3;
   wire FE_OFN1069_dataOut_P_4;
   wire FE_OFN1068_dataOut_P_4;
   wire FE_OFN1067_dataOut_P_5;
   wire FE_OFN1066_dataOut_P_5;
   wire FE_OFN1065_dataOut_P_7;
   wire FE_OFN1064_dataOut_P_7;
   wire FE_OFN1063_dataOut_P_8;
   wire FE_OFN1062_dataOut_P_8;
   wire FE_OFN1059_dataOut_P_12;
   wire FE_OFN1058_dataOut_P_12;
   wire FE_OFN1057_dataOut_P_14;
   wire FE_OFN1056_dataOut_P_14;
   wire FE_OFN1055_dataOut_P_18;
   wire FE_OFN1054_dataOut_P_18;
   wire FE_OFN1051_dataOut_W_2;
   wire FE_OFN1050_dataOut_W_2;
   wire FE_OFN1049_dataOut_W_3;
   wire FE_OFN1048_dataOut_W_3;
   wire FE_OFN1047_dataOut_W_4;
   wire FE_OFN1046_dataOut_W_4;
   wire FE_OFN1045_dataOut_W_5;
   wire FE_OFN1044_dataOut_W_5;
   wire FE_OFN1043_dataOut_W_7;
   wire FE_OFN1042_dataOut_W_7;
   wire FE_OFN1041_dataOut_W_8;
   wire FE_OFN1040_dataOut_W_8;
   wire FE_OFN1037_dataOut_W_12;
   wire FE_OFN1036_dataOut_W_12;
   wire FE_OFN1035_dataOut_W_14;
   wire FE_OFN1034_dataOut_W_14;
   wire FE_OFN1033_dataOut_W_18;
   wire FE_OFN1032_dataOut_W_18;
   wire FE_OFN1027_dataOut_S_2;
   wire FE_OFN1026_dataOut_S_2;
   wire FE_OFN1025_dataOut_S_3;
   wire FE_OFN1024_dataOut_S_3;
   wire FE_OFN1023_dataOut_S_4;
   wire FE_OFN1022_dataOut_S_4;
   wire FE_OFN1021_dataOut_S_5;
   wire FE_OFN1020_dataOut_S_5;
   wire FE_OFN1019_dataOut_S_7;
   wire FE_OFN1018_dataOut_S_7;
   wire FE_OFN1017_dataOut_S_8;
   wire FE_OFN1016_dataOut_S_8;
   wire FE_OFN1015_dataOut_S_9;
   wire FE_OFN1014_dataOut_S_9;
   wire FE_OFN1013_dataOut_S_12;
   wire FE_OFN1012_dataOut_S_12;
   wire FE_OFN1011_dataOut_S_14;
   wire FE_OFN1010_dataOut_S_14;
   wire FE_OFN1009_dataOut_S_18;
   wire FE_OFN1008_dataOut_S_18;
   wire FE_OFN1007_dataOut_S_31;
   wire FE_OFN1006_dataOut_S_31;
   wire FE_OFN1005_dataOut_E_2;
   wire FE_OFN1004_dataOut_E_2;
   wire FE_OFN1003_dataOut_E_3;
   wire FE_OFN1002_dataOut_E_3;
   wire FE_OFN1001_dataOut_E_4;
   wire FE_OFN1000_dataOut_E_4;
   wire FE_OFN999_dataOut_E_5;
   wire FE_OFN998_dataOut_E_5;
   wire FE_OFN997_dataOut_E_7;
   wire FE_OFN996_dataOut_E_7;
   wire FE_OFN993_dataOut_E_9;
   wire FE_OFN992_dataOut_E_9;
   wire FE_OFN991_dataOut_E_12;
   wire FE_OFN990_dataOut_E_12;
   wire FE_OFN989_dataOut_E_14;
   wire FE_OFN988_dataOut_E_14;
   wire FE_OFN987_dataOut_E_18;
   wire FE_OFN986_dataOut_E_18;
   wire FE_OFN981_dataOut_N_2;
   wire FE_OFN980_dataOut_N_2;
   wire FE_OFN979_dataOut_N_3;
   wire FE_OFN978_dataOut_N_3;
   wire FE_OFN977_dataOut_N_4;
   wire FE_OFN976_dataOut_N_4;
   wire FE_OFN975_dataOut_N_5;
   wire FE_OFN974_dataOut_N_5;
   wire FE_OFN973_dataOut_N_7;
   wire FE_OFN972_dataOut_N_7;
   wire FE_OFN971_dataOut_N_8;
   wire FE_OFN970_dataOut_N_8;
   wire FE_OFN969_dataOut_N_9;
   wire FE_OFN968_dataOut_N_9;
   wire FE_OFN967_dataOut_N_12;
   wire FE_OFN966_dataOut_N_12;
   wire FE_OFN965_dataOut_N_14;
   wire FE_OFN964_dataOut_N_14;
   wire FE_OFN963_dataOut_N_18;
   wire FE_OFN962_dataOut_N_18;
   wire FE_OFN959_n25972;
   wire FE_OFN958_n25972;
   wire FE_OFN953_n25916;
   wire FE_OFN952_n25916;
   wire FE_OFN951_n25881;
   wire FE_OFN950_n25881;
   wire FE_OFN947_n25096;
   wire FE_OFN946_n25096;
   wire FE_OFN945_n24998;
   wire FE_OFN943_n24921;
   wire FE_OFN942_n24921;
   wire FE_OFN941_n24921;
   wire FE_OFN940_n24921;
   wire FE_OFN937_n24710;
   wire FE_OFN934_n24710;
   wire FE_OFN923_n23576;
   wire FE_OFN922_n23576;
   wire FE_OFN914_n23246;
   wire FE_OFN913_n23246;
   wire FE_OFN912_n23246;
   wire FE_OFN907_n23046;
   wire FE_OFN906_n21586;
   wire FE_OFN905_n21586;
   wire FE_OFN904_n20750;
   wire FE_OFN903_n20750;
   wire FE_OFN902_n18421;
   wire FE_OFN899_n17770;
   wire FE_OFN896_n17769;
   wire FE_OFN884_dataOut_P_0;
   wire FE_OFN883_dataOut_P_0;
   wire FE_OFN882_dataOut_P_1;
   wire FE_OFN881_dataOut_P_1;
   wire FE_OFN880_dataOut_P_6;
   wire FE_OFN879_dataOut_P_6;
   wire FE_OFN878_dataOut_P_10;
   wire FE_OFN877_dataOut_P_10;
   wire FE_OFN876_dataOut_P_11;
   wire FE_OFN875_dataOut_P_11;
   wire FE_OFN874_dataOut_P_13;
   wire FE_OFN873_dataOut_P_13;
   wire FE_OFN872_dataOut_P_15;
   wire FE_OFN871_dataOut_P_15;
   wire FE_OFN870_dataOut_P_16;
   wire FE_OFN869_dataOut_P_16;
   wire FE_OFN868_dataOut_P_17;
   wire FE_OFN867_dataOut_P_17;
   wire FE_OFN866_dataOut_P_19;
   wire FE_OFN865_dataOut_P_19;
   wire FE_OFN864_dataOut_P_20;
   wire FE_OFN863_dataOut_P_20;
   wire FE_OFN862_dataOut_P_21;
   wire FE_OFN861_dataOut_P_21;
   wire FE_OFN858_dataOut_P_23;
   wire FE_OFN857_dataOut_P_23;
   wire FE_OFN856_dataOut_P_24;
   wire FE_OFN855_dataOut_P_24;
   wire FE_OFN854_dataOut_P_25;
   wire FE_OFN853_dataOut_P_25;
   wire FE_OFN848_dataOut_P_28;
   wire FE_OFN847_dataOut_P_28;
   wire FE_OFN846_dataOut_P_29;
   wire FE_OFN845_dataOut_P_29;
   wire FE_OFN844_dataOut_P_33;
   wire FE_OFN843_dataOut_P_33;
   wire FE_OFN842_dataOut_P_34;
   wire FE_OFN841_dataOut_P_34;
   wire FE_OFN838_dataOut_P_36;
   wire FE_OFN837_dataOut_P_36;
   wire FE_OFN834_dataOut_P_38;
   wire FE_OFN833_dataOut_P_38;
   wire FE_OFN832_dataOut_P_39;
   wire FE_OFN831_dataOut_P_39;
   wire FE_OFN830_dataOut_P_42;
   wire FE_OFN829_dataOut_P_42;
   wire FE_OFN828_dataOut_P_43;
   wire FE_OFN827_dataOut_P_43;
   wire FE_OFN810_dataOut_W_0;
   wire FE_OFN809_dataOut_W_0;
   wire FE_OFN808_dataOut_W_1;
   wire FE_OFN807_dataOut_W_1;
   wire FE_OFN806_dataOut_W_6;
   wire FE_OFN805_dataOut_W_6;
   wire FE_OFN804_dataOut_W_10;
   wire FE_OFN803_dataOut_W_10;
   wire FE_OFN802_dataOut_W_11;
   wire FE_OFN801_dataOut_W_11;
   wire FE_OFN800_dataOut_W_13;
   wire FE_OFN799_dataOut_W_13;
   wire FE_OFN798_dataOut_W_15;
   wire FE_OFN797_dataOut_W_15;
   wire FE_OFN796_dataOut_W_16;
   wire FE_OFN795_dataOut_W_16;
   wire FE_OFN794_dataOut_W_17;
   wire FE_OFN793_dataOut_W_17;
   wire FE_OFN792_dataOut_W_19;
   wire FE_OFN791_dataOut_W_19;
   wire FE_OFN790_dataOut_W_20;
   wire FE_OFN789_dataOut_W_20;
   wire FE_OFN788_dataOut_W_21;
   wire FE_OFN787_dataOut_W_21;
   wire FE_OFN784_dataOut_W_23;
   wire FE_OFN783_dataOut_W_23;
   wire FE_OFN782_dataOut_W_24;
   wire FE_OFN781_dataOut_W_24;
   wire FE_OFN780_dataOut_W_25;
   wire FE_OFN779_dataOut_W_25;
   wire FE_OFN776_dataOut_W_27;
   wire FE_OFN775_dataOut_W_27;
   wire FE_OFN774_dataOut_W_28;
   wire FE_OFN773_dataOut_W_28;
   wire FE_OFN770_dataOut_W_33;
   wire FE_OFN769_dataOut_W_33;
   wire FE_OFN768_dataOut_W_34;
   wire FE_OFN767_dataOut_W_34;
   wire FE_OFN764_dataOut_W_36;
   wire FE_OFN763_dataOut_W_36;
   wire FE_OFN760_dataOut_W_38;
   wire FE_OFN759_dataOut_W_38;
   wire FE_OFN758_dataOut_W_39;
   wire FE_OFN757_dataOut_W_39;
   wire FE_OFN756_dataOut_W_42;
   wire FE_OFN755_dataOut_W_42;
   wire FE_OFN748_dataOut_W_46;
   wire FE_OFN747_dataOut_W_46;
   wire FE_OFN734_dataOut_S_0;
   wire FE_OFN733_dataOut_S_0;
   wire FE_OFN732_dataOut_S_1;
   wire FE_OFN731_dataOut_S_1;
   wire FE_OFN730_dataOut_S_6;
   wire FE_OFN729_dataOut_S_6;
   wire FE_OFN728_dataOut_S_10;
   wire FE_OFN727_dataOut_S_10;
   wire FE_OFN726_dataOut_S_11;
   wire FE_OFN725_dataOut_S_11;
   wire FE_OFN724_dataOut_S_13;
   wire FE_OFN723_dataOut_S_13;
   wire FE_OFN722_dataOut_S_15;
   wire FE_OFN721_dataOut_S_15;
   wire FE_OFN720_dataOut_S_16;
   wire FE_OFN719_dataOut_S_16;
   wire FE_OFN718_dataOut_S_17;
   wire FE_OFN717_dataOut_S_17;
   wire FE_OFN716_dataOut_S_19;
   wire FE_OFN715_dataOut_S_19;
   wire FE_OFN714_dataOut_S_20;
   wire FE_OFN713_dataOut_S_20;
   wire FE_OFN712_dataOut_S_21;
   wire FE_OFN711_dataOut_S_21;
   wire FE_OFN710_dataOut_S_22;
   wire FE_OFN709_dataOut_S_22;
   wire FE_OFN708_dataOut_S_23;
   wire FE_OFN707_dataOut_S_23;
   wire FE_OFN706_dataOut_S_24;
   wire FE_OFN705_dataOut_S_24;
   wire FE_OFN704_dataOut_S_25;
   wire FE_OFN703_dataOut_S_25;
   wire FE_OFN702_dataOut_S_26;
   wire FE_OFN701_dataOut_S_26;
   wire FE_OFN700_dataOut_S_27;
   wire FE_OFN699_dataOut_S_27;
   wire FE_OFN698_dataOut_S_28;
   wire FE_OFN697_dataOut_S_28;
   wire FE_OFN696_dataOut_S_29;
   wire FE_OFN695_dataOut_S_29;
   wire FE_OFN694_dataOut_S_33;
   wire FE_OFN693_dataOut_S_33;
   wire FE_OFN692_dataOut_S_34;
   wire FE_OFN691_dataOut_S_34;
   wire FE_OFN690_dataOut_S_35;
   wire FE_OFN689_dataOut_S_35;
   wire FE_OFN688_dataOut_S_36;
   wire FE_OFN687_dataOut_S_36;
   wire FE_OFN686_dataOut_S_37;
   wire FE_OFN685_dataOut_S_37;
   wire FE_OFN684_dataOut_S_38;
   wire FE_OFN683_dataOut_S_38;
   wire FE_OFN682_dataOut_S_39;
   wire FE_OFN681_dataOut_S_39;
   wire FE_OFN680_dataOut_S_42;
   wire FE_OFN679_dataOut_S_42;
   wire FE_OFN678_dataOut_S_43;
   wire FE_OFN677_dataOut_S_43;
   wire FE_OFN666_dataOut_S_49;
   wire FE_OFN665_dataOut_S_49;
   wire FE_OFN660_dataOut_E_0;
   wire FE_OFN659_dataOut_E_0;
   wire FE_OFN656_dataOut_E_6;
   wire FE_OFN655_dataOut_E_6;
   wire FE_OFN654_dataOut_E_10;
   wire FE_OFN653_dataOut_E_10;
   wire FE_OFN652_dataOut_E_11;
   wire FE_OFN651_dataOut_E_11;
   wire FE_OFN650_dataOut_E_13;
   wire FE_OFN649_dataOut_E_13;
   wire FE_OFN648_dataOut_E_15;
   wire FE_OFN647_dataOut_E_15;
   wire FE_OFN644_dataOut_E_17;
   wire FE_OFN643_dataOut_E_17;
   wire FE_OFN642_dataOut_E_19;
   wire FE_OFN641_dataOut_E_19;
   wire FE_OFN640_dataOut_E_20;
   wire FE_OFN639_dataOut_E_20;
   wire FE_OFN638_dataOut_E_21;
   wire FE_OFN637_dataOut_E_21;
   wire FE_OFN634_dataOut_E_23;
   wire FE_OFN633_dataOut_E_23;
   wire FE_OFN632_dataOut_E_24;
   wire FE_OFN631_dataOut_E_24;
   wire FE_OFN628_dataOut_E_27;
   wire FE_OFN627_dataOut_E_27;
   wire FE_OFN626_dataOut_E_28;
   wire FE_OFN625_dataOut_E_28;
   wire FE_OFN624_dataOut_E_29;
   wire FE_OFN623_dataOut_E_29;
   wire FE_OFN622_dataOut_E_33;
   wire FE_OFN621_dataOut_E_33;
   wire FE_OFN620_dataOut_E_34;
   wire FE_OFN619_dataOut_E_34;
   wire FE_OFN616_dataOut_E_36;
   wire FE_OFN615_dataOut_E_36;
   wire FE_OFN612_dataOut_E_38;
   wire FE_OFN611_dataOut_E_38;
   wire FE_OFN608_dataOut_E_42;
   wire FE_OFN607_dataOut_E_42;
   wire FE_OFN596_dataOut_N_27;
   wire FE_OFN595_dataOut_N_27;
   wire FE_OFN585_n25643;
   wire FE_OFN584_n25643;
   wire FE_OFN582_n25619;
   wire FE_OFN580_n25547;
   wire FE_OFN579_n25511;
   wire FE_OFN578_n25511;
   wire FE_OFN577_n25498;
   wire FE_OFN576_n25498;
   wire FE_OFN575_n25463;
   wire FE_OFN574_n25463;
   wire FE_OFN573_n25463;
   wire FE_OFN572_n25463;
   wire FE_OFN571_n25463;
   wire FE_OFN570_n25395;
   wire FE_OFN569_n25395;
   wire FE_OFN567_n25395;
   wire FE_OFN566_n25395;
   wire FE_OFN565_n25385;
   wire FE_OFN563_n25120;
   wire FE_OFN559_n24969;
   wire FE_OFN558_n24969;
   wire FE_OFN557_n24969;
   wire FE_OFN556_n24761;
   wire FE_OFN555_n24761;
   wire FE_OFN554_n24761;
   wire FE_OFN553_n24761;
   wire FE_OFN546_n24751;
   wire FE_OFN545_n24751;
   wire FE_OFN540_n24743;
   wire FE_OFN539_n24743;
   wire FE_OFN538_n24743;
   wire FE_OFN537_n24743;
   wire FE_OFN536_n24743;
   wire FE_OFN535_n24743;
   wire FE_OFN534_n24743;
   wire FE_OFN533_n24743;
   wire FE_OFN530_n24733;
   wire FE_OFN529_n24733;
   wire FE_OFN528_n24732;
   wire FE_OFN527_n24732;
   wire FE_OFN526_n24731;
   wire FE_OFN525_n24731;
   wire FE_OFN524_n24728;
   wire FE_OFN523_n24728;
   wire FE_OFN522_n24728;
   wire FE_OFN521_n24723;
   wire FE_OFN520_n24723;
   wire FE_OFN517_n24712;
   wire FE_OFN516_n24712;
   wire FE_OFN515_n24702;
   wire FE_OFN514_n24702;
   wire FE_OFN513_n24695;
   wire FE_OFN512_n24695;
   wire FE_OFN499_n24601;
   wire FE_OFN498_n24601;
   wire FE_OFN497_n24586;
   wire FE_OFN496_n24586;
   wire FE_OFN495_n24579;
   wire FE_OFN494_n24579;
   wire FE_OFN493_n24577;
   wire FE_OFN492_n24577;
   wire FE_OFN491_n24022;
   wire FE_OFN490_n24022;
   wire FE_OFN487_n24013;
   wire FE_OFN486_n24013;
   wire FE_OFN485_n24011;
   wire FE_OFN484_n24011;
   wire FE_OFN483_n23987;
   wire FE_OFN482_n23987;
   wire FE_OFN479_n23631;
   wire FE_OFN478_n23631;
   wire FE_OFN477_n23578;
   wire FE_OFN476_n23578;
   wire FE_OFN473_n23560;
   wire FE_OFN472_n23560;
   wire FE_OFN465_n23476;
   wire FE_OFN453_n23262;
   wire FE_OFN452_n23262;
   wire FE_OFN448_n23236;
   wire FE_OFN442_n23051;
   wire FE_OFN440_n23051;
   wire FE_OFN438_n22958;
   wire FE_OFN437_n22958;
   wire FE_OFN436_n22958;
   wire FE_OFN435_n22958;
   wire FE_OFN434_n22958;
   wire FE_OFN433_n22945;
   wire FE_OFN432_n22945;
   wire FE_OFN431_n22945;
   wire FE_OFN430_n22945;
   wire FE_OFN428_n22902;
   wire FE_OFN427_n22778;
   wire FE_OFN426_n22778;
   wire FE_OFN425_n22778;
   wire FE_OFN424_n22766;
   wire FE_OFN423_n22766;
   wire FE_OFN418_n22535;
   wire FE_OFN417_n22535;
   wire FE_OFN416_n22085;
   wire FE_OFN412_n21671;
   wire FE_OFN411_n21671;
   wire FE_OFN408_n21421;
   wire FE_OFN407_n21421;
   wire FE_OFN403_n20815;
   wire FE_OFN396_n19493;
   wire FE_OFN395_n19493;
   wire FE_OFN394_n19446;
   wire FE_OFN393_n19446;
   wire FE_OFN391_n19446;
   wire FE_OFN390_n19446;
   wire FE_OFN389_n17786;
   wire FE_OFN388_n17786;
   wire FE_OFN387_n17783;
   wire FE_OFN386_n17783;
   wire FE_OFN382_n17772;
   wire FE_OFN381_n17772;
   wire FE_OFN380_n17772;
   wire FE_OFN374_n17762;
   wire FE_OFN373_n17762;
   wire FE_OFN370_n17761;
   wire FE_OFN369_n17761;
   wire FE_OFN368_n17761;
   wire FE_OFN366_n17753;
   wire FE_OFN365_dataOut_P_40;
   wire FE_OFN364_dataOut_P_40;
   wire FE_OFN363_dataOut_W_40;
   wire FE_OFN362_dataOut_W_40;
   wire FE_OFN361_dataOut_S_40;
   wire FE_OFN360_dataOut_S_40;
   wire FE_OFN355_dataOut_E_40;
   wire FE_OFN354_dataOut_E_40;
   wire FE_OFN353_dataOut_E_43;
   wire FE_OFN352_dataOut_E_43;
   wire FE_OFN343_dataOut_N_0;
   wire FE_OFN342_dataOut_N_0;
   wire FE_OFN341_dataOut_N_1;
   wire FE_OFN340_dataOut_N_1;
   wire FE_OFN339_dataOut_N_6;
   wire FE_OFN338_dataOut_N_6;
   wire FE_OFN337_dataOut_N_10;
   wire FE_OFN336_dataOut_N_10;
   wire FE_OFN335_dataOut_N_11;
   wire FE_OFN334_dataOut_N_11;
   wire FE_OFN333_dataOut_N_13;
   wire FE_OFN332_dataOut_N_13;
   wire FE_OFN331_dataOut_N_15;
   wire FE_OFN330_dataOut_N_15;
   wire FE_OFN329_dataOut_N_16;
   wire FE_OFN328_dataOut_N_16;
   wire FE_OFN327_dataOut_N_17;
   wire FE_OFN326_dataOut_N_17;
   wire FE_OFN325_dataOut_N_19;
   wire FE_OFN324_dataOut_N_19;
   wire FE_OFN323_dataOut_N_20;
   wire FE_OFN322_dataOut_N_20;
   wire FE_OFN321_dataOut_N_21;
   wire FE_OFN320_dataOut_N_21;
   wire FE_OFN317_dataOut_N_23;
   wire FE_OFN316_dataOut_N_23;
   wire FE_OFN315_dataOut_N_24;
   wire FE_OFN314_dataOut_N_24;
   wire FE_OFN313_dataOut_N_25;
   wire FE_OFN312_dataOut_N_25;
   wire FE_OFN311_dataOut_N_28;
   wire FE_OFN310_dataOut_N_28;
   wire FE_OFN309_dataOut_N_29;
   wire FE_OFN308_dataOut_N_29;
   wire FE_OFN305_dataOut_N_33;
   wire FE_OFN304_dataOut_N_33;
   wire FE_OFN303_dataOut_N_34;
   wire FE_OFN302_dataOut_N_34;
   wire FE_OFN299_dataOut_N_36;
   wire FE_OFN298_dataOut_N_36;
   wire FE_OFN295_dataOut_N_38;
   wire FE_OFN294_dataOut_N_38;
   wire FE_OFN293_dataOut_N_39;
   wire FE_OFN292_dataOut_N_39;
   wire FE_OFN291_dataOut_N_42;
   wire FE_OFN290_dataOut_N_42;
   wire FE_OFN289_dataOut_N_43;
   wire FE_OFN288_dataOut_N_43;
   wire FE_OFN272_n25595;
   wire FE_OFN269_n25506;
   wire FE_OFN268_n25506;
   wire FE_OFN266_n25499;
   wire FE_OFN265_n25427;
   wire FE_OFN264_n25427;
   wire FE_OFN262_n25301;
   wire FE_OFN261_n25301;
   wire FE_OFN260_n25295;
   wire FE_OFN259_n25295;
   wire FE_OFN258_n25295;
   wire FE_OFN257_n25294;
   wire FE_OFN256_n25294;
   wire FE_OFN255_n25247;
   wire FE_OFN254_n25247;
   wire FE_OFN253_n25241;
   wire FE_OFN252_n25241;
   wire FE_OFN251_n25152;
   wire FE_OFN250_n25152;
   wire FE_OFN249_n25152;
   wire FE_OFN248_n25152;
   wire FE_OFN247_n24982;
   wire FE_OFN246_n24982;
   wire FE_OFN242_n24744;
   wire FE_OFN241_n24744;
   wire FE_OFN239_n24739;
   wire FE_OFN238_n24739;
   wire FE_OFN237_n24730;
   wire FE_OFN236_n24730;
   wire FE_OFN235_n24729;
   wire FE_OFN234_n24729;
   wire FE_OFN233_n24719;
   wire FE_OFN232_n24719;
   wire FE_OFN231_n24704;
   wire FE_OFN230_n24704;
   wire FE_OFN229_n24684;
   wire FE_OFN228_n24684;
   wire FE_OFN227_n24677;
   wire FE_OFN226_n24677;
   wire FE_OFN223_n24664;
   wire FE_OFN222_n24664;
   wire FE_OFN221_n24662;
   wire FE_OFN220_n24662;
   wire FE_OFN219_n24645;
   wire FE_OFN218_n24645;
   wire FE_OFN217_n24637;
   wire FE_OFN216_n24637;
   wire FE_OFN215_n24636;
   wire FE_OFN214_n24636;
   wire FE_OFN211_n24630;
   wire FE_OFN210_n24630;
   wire FE_OFN207_n24619;
   wire FE_OFN206_n24619;
   wire FE_OFN203_n24600;
   wire FE_OFN202_n24600;
   wire FE_OFN201_n24584;
   wire FE_OFN200_n24584;
   wire FE_OFN191_n24454;
   wire FE_OFN188_n24453;
   wire FE_OFN186_n24453;
   wire FE_OFN183_n24390;
   wire FE_OFN178_n24364;
   wire FE_OFN177_n24364;
   wire FE_OFN176_n24364;
   wire FE_OFN170_n24343;
   wire FE_OFN169_n24343;
   wire FE_OFN168_n24343;
   wire FE_OFN167_n24343;
   wire FE_OFN165_n24129;
   wire FE_OFN161_n24129;
   wire FE_OFN156_n24129;
   wire FE_OFN155_n24036;
   wire FE_OFN154_n24036;
   wire FE_OFN153_n24027;
   wire FE_OFN152_n24027;
   wire FE_OFN151_n24019;
   wire FE_OFN150_n24019;
   wire FE_OFN146_n24010;
   wire FE_OFN145_n24010;
   wire FE_OFN144_n23991;
   wire FE_OFN143_n23991;
   wire FE_OFN142_n23964;
   wire FE_OFN141_n23964;
   wire FE_OFN140_n23959;
   wire FE_OFN139_n23959;
   wire FE_OFN138_n23948;
   wire FE_OFN137_n23948;
   wire FE_OFN136_n23623;
   wire FE_OFN135_n23623;
   wire FE_OFN134_n23594;
   wire FE_OFN133_n23594;
   wire FE_OFN130_n23559;
   wire FE_OFN129_n23559;
   wire FE_OFN128_n23536;
   wire FE_OFN127_n23536;
   wire FE_OFN122_n23520;
   wire FE_OFN120_n23482;
   wire FE_OFN119_n23482;
   wire FE_OFN116_n23148;
   wire FE_OFN115_n23148;
   wire FE_OFN114_n23102;
   wire FE_OFN113_n23102;
   wire FE_OFN112_n22773;
   wire FE_OFN111_n22773;
   wire FE_OFN110_n22771;
   wire FE_OFN109_n22771;
   wire FE_OFN108_n22518;
   wire FE_OFN107_n22518;
   wire FE_OFN106_n22517;
   wire FE_OFN105_n22517;
   wire FE_OFN104_n22140;
   wire FE_OFN103_n22140;
   wire FE_OFN101_n22098;
   wire FE_OFN100_n21907;
   wire FE_OFN99_n21907;
   wire FE_OFN97_n21865;
   wire FE_OFN96_n21865;
   wire FE_OFN94_n21695;
   wire FE_OFN93_n21667;
   wire FE_OFN92_n21667;
   wire FE_OFN91_n21590;
   wire FE_OFN90_n21590;
   wire FE_OFN88_n21220;
   wire FE_OFN86_n21175;
   wire FE_OFN84_n20972;
   wire FE_OFN83_n20814;
   wire FE_OFN82_n20814;
   wire FE_OFN79_n20501;
   wire FE_OFN78_n20501;
   wire FE_OFN73_n19631;
   wire FE_OFN67_n19548;
   wire FE_OFN65_n19542;
   wire FE_OFN63_n19518;
   wire FE_OFN62_n19518;
   wire FE_OFN61_n19435;
   wire FE_OFN60_n19435;
   wire FE_OFN59_n19435;
   wire FE_OFN58_n19435;
   wire FE_OFN53_n19355;
   wire FE_OFN51_n19193;
   wire FE_OFN48_n19193;
   wire FE_OFN47_n19056;
   wire FE_OFN46_n19056;
   wire FE_OFN45_n19054;
   wire FE_OFN44_n19054;
   wire FE_OFN43_n19054;
   wire FE_OFN42_n19022;
   wire FE_OFN41_n19022;
   wire FE_OFN35_n19017;
   wire FE_OFN34_n19017;
   wire FE_OFN30_n18974;
   wire FE_OFN28_n18974;
   wire FE_OFN27_n18974;
   wire FE_OFN26_n18974;
   wire FE_OFN25_n17787;
   wire FE_OFN24_n17787;
   wire FE_OFN20_n17779;
   wire FE_OFN15_south_input_NIB_head_ptr_f_1;
   wire FE_OFN8_reset;
   wire FE_OFN5_reset;
   wire FE_OFN4_reset;
   wire FE_OFN3_reset;
   wire FE_OFN2_reset;
   wire FE_OFN1_dataOut_N_40;
   wire FE_OFN0_dataOut_N_40;
   wire ec_thanks_n_to_n_reg;
   wire ec_thanks_n_to_e_reg;
   wire ec_thanks_n_to_s_reg;
   wire ec_thanks_n_to_w_reg;
   wire ec_thanks_n_to_p_reg;
   wire ec_thanks_e_to_n_reg;
   wire ec_thanks_e_to_e_reg;
   wire ec_thanks_e_to_s_reg;
   wire ec_thanks_e_to_w_reg;
   wire ec_thanks_e_to_p_reg;
   wire ec_thanks_s_to_n_reg;
   wire ec_thanks_s_to_e_reg;
   wire ec_thanks_s_to_s_reg;
   wire ec_thanks_s_to_w_reg;
   wire ec_thanks_s_to_p_reg;
   wire ec_thanks_w_to_n_reg;
   wire ec_thanks_w_to_e_reg;
   wire ec_thanks_w_to_s_reg;
   wire ec_thanks_w_to_w_reg;
   wire ec_thanks_w_to_p_reg;
   wire ec_thanks_p_to_n_reg;
   wire ec_thanks_p_to_e_reg;
   wire ec_thanks_p_to_s_reg;
   wire ec_thanks_p_to_w_reg;
   wire ec_thanks_p_to_p_reg;
   wire ec_north_input_valid_reg;
   wire north_input_valid;
   wire ec_east_input_valid_reg;
   wire east_input_valid;
   wire ec_south_input_valid_reg;
   wire south_input_valid;
   wire ec_west_input_valid_reg;
   wire west_input_valid;
   wire ec_proc_input_valid_reg;
   wire proc_input_valid;
   wire ec_wants_to_send_but_cannot_N;
   wire ec_wants_to_send_but_cannot_E;
   wire ec_wants_to_send_but_cannot_S;
   wire ec_wants_to_send_but_cannot_W;
   wire ec_wants_to_send_but_cannot_P;
   wire reset;
   wire myLocY_f_7_;
   wire myLocY_f_6_;
   wire myLocY_f_5_;
   wire myLocY_f_4_;
   wire myLocY_f_3_;
   wire myLocY_f_2_;
   wire myLocY_f_1_;
   wire myLocY_f_0_;
   wire myLocX_f_7_;
   wire myLocX_f_6_;
   wire myLocX_f_5_;
   wire myLocX_f_4_;
   wire myLocX_f_3_;
   wire myLocX_f_2_;
   wire myLocX_f_1_;
   wire myLocX_f_0_;
   wire myChipID_f_13_;
   wire myChipID_f_12_;
   wire myChipID_f_11_;
   wire myChipID_f_10_;
   wire myChipID_f_9_;
   wire myChipID_f_8_;
   wire myChipID_f_7_;
   wire myChipID_f_6_;
   wire myChipID_f_5_;
   wire myChipID_f_4_;
   wire myChipID_f_3_;
   wire myChipID_f_2_;
   wire myChipID_f_1_;
   wire myChipID_f_0_;
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N33;
   wire north_input_NIB_tail_ptr_f_0_;
   wire north_input_NIB_tail_ptr_f_1_;
   wire north_input_NIB_elements_in_array_f_0_;
   wire north_input_NIB_elements_in_array_f_1_;
   wire north_input_NIB_elements_in_array_f_2_;
   wire north_input_NIB_storage_data_f_3__0_;
   wire north_input_NIB_storage_data_f_3__1_;
   wire north_input_NIB_storage_data_f_3__2_;
   wire north_input_NIB_storage_data_f_3__3_;
   wire north_input_NIB_storage_data_f_3__4_;
   wire north_input_NIB_storage_data_f_3__5_;
   wire north_input_NIB_storage_data_f_3__6_;
   wire north_input_NIB_storage_data_f_3__7_;
   wire north_input_NIB_storage_data_f_3__8_;
   wire north_input_NIB_storage_data_f_3__9_;
   wire north_input_NIB_storage_data_f_3__10_;
   wire north_input_NIB_storage_data_f_3__11_;
   wire north_input_NIB_storage_data_f_3__12_;
   wire north_input_NIB_storage_data_f_3__13_;
   wire north_input_NIB_storage_data_f_3__14_;
   wire north_input_NIB_storage_data_f_3__15_;
   wire north_input_NIB_storage_data_f_3__16_;
   wire north_input_NIB_storage_data_f_3__17_;
   wire north_input_NIB_storage_data_f_3__18_;
   wire north_input_NIB_storage_data_f_3__19_;
   wire north_input_NIB_storage_data_f_3__20_;
   wire north_input_NIB_storage_data_f_3__21_;
   wire north_input_NIB_storage_data_f_3__22_;
   wire north_input_NIB_storage_data_f_3__23_;
   wire north_input_NIB_storage_data_f_3__24_;
   wire north_input_NIB_storage_data_f_3__25_;
   wire north_input_NIB_storage_data_f_3__26_;
   wire north_input_NIB_storage_data_f_3__27_;
   wire north_input_NIB_storage_data_f_3__28_;
   wire north_input_NIB_storage_data_f_3__29_;
   wire north_input_NIB_storage_data_f_3__30_;
   wire north_input_NIB_storage_data_f_3__31_;
   wire north_input_NIB_storage_data_f_3__32_;
   wire north_input_NIB_storage_data_f_3__33_;
   wire north_input_NIB_storage_data_f_3__34_;
   wire north_input_NIB_storage_data_f_3__35_;
   wire north_input_NIB_storage_data_f_3__36_;
   wire north_input_NIB_storage_data_f_3__37_;
   wire north_input_NIB_storage_data_f_3__38_;
   wire north_input_NIB_storage_data_f_3__39_;
   wire north_input_NIB_storage_data_f_3__40_;
   wire north_input_NIB_storage_data_f_3__41_;
   wire north_input_NIB_storage_data_f_3__42_;
   wire north_input_NIB_storage_data_f_3__43_;
   wire north_input_NIB_storage_data_f_3__44_;
   wire north_input_NIB_storage_data_f_3__45_;
   wire north_input_NIB_storage_data_f_3__46_;
   wire north_input_NIB_storage_data_f_3__47_;
   wire north_input_NIB_storage_data_f_3__48_;
   wire north_input_NIB_storage_data_f_3__49_;
   wire north_input_NIB_storage_data_f_3__50_;
   wire north_input_NIB_storage_data_f_3__51_;
   wire north_input_NIB_storage_data_f_3__52_;
   wire north_input_NIB_storage_data_f_3__53_;
   wire north_input_NIB_storage_data_f_3__54_;
   wire north_input_NIB_storage_data_f_3__55_;
   wire north_input_NIB_storage_data_f_3__56_;
   wire north_input_NIB_storage_data_f_3__57_;
   wire north_input_NIB_storage_data_f_3__58_;
   wire north_input_NIB_storage_data_f_3__59_;
   wire north_input_NIB_storage_data_f_3__60_;
   wire north_input_NIB_storage_data_f_3__61_;
   wire north_input_NIB_storage_data_f_3__62_;
   wire north_input_NIB_storage_data_f_3__63_;
   wire north_input_NIB_storage_data_f_2__0_;
   wire north_input_NIB_storage_data_f_2__1_;
   wire north_input_NIB_storage_data_f_2__2_;
   wire north_input_NIB_storage_data_f_2__3_;
   wire north_input_NIB_storage_data_f_2__4_;
   wire north_input_NIB_storage_data_f_2__5_;
   wire north_input_NIB_storage_data_f_2__6_;
   wire north_input_NIB_storage_data_f_2__7_;
   wire north_input_NIB_storage_data_f_2__8_;
   wire north_input_NIB_storage_data_f_2__9_;
   wire north_input_NIB_storage_data_f_2__10_;
   wire north_input_NIB_storage_data_f_2__11_;
   wire north_input_NIB_storage_data_f_2__12_;
   wire north_input_NIB_storage_data_f_2__13_;
   wire north_input_NIB_storage_data_f_2__14_;
   wire north_input_NIB_storage_data_f_2__15_;
   wire north_input_NIB_storage_data_f_2__16_;
   wire north_input_NIB_storage_data_f_2__17_;
   wire north_input_NIB_storage_data_f_2__18_;
   wire north_input_NIB_storage_data_f_2__19_;
   wire north_input_NIB_storage_data_f_2__20_;
   wire north_input_NIB_storage_data_f_2__21_;
   wire north_input_NIB_storage_data_f_2__22_;
   wire north_input_NIB_storage_data_f_2__23_;
   wire north_input_NIB_storage_data_f_2__24_;
   wire north_input_NIB_storage_data_f_2__25_;
   wire north_input_NIB_storage_data_f_2__26_;
   wire north_input_NIB_storage_data_f_2__27_;
   wire north_input_NIB_storage_data_f_2__28_;
   wire north_input_NIB_storage_data_f_2__29_;
   wire north_input_NIB_storage_data_f_2__30_;
   wire north_input_NIB_storage_data_f_2__31_;
   wire north_input_NIB_storage_data_f_2__32_;
   wire north_input_NIB_storage_data_f_2__33_;
   wire north_input_NIB_storage_data_f_2__34_;
   wire north_input_NIB_storage_data_f_2__35_;
   wire north_input_NIB_storage_data_f_2__36_;
   wire north_input_NIB_storage_data_f_2__37_;
   wire north_input_NIB_storage_data_f_2__38_;
   wire north_input_NIB_storage_data_f_2__39_;
   wire north_input_NIB_storage_data_f_2__40_;
   wire north_input_NIB_storage_data_f_2__41_;
   wire north_input_NIB_storage_data_f_2__42_;
   wire north_input_NIB_storage_data_f_2__43_;
   wire north_input_NIB_storage_data_f_2__44_;
   wire north_input_NIB_storage_data_f_2__45_;
   wire north_input_NIB_storage_data_f_2__46_;
   wire north_input_NIB_storage_data_f_2__47_;
   wire north_input_NIB_storage_data_f_2__48_;
   wire north_input_NIB_storage_data_f_2__49_;
   wire north_input_NIB_storage_data_f_2__50_;
   wire north_input_NIB_storage_data_f_2__51_;
   wire north_input_NIB_storage_data_f_2__52_;
   wire north_input_NIB_storage_data_f_2__53_;
   wire north_input_NIB_storage_data_f_2__54_;
   wire north_input_NIB_storage_data_f_2__55_;
   wire north_input_NIB_storage_data_f_2__56_;
   wire north_input_NIB_storage_data_f_2__57_;
   wire north_input_NIB_storage_data_f_2__58_;
   wire north_input_NIB_storage_data_f_2__59_;
   wire north_input_NIB_storage_data_f_2__60_;
   wire north_input_NIB_storage_data_f_2__61_;
   wire north_input_NIB_storage_data_f_2__62_;
   wire north_input_NIB_storage_data_f_2__63_;
   wire north_input_NIB_storage_data_f_1__0_;
   wire north_input_NIB_storage_data_f_1__1_;
   wire north_input_NIB_storage_data_f_1__2_;
   wire north_input_NIB_storage_data_f_1__3_;
   wire north_input_NIB_storage_data_f_1__4_;
   wire north_input_NIB_storage_data_f_1__5_;
   wire north_input_NIB_storage_data_f_1__6_;
   wire north_input_NIB_storage_data_f_1__7_;
   wire north_input_NIB_storage_data_f_1__8_;
   wire north_input_NIB_storage_data_f_1__9_;
   wire north_input_NIB_storage_data_f_1__10_;
   wire north_input_NIB_storage_data_f_1__11_;
   wire north_input_NIB_storage_data_f_1__12_;
   wire north_input_NIB_storage_data_f_1__13_;
   wire north_input_NIB_storage_data_f_1__14_;
   wire north_input_NIB_storage_data_f_1__15_;
   wire north_input_NIB_storage_data_f_1__16_;
   wire north_input_NIB_storage_data_f_1__17_;
   wire north_input_NIB_storage_data_f_1__18_;
   wire north_input_NIB_storage_data_f_1__19_;
   wire north_input_NIB_storage_data_f_1__20_;
   wire north_input_NIB_storage_data_f_1__21_;
   wire north_input_NIB_storage_data_f_1__22_;
   wire north_input_NIB_storage_data_f_1__23_;
   wire north_input_NIB_storage_data_f_1__24_;
   wire north_input_NIB_storage_data_f_1__25_;
   wire north_input_NIB_storage_data_f_1__26_;
   wire north_input_NIB_storage_data_f_1__27_;
   wire north_input_NIB_storage_data_f_1__28_;
   wire north_input_NIB_storage_data_f_1__29_;
   wire north_input_NIB_storage_data_f_1__30_;
   wire north_input_NIB_storage_data_f_1__31_;
   wire north_input_NIB_storage_data_f_1__32_;
   wire north_input_NIB_storage_data_f_1__33_;
   wire north_input_NIB_storage_data_f_1__34_;
   wire north_input_NIB_storage_data_f_1__35_;
   wire north_input_NIB_storage_data_f_1__36_;
   wire north_input_NIB_storage_data_f_1__37_;
   wire north_input_NIB_storage_data_f_1__38_;
   wire north_input_NIB_storage_data_f_1__39_;
   wire north_input_NIB_storage_data_f_1__40_;
   wire north_input_NIB_storage_data_f_1__41_;
   wire north_input_NIB_storage_data_f_1__42_;
   wire north_input_NIB_storage_data_f_1__43_;
   wire north_input_NIB_storage_data_f_1__44_;
   wire north_input_NIB_storage_data_f_1__45_;
   wire north_input_NIB_storage_data_f_1__46_;
   wire north_input_NIB_storage_data_f_1__47_;
   wire north_input_NIB_storage_data_f_1__48_;
   wire north_input_NIB_storage_data_f_1__49_;
   wire north_input_NIB_storage_data_f_1__50_;
   wire north_input_NIB_storage_data_f_1__51_;
   wire north_input_NIB_storage_data_f_1__52_;
   wire north_input_NIB_storage_data_f_1__53_;
   wire north_input_NIB_storage_data_f_1__54_;
   wire north_input_NIB_storage_data_f_1__55_;
   wire north_input_NIB_storage_data_f_1__56_;
   wire north_input_NIB_storage_data_f_1__57_;
   wire north_input_NIB_storage_data_f_1__58_;
   wire north_input_NIB_storage_data_f_1__59_;
   wire north_input_NIB_storage_data_f_1__60_;
   wire north_input_NIB_storage_data_f_1__61_;
   wire north_input_NIB_storage_data_f_1__62_;
   wire north_input_NIB_storage_data_f_1__63_;
   wire north_input_NIB_storage_data_f_0__0_;
   wire north_input_NIB_storage_data_f_0__1_;
   wire north_input_NIB_storage_data_f_0__2_;
   wire north_input_NIB_storage_data_f_0__3_;
   wire north_input_NIB_storage_data_f_0__4_;
   wire north_input_NIB_storage_data_f_0__5_;
   wire north_input_NIB_storage_data_f_0__6_;
   wire north_input_NIB_storage_data_f_0__7_;
   wire north_input_NIB_storage_data_f_0__8_;
   wire north_input_NIB_storage_data_f_0__9_;
   wire north_input_NIB_storage_data_f_0__10_;
   wire north_input_NIB_storage_data_f_0__11_;
   wire north_input_NIB_storage_data_f_0__12_;
   wire north_input_NIB_storage_data_f_0__13_;
   wire north_input_NIB_storage_data_f_0__14_;
   wire north_input_NIB_storage_data_f_0__15_;
   wire north_input_NIB_storage_data_f_0__16_;
   wire north_input_NIB_storage_data_f_0__17_;
   wire north_input_NIB_storage_data_f_0__18_;
   wire north_input_NIB_storage_data_f_0__19_;
   wire north_input_NIB_storage_data_f_0__20_;
   wire north_input_NIB_storage_data_f_0__21_;
   wire north_input_NIB_storage_data_f_0__22_;
   wire north_input_NIB_storage_data_f_0__23_;
   wire north_input_NIB_storage_data_f_0__24_;
   wire north_input_NIB_storage_data_f_0__25_;
   wire north_input_NIB_storage_data_f_0__26_;
   wire north_input_NIB_storage_data_f_0__27_;
   wire north_input_NIB_storage_data_f_0__28_;
   wire north_input_NIB_storage_data_f_0__29_;
   wire north_input_NIB_storage_data_f_0__30_;
   wire north_input_NIB_storage_data_f_0__31_;
   wire north_input_NIB_storage_data_f_0__32_;
   wire north_input_NIB_storage_data_f_0__33_;
   wire north_input_NIB_storage_data_f_0__34_;
   wire north_input_NIB_storage_data_f_0__35_;
   wire north_input_NIB_storage_data_f_0__36_;
   wire north_input_NIB_storage_data_f_0__37_;
   wire north_input_NIB_storage_data_f_0__38_;
   wire north_input_NIB_storage_data_f_0__39_;
   wire north_input_NIB_storage_data_f_0__40_;
   wire north_input_NIB_storage_data_f_0__41_;
   wire north_input_NIB_storage_data_f_0__42_;
   wire north_input_NIB_storage_data_f_0__43_;
   wire north_input_NIB_storage_data_f_0__44_;
   wire north_input_NIB_storage_data_f_0__45_;
   wire north_input_NIB_storage_data_f_0__46_;
   wire north_input_NIB_storage_data_f_0__47_;
   wire north_input_NIB_storage_data_f_0__48_;
   wire north_input_NIB_storage_data_f_0__49_;
   wire north_input_NIB_storage_data_f_0__50_;
   wire north_input_NIB_storage_data_f_0__51_;
   wire north_input_NIB_storage_data_f_0__52_;
   wire north_input_NIB_storage_data_f_0__53_;
   wire north_input_NIB_storage_data_f_0__54_;
   wire north_input_NIB_storage_data_f_0__55_;
   wire north_input_NIB_storage_data_f_0__56_;
   wire north_input_NIB_storage_data_f_0__57_;
   wire north_input_NIB_storage_data_f_0__58_;
   wire north_input_NIB_storage_data_f_0__59_;
   wire north_input_NIB_storage_data_f_0__60_;
   wire north_input_NIB_storage_data_f_0__61_;
   wire north_input_NIB_storage_data_f_0__62_;
   wire north_input_NIB_storage_data_f_0__63_;
   wire north_input_NIB_head_ptr_f_0_;
   wire north_input_NIB_head_ptr_f_1_;
   wire east_input_NIB_tail_ptr_f_0_;
   wire east_input_NIB_tail_ptr_f_1_;
   wire east_input_NIB_elements_in_array_f_0_;
   wire east_input_NIB_elements_in_array_f_1_;
   wire east_input_NIB_elements_in_array_f_2_;
   wire east_input_NIB_storage_data_f_3__0_;
   wire east_input_NIB_storage_data_f_3__1_;
   wire east_input_NIB_storage_data_f_3__2_;
   wire east_input_NIB_storage_data_f_3__3_;
   wire east_input_NIB_storage_data_f_3__4_;
   wire east_input_NIB_storage_data_f_3__5_;
   wire east_input_NIB_storage_data_f_3__6_;
   wire east_input_NIB_storage_data_f_3__7_;
   wire east_input_NIB_storage_data_f_3__8_;
   wire east_input_NIB_storage_data_f_3__9_;
   wire east_input_NIB_storage_data_f_3__10_;
   wire east_input_NIB_storage_data_f_3__11_;
   wire east_input_NIB_storage_data_f_3__12_;
   wire east_input_NIB_storage_data_f_3__13_;
   wire east_input_NIB_storage_data_f_3__14_;
   wire east_input_NIB_storage_data_f_3__15_;
   wire east_input_NIB_storage_data_f_3__16_;
   wire east_input_NIB_storage_data_f_3__17_;
   wire east_input_NIB_storage_data_f_3__18_;
   wire east_input_NIB_storage_data_f_3__19_;
   wire east_input_NIB_storage_data_f_3__20_;
   wire east_input_NIB_storage_data_f_3__21_;
   wire east_input_NIB_storage_data_f_3__22_;
   wire east_input_NIB_storage_data_f_3__23_;
   wire east_input_NIB_storage_data_f_3__24_;
   wire east_input_NIB_storage_data_f_3__25_;
   wire east_input_NIB_storage_data_f_3__26_;
   wire east_input_NIB_storage_data_f_3__27_;
   wire east_input_NIB_storage_data_f_3__28_;
   wire east_input_NIB_storage_data_f_3__29_;
   wire east_input_NIB_storage_data_f_3__30_;
   wire east_input_NIB_storage_data_f_3__31_;
   wire east_input_NIB_storage_data_f_3__32_;
   wire east_input_NIB_storage_data_f_3__33_;
   wire east_input_NIB_storage_data_f_3__34_;
   wire east_input_NIB_storage_data_f_3__35_;
   wire east_input_NIB_storage_data_f_3__36_;
   wire east_input_NIB_storage_data_f_3__37_;
   wire east_input_NIB_storage_data_f_3__38_;
   wire east_input_NIB_storage_data_f_3__39_;
   wire east_input_NIB_storage_data_f_3__40_;
   wire east_input_NIB_storage_data_f_3__41_;
   wire east_input_NIB_storage_data_f_3__42_;
   wire east_input_NIB_storage_data_f_3__43_;
   wire east_input_NIB_storage_data_f_3__44_;
   wire east_input_NIB_storage_data_f_3__45_;
   wire east_input_NIB_storage_data_f_3__46_;
   wire east_input_NIB_storage_data_f_3__47_;
   wire east_input_NIB_storage_data_f_3__48_;
   wire east_input_NIB_storage_data_f_3__49_;
   wire east_input_NIB_storage_data_f_3__50_;
   wire east_input_NIB_storage_data_f_3__51_;
   wire east_input_NIB_storage_data_f_3__52_;
   wire east_input_NIB_storage_data_f_3__53_;
   wire east_input_NIB_storage_data_f_3__54_;
   wire east_input_NIB_storage_data_f_3__55_;
   wire east_input_NIB_storage_data_f_3__56_;
   wire east_input_NIB_storage_data_f_3__57_;
   wire east_input_NIB_storage_data_f_3__58_;
   wire east_input_NIB_storage_data_f_3__59_;
   wire east_input_NIB_storage_data_f_3__60_;
   wire east_input_NIB_storage_data_f_3__61_;
   wire east_input_NIB_storage_data_f_3__62_;
   wire east_input_NIB_storage_data_f_3__63_;
   wire east_input_NIB_storage_data_f_2__0_;
   wire east_input_NIB_storage_data_f_2__1_;
   wire east_input_NIB_storage_data_f_2__2_;
   wire east_input_NIB_storage_data_f_2__3_;
   wire east_input_NIB_storage_data_f_2__4_;
   wire east_input_NIB_storage_data_f_2__5_;
   wire east_input_NIB_storage_data_f_2__6_;
   wire east_input_NIB_storage_data_f_2__7_;
   wire east_input_NIB_storage_data_f_2__8_;
   wire east_input_NIB_storage_data_f_2__9_;
   wire east_input_NIB_storage_data_f_2__10_;
   wire east_input_NIB_storage_data_f_2__11_;
   wire east_input_NIB_storage_data_f_2__12_;
   wire east_input_NIB_storage_data_f_2__13_;
   wire east_input_NIB_storage_data_f_2__14_;
   wire east_input_NIB_storage_data_f_2__15_;
   wire east_input_NIB_storage_data_f_2__16_;
   wire east_input_NIB_storage_data_f_2__17_;
   wire east_input_NIB_storage_data_f_2__18_;
   wire east_input_NIB_storage_data_f_2__19_;
   wire east_input_NIB_storage_data_f_2__20_;
   wire east_input_NIB_storage_data_f_2__21_;
   wire east_input_NIB_storage_data_f_2__22_;
   wire east_input_NIB_storage_data_f_2__23_;
   wire east_input_NIB_storage_data_f_2__24_;
   wire east_input_NIB_storage_data_f_2__25_;
   wire east_input_NIB_storage_data_f_2__26_;
   wire east_input_NIB_storage_data_f_2__27_;
   wire east_input_NIB_storage_data_f_2__28_;
   wire east_input_NIB_storage_data_f_2__29_;
   wire east_input_NIB_storage_data_f_2__30_;
   wire east_input_NIB_storage_data_f_2__31_;
   wire east_input_NIB_storage_data_f_2__32_;
   wire east_input_NIB_storage_data_f_2__33_;
   wire east_input_NIB_storage_data_f_2__34_;
   wire east_input_NIB_storage_data_f_2__35_;
   wire east_input_NIB_storage_data_f_2__36_;
   wire east_input_NIB_storage_data_f_2__37_;
   wire east_input_NIB_storage_data_f_2__38_;
   wire east_input_NIB_storage_data_f_2__39_;
   wire east_input_NIB_storage_data_f_2__40_;
   wire east_input_NIB_storage_data_f_2__41_;
   wire east_input_NIB_storage_data_f_2__42_;
   wire east_input_NIB_storage_data_f_2__43_;
   wire east_input_NIB_storage_data_f_2__44_;
   wire east_input_NIB_storage_data_f_2__45_;
   wire east_input_NIB_storage_data_f_2__46_;
   wire east_input_NIB_storage_data_f_2__47_;
   wire east_input_NIB_storage_data_f_2__48_;
   wire east_input_NIB_storage_data_f_2__49_;
   wire east_input_NIB_storage_data_f_2__50_;
   wire east_input_NIB_storage_data_f_2__51_;
   wire east_input_NIB_storage_data_f_2__52_;
   wire east_input_NIB_storage_data_f_2__53_;
   wire east_input_NIB_storage_data_f_2__54_;
   wire east_input_NIB_storage_data_f_2__55_;
   wire east_input_NIB_storage_data_f_2__56_;
   wire east_input_NIB_storage_data_f_2__57_;
   wire east_input_NIB_storage_data_f_2__58_;
   wire east_input_NIB_storage_data_f_2__59_;
   wire east_input_NIB_storage_data_f_2__60_;
   wire east_input_NIB_storage_data_f_2__61_;
   wire east_input_NIB_storage_data_f_2__62_;
   wire east_input_NIB_storage_data_f_2__63_;
   wire east_input_NIB_storage_data_f_1__0_;
   wire east_input_NIB_storage_data_f_1__1_;
   wire east_input_NIB_storage_data_f_1__2_;
   wire east_input_NIB_storage_data_f_1__3_;
   wire east_input_NIB_storage_data_f_1__4_;
   wire east_input_NIB_storage_data_f_1__5_;
   wire east_input_NIB_storage_data_f_1__6_;
   wire east_input_NIB_storage_data_f_1__7_;
   wire east_input_NIB_storage_data_f_1__8_;
   wire east_input_NIB_storage_data_f_1__9_;
   wire east_input_NIB_storage_data_f_1__10_;
   wire east_input_NIB_storage_data_f_1__11_;
   wire east_input_NIB_storage_data_f_1__12_;
   wire east_input_NIB_storage_data_f_1__13_;
   wire east_input_NIB_storage_data_f_1__14_;
   wire east_input_NIB_storage_data_f_1__15_;
   wire east_input_NIB_storage_data_f_1__16_;
   wire east_input_NIB_storage_data_f_1__17_;
   wire east_input_NIB_storage_data_f_1__18_;
   wire east_input_NIB_storage_data_f_1__19_;
   wire east_input_NIB_storage_data_f_1__20_;
   wire east_input_NIB_storage_data_f_1__21_;
   wire east_input_NIB_storage_data_f_1__22_;
   wire east_input_NIB_storage_data_f_1__23_;
   wire east_input_NIB_storage_data_f_1__24_;
   wire east_input_NIB_storage_data_f_1__25_;
   wire east_input_NIB_storage_data_f_1__26_;
   wire east_input_NIB_storage_data_f_1__27_;
   wire east_input_NIB_storage_data_f_1__28_;
   wire east_input_NIB_storage_data_f_1__29_;
   wire east_input_NIB_storage_data_f_1__30_;
   wire east_input_NIB_storage_data_f_1__31_;
   wire east_input_NIB_storage_data_f_1__32_;
   wire east_input_NIB_storage_data_f_1__33_;
   wire east_input_NIB_storage_data_f_1__34_;
   wire east_input_NIB_storage_data_f_1__35_;
   wire east_input_NIB_storage_data_f_1__36_;
   wire east_input_NIB_storage_data_f_1__37_;
   wire east_input_NIB_storage_data_f_1__38_;
   wire east_input_NIB_storage_data_f_1__39_;
   wire east_input_NIB_storage_data_f_1__40_;
   wire east_input_NIB_storage_data_f_1__41_;
   wire east_input_NIB_storage_data_f_1__42_;
   wire east_input_NIB_storage_data_f_1__43_;
   wire east_input_NIB_storage_data_f_1__44_;
   wire east_input_NIB_storage_data_f_1__45_;
   wire east_input_NIB_storage_data_f_1__46_;
   wire east_input_NIB_storage_data_f_1__47_;
   wire east_input_NIB_storage_data_f_1__48_;
   wire east_input_NIB_storage_data_f_1__49_;
   wire east_input_NIB_storage_data_f_1__50_;
   wire east_input_NIB_storage_data_f_1__51_;
   wire east_input_NIB_storage_data_f_1__52_;
   wire east_input_NIB_storage_data_f_1__53_;
   wire east_input_NIB_storage_data_f_1__54_;
   wire east_input_NIB_storage_data_f_1__55_;
   wire east_input_NIB_storage_data_f_1__56_;
   wire east_input_NIB_storage_data_f_1__57_;
   wire east_input_NIB_storage_data_f_1__58_;
   wire east_input_NIB_storage_data_f_1__59_;
   wire east_input_NIB_storage_data_f_1__60_;
   wire east_input_NIB_storage_data_f_1__61_;
   wire east_input_NIB_storage_data_f_1__62_;
   wire east_input_NIB_storage_data_f_1__63_;
   wire east_input_NIB_storage_data_f_0__0_;
   wire east_input_NIB_storage_data_f_0__1_;
   wire east_input_NIB_storage_data_f_0__2_;
   wire east_input_NIB_storage_data_f_0__3_;
   wire east_input_NIB_storage_data_f_0__4_;
   wire east_input_NIB_storage_data_f_0__5_;
   wire east_input_NIB_storage_data_f_0__6_;
   wire east_input_NIB_storage_data_f_0__7_;
   wire east_input_NIB_storage_data_f_0__8_;
   wire east_input_NIB_storage_data_f_0__9_;
   wire east_input_NIB_storage_data_f_0__10_;
   wire east_input_NIB_storage_data_f_0__11_;
   wire east_input_NIB_storage_data_f_0__12_;
   wire east_input_NIB_storage_data_f_0__13_;
   wire east_input_NIB_storage_data_f_0__14_;
   wire east_input_NIB_storage_data_f_0__15_;
   wire east_input_NIB_storage_data_f_0__16_;
   wire east_input_NIB_storage_data_f_0__17_;
   wire east_input_NIB_storage_data_f_0__18_;
   wire east_input_NIB_storage_data_f_0__19_;
   wire east_input_NIB_storage_data_f_0__20_;
   wire east_input_NIB_storage_data_f_0__21_;
   wire east_input_NIB_storage_data_f_0__22_;
   wire east_input_NIB_storage_data_f_0__23_;
   wire east_input_NIB_storage_data_f_0__24_;
   wire east_input_NIB_storage_data_f_0__25_;
   wire east_input_NIB_storage_data_f_0__26_;
   wire east_input_NIB_storage_data_f_0__27_;
   wire east_input_NIB_storage_data_f_0__28_;
   wire east_input_NIB_storage_data_f_0__29_;
   wire east_input_NIB_storage_data_f_0__30_;
   wire east_input_NIB_storage_data_f_0__31_;
   wire east_input_NIB_storage_data_f_0__32_;
   wire east_input_NIB_storage_data_f_0__33_;
   wire east_input_NIB_storage_data_f_0__34_;
   wire east_input_NIB_storage_data_f_0__35_;
   wire east_input_NIB_storage_data_f_0__36_;
   wire east_input_NIB_storage_data_f_0__37_;
   wire east_input_NIB_storage_data_f_0__38_;
   wire east_input_NIB_storage_data_f_0__39_;
   wire east_input_NIB_storage_data_f_0__40_;
   wire east_input_NIB_storage_data_f_0__41_;
   wire east_input_NIB_storage_data_f_0__42_;
   wire east_input_NIB_storage_data_f_0__43_;
   wire east_input_NIB_storage_data_f_0__44_;
   wire east_input_NIB_storage_data_f_0__45_;
   wire east_input_NIB_storage_data_f_0__46_;
   wire east_input_NIB_storage_data_f_0__47_;
   wire east_input_NIB_storage_data_f_0__48_;
   wire east_input_NIB_storage_data_f_0__49_;
   wire east_input_NIB_storage_data_f_0__50_;
   wire east_input_NIB_storage_data_f_0__51_;
   wire east_input_NIB_storage_data_f_0__52_;
   wire east_input_NIB_storage_data_f_0__53_;
   wire east_input_NIB_storage_data_f_0__54_;
   wire east_input_NIB_storage_data_f_0__55_;
   wire east_input_NIB_storage_data_f_0__56_;
   wire east_input_NIB_storage_data_f_0__57_;
   wire east_input_NIB_storage_data_f_0__58_;
   wire east_input_NIB_storage_data_f_0__59_;
   wire east_input_NIB_storage_data_f_0__60_;
   wire east_input_NIB_storage_data_f_0__61_;
   wire east_input_NIB_storage_data_f_0__62_;
   wire east_input_NIB_storage_data_f_0__63_;
   wire east_input_NIB_head_ptr_f_0_;
   wire east_input_NIB_head_ptr_f_1_;
   wire south_input_NIB_tail_ptr_f_0_;
   wire south_input_NIB_tail_ptr_f_1_;
   wire south_input_NIB_elements_in_array_f_0_;
   wire south_input_NIB_elements_in_array_f_1_;
   wire south_input_NIB_elements_in_array_f_2_;
   wire south_input_NIB_storage_data_f_3__0_;
   wire south_input_NIB_storage_data_f_3__1_;
   wire south_input_NIB_storage_data_f_3__2_;
   wire south_input_NIB_storage_data_f_3__3_;
   wire south_input_NIB_storage_data_f_3__4_;
   wire south_input_NIB_storage_data_f_3__5_;
   wire south_input_NIB_storage_data_f_3__6_;
   wire south_input_NIB_storage_data_f_3__7_;
   wire south_input_NIB_storage_data_f_3__8_;
   wire south_input_NIB_storage_data_f_3__9_;
   wire south_input_NIB_storage_data_f_3__10_;
   wire south_input_NIB_storage_data_f_3__11_;
   wire south_input_NIB_storage_data_f_3__12_;
   wire south_input_NIB_storage_data_f_3__13_;
   wire south_input_NIB_storage_data_f_3__14_;
   wire south_input_NIB_storage_data_f_3__15_;
   wire south_input_NIB_storage_data_f_3__16_;
   wire south_input_NIB_storage_data_f_3__17_;
   wire south_input_NIB_storage_data_f_3__18_;
   wire south_input_NIB_storage_data_f_3__19_;
   wire south_input_NIB_storage_data_f_3__20_;
   wire south_input_NIB_storage_data_f_3__21_;
   wire south_input_NIB_storage_data_f_3__22_;
   wire south_input_NIB_storage_data_f_3__23_;
   wire south_input_NIB_storage_data_f_3__24_;
   wire south_input_NIB_storage_data_f_3__25_;
   wire south_input_NIB_storage_data_f_3__26_;
   wire south_input_NIB_storage_data_f_3__27_;
   wire south_input_NIB_storage_data_f_3__28_;
   wire south_input_NIB_storage_data_f_3__29_;
   wire south_input_NIB_storage_data_f_3__30_;
   wire south_input_NIB_storage_data_f_3__31_;
   wire south_input_NIB_storage_data_f_3__32_;
   wire south_input_NIB_storage_data_f_3__33_;
   wire south_input_NIB_storage_data_f_3__34_;
   wire south_input_NIB_storage_data_f_3__35_;
   wire south_input_NIB_storage_data_f_3__36_;
   wire south_input_NIB_storage_data_f_3__37_;
   wire south_input_NIB_storage_data_f_3__38_;
   wire south_input_NIB_storage_data_f_3__39_;
   wire south_input_NIB_storage_data_f_3__40_;
   wire south_input_NIB_storage_data_f_3__41_;
   wire south_input_NIB_storage_data_f_3__42_;
   wire south_input_NIB_storage_data_f_3__43_;
   wire south_input_NIB_storage_data_f_3__44_;
   wire south_input_NIB_storage_data_f_3__45_;
   wire south_input_NIB_storage_data_f_3__46_;
   wire south_input_NIB_storage_data_f_3__47_;
   wire south_input_NIB_storage_data_f_3__48_;
   wire south_input_NIB_storage_data_f_3__49_;
   wire south_input_NIB_storage_data_f_3__50_;
   wire south_input_NIB_storage_data_f_3__51_;
   wire south_input_NIB_storage_data_f_3__52_;
   wire south_input_NIB_storage_data_f_3__53_;
   wire south_input_NIB_storage_data_f_3__54_;
   wire south_input_NIB_storage_data_f_3__55_;
   wire south_input_NIB_storage_data_f_3__56_;
   wire south_input_NIB_storage_data_f_3__57_;
   wire south_input_NIB_storage_data_f_3__58_;
   wire south_input_NIB_storage_data_f_3__59_;
   wire south_input_NIB_storage_data_f_3__60_;
   wire south_input_NIB_storage_data_f_3__61_;
   wire south_input_NIB_storage_data_f_3__62_;
   wire south_input_NIB_storage_data_f_3__63_;
   wire south_input_NIB_storage_data_f_2__0_;
   wire south_input_NIB_storage_data_f_2__1_;
   wire south_input_NIB_storage_data_f_2__2_;
   wire south_input_NIB_storage_data_f_2__3_;
   wire south_input_NIB_storage_data_f_2__4_;
   wire south_input_NIB_storage_data_f_2__5_;
   wire south_input_NIB_storage_data_f_2__6_;
   wire south_input_NIB_storage_data_f_2__7_;
   wire south_input_NIB_storage_data_f_2__8_;
   wire south_input_NIB_storage_data_f_2__9_;
   wire south_input_NIB_storage_data_f_2__10_;
   wire south_input_NIB_storage_data_f_2__11_;
   wire south_input_NIB_storage_data_f_2__12_;
   wire south_input_NIB_storage_data_f_2__13_;
   wire south_input_NIB_storage_data_f_2__14_;
   wire south_input_NIB_storage_data_f_2__15_;
   wire south_input_NIB_storage_data_f_2__16_;
   wire south_input_NIB_storage_data_f_2__17_;
   wire south_input_NIB_storage_data_f_2__18_;
   wire south_input_NIB_storage_data_f_2__19_;
   wire south_input_NIB_storage_data_f_2__20_;
   wire south_input_NIB_storage_data_f_2__21_;
   wire south_input_NIB_storage_data_f_2__22_;
   wire south_input_NIB_storage_data_f_2__23_;
   wire south_input_NIB_storage_data_f_2__24_;
   wire south_input_NIB_storage_data_f_2__25_;
   wire south_input_NIB_storage_data_f_2__26_;
   wire south_input_NIB_storage_data_f_2__27_;
   wire south_input_NIB_storage_data_f_2__28_;
   wire south_input_NIB_storage_data_f_2__29_;
   wire south_input_NIB_storage_data_f_2__30_;
   wire south_input_NIB_storage_data_f_2__31_;
   wire south_input_NIB_storage_data_f_2__32_;
   wire south_input_NIB_storage_data_f_2__33_;
   wire south_input_NIB_storage_data_f_2__34_;
   wire south_input_NIB_storage_data_f_2__35_;
   wire south_input_NIB_storage_data_f_2__36_;
   wire south_input_NIB_storage_data_f_2__37_;
   wire south_input_NIB_storage_data_f_2__38_;
   wire south_input_NIB_storage_data_f_2__39_;
   wire south_input_NIB_storage_data_f_2__40_;
   wire south_input_NIB_storage_data_f_2__41_;
   wire south_input_NIB_storage_data_f_2__42_;
   wire south_input_NIB_storage_data_f_2__43_;
   wire south_input_NIB_storage_data_f_2__44_;
   wire south_input_NIB_storage_data_f_2__45_;
   wire south_input_NIB_storage_data_f_2__46_;
   wire south_input_NIB_storage_data_f_2__47_;
   wire south_input_NIB_storage_data_f_2__48_;
   wire south_input_NIB_storage_data_f_2__49_;
   wire south_input_NIB_storage_data_f_2__50_;
   wire south_input_NIB_storage_data_f_2__51_;
   wire south_input_NIB_storage_data_f_2__52_;
   wire south_input_NIB_storage_data_f_2__53_;
   wire south_input_NIB_storage_data_f_2__54_;
   wire south_input_NIB_storage_data_f_2__55_;
   wire south_input_NIB_storage_data_f_2__56_;
   wire south_input_NIB_storage_data_f_2__57_;
   wire south_input_NIB_storage_data_f_2__58_;
   wire south_input_NIB_storage_data_f_2__59_;
   wire south_input_NIB_storage_data_f_2__60_;
   wire south_input_NIB_storage_data_f_2__61_;
   wire south_input_NIB_storage_data_f_2__62_;
   wire south_input_NIB_storage_data_f_2__63_;
   wire south_input_NIB_storage_data_f_1__0_;
   wire south_input_NIB_storage_data_f_1__1_;
   wire south_input_NIB_storage_data_f_1__2_;
   wire south_input_NIB_storage_data_f_1__3_;
   wire south_input_NIB_storage_data_f_1__4_;
   wire south_input_NIB_storage_data_f_1__5_;
   wire south_input_NIB_storage_data_f_1__6_;
   wire south_input_NIB_storage_data_f_1__7_;
   wire south_input_NIB_storage_data_f_1__8_;
   wire south_input_NIB_storage_data_f_1__9_;
   wire south_input_NIB_storage_data_f_1__10_;
   wire south_input_NIB_storage_data_f_1__11_;
   wire south_input_NIB_storage_data_f_1__12_;
   wire south_input_NIB_storage_data_f_1__13_;
   wire south_input_NIB_storage_data_f_1__14_;
   wire south_input_NIB_storage_data_f_1__15_;
   wire south_input_NIB_storage_data_f_1__16_;
   wire south_input_NIB_storage_data_f_1__17_;
   wire south_input_NIB_storage_data_f_1__18_;
   wire south_input_NIB_storage_data_f_1__19_;
   wire south_input_NIB_storage_data_f_1__20_;
   wire south_input_NIB_storage_data_f_1__21_;
   wire south_input_NIB_storage_data_f_1__22_;
   wire south_input_NIB_storage_data_f_1__23_;
   wire south_input_NIB_storage_data_f_1__24_;
   wire south_input_NIB_storage_data_f_1__25_;
   wire south_input_NIB_storage_data_f_1__26_;
   wire south_input_NIB_storage_data_f_1__27_;
   wire south_input_NIB_storage_data_f_1__28_;
   wire south_input_NIB_storage_data_f_1__29_;
   wire south_input_NIB_storage_data_f_1__30_;
   wire south_input_NIB_storage_data_f_1__31_;
   wire south_input_NIB_storage_data_f_1__32_;
   wire south_input_NIB_storage_data_f_1__33_;
   wire south_input_NIB_storage_data_f_1__34_;
   wire south_input_NIB_storage_data_f_1__35_;
   wire south_input_NIB_storage_data_f_1__36_;
   wire south_input_NIB_storage_data_f_1__37_;
   wire south_input_NIB_storage_data_f_1__38_;
   wire south_input_NIB_storage_data_f_1__39_;
   wire south_input_NIB_storage_data_f_1__40_;
   wire south_input_NIB_storage_data_f_1__41_;
   wire south_input_NIB_storage_data_f_1__42_;
   wire south_input_NIB_storage_data_f_1__43_;
   wire south_input_NIB_storage_data_f_1__44_;
   wire south_input_NIB_storage_data_f_1__45_;
   wire south_input_NIB_storage_data_f_1__46_;
   wire south_input_NIB_storage_data_f_1__47_;
   wire south_input_NIB_storage_data_f_1__48_;
   wire south_input_NIB_storage_data_f_1__49_;
   wire south_input_NIB_storage_data_f_1__50_;
   wire south_input_NIB_storage_data_f_1__51_;
   wire south_input_NIB_storage_data_f_1__52_;
   wire south_input_NIB_storage_data_f_1__53_;
   wire south_input_NIB_storage_data_f_1__54_;
   wire south_input_NIB_storage_data_f_1__55_;
   wire south_input_NIB_storage_data_f_1__56_;
   wire south_input_NIB_storage_data_f_1__57_;
   wire south_input_NIB_storage_data_f_1__58_;
   wire south_input_NIB_storage_data_f_1__59_;
   wire south_input_NIB_storage_data_f_1__60_;
   wire south_input_NIB_storage_data_f_1__61_;
   wire south_input_NIB_storage_data_f_1__62_;
   wire south_input_NIB_storage_data_f_1__63_;
   wire south_input_NIB_storage_data_f_0__0_;
   wire south_input_NIB_storage_data_f_0__1_;
   wire south_input_NIB_storage_data_f_0__2_;
   wire south_input_NIB_storage_data_f_0__3_;
   wire south_input_NIB_storage_data_f_0__4_;
   wire south_input_NIB_storage_data_f_0__5_;
   wire south_input_NIB_storage_data_f_0__6_;
   wire south_input_NIB_storage_data_f_0__7_;
   wire south_input_NIB_storage_data_f_0__8_;
   wire south_input_NIB_storage_data_f_0__9_;
   wire south_input_NIB_storage_data_f_0__10_;
   wire south_input_NIB_storage_data_f_0__11_;
   wire south_input_NIB_storage_data_f_0__12_;
   wire south_input_NIB_storage_data_f_0__13_;
   wire south_input_NIB_storage_data_f_0__14_;
   wire south_input_NIB_storage_data_f_0__15_;
   wire south_input_NIB_storage_data_f_0__16_;
   wire south_input_NIB_storage_data_f_0__17_;
   wire south_input_NIB_storage_data_f_0__18_;
   wire south_input_NIB_storage_data_f_0__19_;
   wire south_input_NIB_storage_data_f_0__20_;
   wire south_input_NIB_storage_data_f_0__21_;
   wire south_input_NIB_storage_data_f_0__22_;
   wire south_input_NIB_storage_data_f_0__23_;
   wire south_input_NIB_storage_data_f_0__24_;
   wire south_input_NIB_storage_data_f_0__25_;
   wire south_input_NIB_storage_data_f_0__26_;
   wire south_input_NIB_storage_data_f_0__27_;
   wire south_input_NIB_storage_data_f_0__28_;
   wire south_input_NIB_storage_data_f_0__29_;
   wire south_input_NIB_storage_data_f_0__30_;
   wire south_input_NIB_storage_data_f_0__31_;
   wire south_input_NIB_storage_data_f_0__32_;
   wire south_input_NIB_storage_data_f_0__33_;
   wire south_input_NIB_storage_data_f_0__34_;
   wire south_input_NIB_storage_data_f_0__35_;
   wire south_input_NIB_storage_data_f_0__36_;
   wire south_input_NIB_storage_data_f_0__37_;
   wire south_input_NIB_storage_data_f_0__38_;
   wire south_input_NIB_storage_data_f_0__39_;
   wire south_input_NIB_storage_data_f_0__40_;
   wire south_input_NIB_storage_data_f_0__41_;
   wire south_input_NIB_storage_data_f_0__42_;
   wire south_input_NIB_storage_data_f_0__43_;
   wire south_input_NIB_storage_data_f_0__44_;
   wire south_input_NIB_storage_data_f_0__45_;
   wire south_input_NIB_storage_data_f_0__46_;
   wire south_input_NIB_storage_data_f_0__47_;
   wire south_input_NIB_storage_data_f_0__48_;
   wire south_input_NIB_storage_data_f_0__49_;
   wire south_input_NIB_storage_data_f_0__50_;
   wire south_input_NIB_storage_data_f_0__51_;
   wire south_input_NIB_storage_data_f_0__52_;
   wire south_input_NIB_storage_data_f_0__53_;
   wire south_input_NIB_storage_data_f_0__54_;
   wire south_input_NIB_storage_data_f_0__55_;
   wire south_input_NIB_storage_data_f_0__56_;
   wire south_input_NIB_storage_data_f_0__57_;
   wire south_input_NIB_storage_data_f_0__58_;
   wire south_input_NIB_storage_data_f_0__59_;
   wire south_input_NIB_storage_data_f_0__60_;
   wire south_input_NIB_storage_data_f_0__61_;
   wire south_input_NIB_storage_data_f_0__62_;
   wire south_input_NIB_storage_data_f_0__63_;
   wire south_input_NIB_head_ptr_f_0_;
   wire south_input_NIB_head_ptr_f_1_;
   wire west_input_NIB_tail_ptr_f_0_;
   wire west_input_NIB_tail_ptr_f_1_;
   wire west_input_NIB_elements_in_array_f_0_;
   wire west_input_NIB_elements_in_array_f_1_;
   wire west_input_NIB_elements_in_array_f_2_;
   wire west_input_NIB_storage_data_f_3__0_;
   wire west_input_NIB_storage_data_f_3__1_;
   wire west_input_NIB_storage_data_f_3__2_;
   wire west_input_NIB_storage_data_f_3__3_;
   wire west_input_NIB_storage_data_f_3__4_;
   wire west_input_NIB_storage_data_f_3__5_;
   wire west_input_NIB_storage_data_f_3__6_;
   wire west_input_NIB_storage_data_f_3__7_;
   wire west_input_NIB_storage_data_f_3__8_;
   wire west_input_NIB_storage_data_f_3__9_;
   wire west_input_NIB_storage_data_f_3__10_;
   wire west_input_NIB_storage_data_f_3__11_;
   wire west_input_NIB_storage_data_f_3__12_;
   wire west_input_NIB_storage_data_f_3__13_;
   wire west_input_NIB_storage_data_f_3__14_;
   wire west_input_NIB_storage_data_f_3__15_;
   wire west_input_NIB_storage_data_f_3__16_;
   wire west_input_NIB_storage_data_f_3__17_;
   wire west_input_NIB_storage_data_f_3__18_;
   wire west_input_NIB_storage_data_f_3__19_;
   wire west_input_NIB_storage_data_f_3__20_;
   wire west_input_NIB_storage_data_f_3__21_;
   wire west_input_NIB_storage_data_f_3__22_;
   wire west_input_NIB_storage_data_f_3__23_;
   wire west_input_NIB_storage_data_f_3__24_;
   wire west_input_NIB_storage_data_f_3__25_;
   wire west_input_NIB_storage_data_f_3__26_;
   wire west_input_NIB_storage_data_f_3__27_;
   wire west_input_NIB_storage_data_f_3__28_;
   wire west_input_NIB_storage_data_f_3__29_;
   wire west_input_NIB_storage_data_f_3__30_;
   wire west_input_NIB_storage_data_f_3__31_;
   wire west_input_NIB_storage_data_f_3__32_;
   wire west_input_NIB_storage_data_f_3__33_;
   wire west_input_NIB_storage_data_f_3__34_;
   wire west_input_NIB_storage_data_f_3__35_;
   wire west_input_NIB_storage_data_f_3__36_;
   wire west_input_NIB_storage_data_f_3__37_;
   wire west_input_NIB_storage_data_f_3__38_;
   wire west_input_NIB_storage_data_f_3__39_;
   wire west_input_NIB_storage_data_f_3__40_;
   wire west_input_NIB_storage_data_f_3__41_;
   wire west_input_NIB_storage_data_f_3__42_;
   wire west_input_NIB_storage_data_f_3__43_;
   wire west_input_NIB_storage_data_f_3__44_;
   wire west_input_NIB_storage_data_f_3__45_;
   wire west_input_NIB_storage_data_f_3__46_;
   wire west_input_NIB_storage_data_f_3__47_;
   wire west_input_NIB_storage_data_f_3__48_;
   wire west_input_NIB_storage_data_f_3__49_;
   wire west_input_NIB_storage_data_f_3__50_;
   wire west_input_NIB_storage_data_f_3__51_;
   wire west_input_NIB_storage_data_f_3__52_;
   wire west_input_NIB_storage_data_f_3__53_;
   wire west_input_NIB_storage_data_f_3__54_;
   wire west_input_NIB_storage_data_f_3__55_;
   wire west_input_NIB_storage_data_f_3__56_;
   wire west_input_NIB_storage_data_f_3__57_;
   wire west_input_NIB_storage_data_f_3__58_;
   wire west_input_NIB_storage_data_f_3__59_;
   wire west_input_NIB_storage_data_f_3__60_;
   wire west_input_NIB_storage_data_f_3__61_;
   wire west_input_NIB_storage_data_f_3__62_;
   wire west_input_NIB_storage_data_f_3__63_;
   wire west_input_NIB_storage_data_f_2__0_;
   wire west_input_NIB_storage_data_f_2__1_;
   wire west_input_NIB_storage_data_f_2__2_;
   wire west_input_NIB_storage_data_f_2__3_;
   wire west_input_NIB_storage_data_f_2__4_;
   wire west_input_NIB_storage_data_f_2__5_;
   wire west_input_NIB_storage_data_f_2__6_;
   wire west_input_NIB_storage_data_f_2__7_;
   wire west_input_NIB_storage_data_f_2__8_;
   wire west_input_NIB_storage_data_f_2__9_;
   wire west_input_NIB_storage_data_f_2__10_;
   wire west_input_NIB_storage_data_f_2__11_;
   wire west_input_NIB_storage_data_f_2__12_;
   wire west_input_NIB_storage_data_f_2__13_;
   wire west_input_NIB_storage_data_f_2__14_;
   wire west_input_NIB_storage_data_f_2__15_;
   wire west_input_NIB_storage_data_f_2__16_;
   wire west_input_NIB_storage_data_f_2__17_;
   wire west_input_NIB_storage_data_f_2__18_;
   wire west_input_NIB_storage_data_f_2__19_;
   wire west_input_NIB_storage_data_f_2__20_;
   wire west_input_NIB_storage_data_f_2__21_;
   wire west_input_NIB_storage_data_f_2__22_;
   wire west_input_NIB_storage_data_f_2__23_;
   wire west_input_NIB_storage_data_f_2__24_;
   wire west_input_NIB_storage_data_f_2__25_;
   wire west_input_NIB_storage_data_f_2__26_;
   wire west_input_NIB_storage_data_f_2__27_;
   wire west_input_NIB_storage_data_f_2__28_;
   wire west_input_NIB_storage_data_f_2__29_;
   wire west_input_NIB_storage_data_f_2__30_;
   wire west_input_NIB_storage_data_f_2__31_;
   wire west_input_NIB_storage_data_f_2__32_;
   wire west_input_NIB_storage_data_f_2__33_;
   wire west_input_NIB_storage_data_f_2__34_;
   wire west_input_NIB_storage_data_f_2__35_;
   wire west_input_NIB_storage_data_f_2__36_;
   wire west_input_NIB_storage_data_f_2__37_;
   wire west_input_NIB_storage_data_f_2__38_;
   wire west_input_NIB_storage_data_f_2__39_;
   wire west_input_NIB_storage_data_f_2__40_;
   wire west_input_NIB_storage_data_f_2__41_;
   wire west_input_NIB_storage_data_f_2__42_;
   wire west_input_NIB_storage_data_f_2__43_;
   wire west_input_NIB_storage_data_f_2__44_;
   wire west_input_NIB_storage_data_f_2__45_;
   wire west_input_NIB_storage_data_f_2__46_;
   wire west_input_NIB_storage_data_f_2__47_;
   wire west_input_NIB_storage_data_f_2__48_;
   wire west_input_NIB_storage_data_f_2__49_;
   wire west_input_NIB_storage_data_f_2__50_;
   wire west_input_NIB_storage_data_f_2__51_;
   wire west_input_NIB_storage_data_f_2__52_;
   wire west_input_NIB_storage_data_f_2__53_;
   wire west_input_NIB_storage_data_f_2__54_;
   wire west_input_NIB_storage_data_f_2__55_;
   wire west_input_NIB_storage_data_f_2__56_;
   wire west_input_NIB_storage_data_f_2__57_;
   wire west_input_NIB_storage_data_f_2__58_;
   wire west_input_NIB_storage_data_f_2__59_;
   wire west_input_NIB_storage_data_f_2__60_;
   wire west_input_NIB_storage_data_f_2__61_;
   wire west_input_NIB_storage_data_f_2__62_;
   wire west_input_NIB_storage_data_f_2__63_;
   wire west_input_NIB_storage_data_f_1__0_;
   wire west_input_NIB_storage_data_f_1__1_;
   wire west_input_NIB_storage_data_f_1__2_;
   wire west_input_NIB_storage_data_f_1__3_;
   wire west_input_NIB_storage_data_f_1__4_;
   wire west_input_NIB_storage_data_f_1__5_;
   wire west_input_NIB_storage_data_f_1__6_;
   wire west_input_NIB_storage_data_f_1__7_;
   wire west_input_NIB_storage_data_f_1__8_;
   wire west_input_NIB_storage_data_f_1__9_;
   wire west_input_NIB_storage_data_f_1__10_;
   wire west_input_NIB_storage_data_f_1__11_;
   wire west_input_NIB_storage_data_f_1__12_;
   wire west_input_NIB_storage_data_f_1__13_;
   wire west_input_NIB_storage_data_f_1__14_;
   wire west_input_NIB_storage_data_f_1__15_;
   wire west_input_NIB_storage_data_f_1__16_;
   wire west_input_NIB_storage_data_f_1__17_;
   wire west_input_NIB_storage_data_f_1__18_;
   wire west_input_NIB_storage_data_f_1__19_;
   wire west_input_NIB_storage_data_f_1__20_;
   wire west_input_NIB_storage_data_f_1__21_;
   wire west_input_NIB_storage_data_f_1__22_;
   wire west_input_NIB_storage_data_f_1__23_;
   wire west_input_NIB_storage_data_f_1__24_;
   wire west_input_NIB_storage_data_f_1__25_;
   wire west_input_NIB_storage_data_f_1__26_;
   wire west_input_NIB_storage_data_f_1__27_;
   wire west_input_NIB_storage_data_f_1__28_;
   wire west_input_NIB_storage_data_f_1__29_;
   wire west_input_NIB_storage_data_f_1__30_;
   wire west_input_NIB_storage_data_f_1__31_;
   wire west_input_NIB_storage_data_f_1__32_;
   wire west_input_NIB_storage_data_f_1__33_;
   wire west_input_NIB_storage_data_f_1__34_;
   wire west_input_NIB_storage_data_f_1__35_;
   wire west_input_NIB_storage_data_f_1__36_;
   wire west_input_NIB_storage_data_f_1__37_;
   wire west_input_NIB_storage_data_f_1__38_;
   wire west_input_NIB_storage_data_f_1__39_;
   wire west_input_NIB_storage_data_f_1__40_;
   wire west_input_NIB_storage_data_f_1__41_;
   wire west_input_NIB_storage_data_f_1__42_;
   wire west_input_NIB_storage_data_f_1__43_;
   wire west_input_NIB_storage_data_f_1__44_;
   wire west_input_NIB_storage_data_f_1__45_;
   wire west_input_NIB_storage_data_f_1__46_;
   wire west_input_NIB_storage_data_f_1__47_;
   wire west_input_NIB_storage_data_f_1__48_;
   wire west_input_NIB_storage_data_f_1__49_;
   wire west_input_NIB_storage_data_f_1__50_;
   wire west_input_NIB_storage_data_f_1__51_;
   wire west_input_NIB_storage_data_f_1__52_;
   wire west_input_NIB_storage_data_f_1__53_;
   wire west_input_NIB_storage_data_f_1__54_;
   wire west_input_NIB_storage_data_f_1__55_;
   wire west_input_NIB_storage_data_f_1__56_;
   wire west_input_NIB_storage_data_f_1__57_;
   wire west_input_NIB_storage_data_f_1__58_;
   wire west_input_NIB_storage_data_f_1__59_;
   wire west_input_NIB_storage_data_f_1__60_;
   wire west_input_NIB_storage_data_f_1__61_;
   wire west_input_NIB_storage_data_f_1__62_;
   wire west_input_NIB_storage_data_f_1__63_;
   wire west_input_NIB_storage_data_f_0__0_;
   wire west_input_NIB_storage_data_f_0__1_;
   wire west_input_NIB_storage_data_f_0__2_;
   wire west_input_NIB_storage_data_f_0__3_;
   wire west_input_NIB_storage_data_f_0__4_;
   wire west_input_NIB_storage_data_f_0__5_;
   wire west_input_NIB_storage_data_f_0__6_;
   wire west_input_NIB_storage_data_f_0__7_;
   wire west_input_NIB_storage_data_f_0__8_;
   wire west_input_NIB_storage_data_f_0__9_;
   wire west_input_NIB_storage_data_f_0__10_;
   wire west_input_NIB_storage_data_f_0__11_;
   wire west_input_NIB_storage_data_f_0__12_;
   wire west_input_NIB_storage_data_f_0__13_;
   wire west_input_NIB_storage_data_f_0__14_;
   wire west_input_NIB_storage_data_f_0__15_;
   wire west_input_NIB_storage_data_f_0__16_;
   wire west_input_NIB_storage_data_f_0__17_;
   wire west_input_NIB_storage_data_f_0__18_;
   wire west_input_NIB_storage_data_f_0__19_;
   wire west_input_NIB_storage_data_f_0__20_;
   wire west_input_NIB_storage_data_f_0__21_;
   wire west_input_NIB_storage_data_f_0__22_;
   wire west_input_NIB_storage_data_f_0__23_;
   wire west_input_NIB_storage_data_f_0__24_;
   wire west_input_NIB_storage_data_f_0__25_;
   wire west_input_NIB_storage_data_f_0__26_;
   wire west_input_NIB_storage_data_f_0__27_;
   wire west_input_NIB_storage_data_f_0__28_;
   wire west_input_NIB_storage_data_f_0__29_;
   wire west_input_NIB_storage_data_f_0__30_;
   wire west_input_NIB_storage_data_f_0__31_;
   wire west_input_NIB_storage_data_f_0__32_;
   wire west_input_NIB_storage_data_f_0__33_;
   wire west_input_NIB_storage_data_f_0__34_;
   wire west_input_NIB_storage_data_f_0__35_;
   wire west_input_NIB_storage_data_f_0__36_;
   wire west_input_NIB_storage_data_f_0__37_;
   wire west_input_NIB_storage_data_f_0__38_;
   wire west_input_NIB_storage_data_f_0__39_;
   wire west_input_NIB_storage_data_f_0__40_;
   wire west_input_NIB_storage_data_f_0__41_;
   wire west_input_NIB_storage_data_f_0__42_;
   wire west_input_NIB_storage_data_f_0__43_;
   wire west_input_NIB_storage_data_f_0__44_;
   wire west_input_NIB_storage_data_f_0__45_;
   wire west_input_NIB_storage_data_f_0__46_;
   wire west_input_NIB_storage_data_f_0__47_;
   wire west_input_NIB_storage_data_f_0__48_;
   wire west_input_NIB_storage_data_f_0__49_;
   wire west_input_NIB_storage_data_f_0__50_;
   wire west_input_NIB_storage_data_f_0__51_;
   wire west_input_NIB_storage_data_f_0__52_;
   wire west_input_NIB_storage_data_f_0__53_;
   wire west_input_NIB_storage_data_f_0__54_;
   wire west_input_NIB_storage_data_f_0__55_;
   wire west_input_NIB_storage_data_f_0__56_;
   wire west_input_NIB_storage_data_f_0__57_;
   wire west_input_NIB_storage_data_f_0__58_;
   wire west_input_NIB_storage_data_f_0__59_;
   wire west_input_NIB_storage_data_f_0__60_;
   wire west_input_NIB_storage_data_f_0__61_;
   wire west_input_NIB_storage_data_f_0__62_;
   wire west_input_NIB_storage_data_f_0__63_;
   wire west_input_NIB_head_ptr_f_0_;
   wire west_input_NIB_head_ptr_f_1_;
   wire proc_input_NIB_tail_ptr_f_0_;
   wire proc_input_NIB_tail_ptr_f_1_;
   wire proc_input_NIB_tail_ptr_f_2_;
   wire proc_input_NIB_tail_ptr_f_3_;
   wire proc_input_NIB_elements_in_array_f_0_;
   wire proc_input_NIB_elements_in_array_f_1_;
   wire proc_input_NIB_elements_in_array_f_2_;
   wire proc_input_NIB_elements_in_array_f_3_;
   wire proc_input_NIB_elements_in_array_f_4_;
   wire proc_input_NIB_storage_data_f_15__0_;
   wire proc_input_NIB_storage_data_f_15__1_;
   wire proc_input_NIB_storage_data_f_15__2_;
   wire proc_input_NIB_storage_data_f_15__3_;
   wire proc_input_NIB_storage_data_f_15__4_;
   wire proc_input_NIB_storage_data_f_15__5_;
   wire proc_input_NIB_storage_data_f_15__6_;
   wire proc_input_NIB_storage_data_f_15__7_;
   wire proc_input_NIB_storage_data_f_15__8_;
   wire proc_input_NIB_storage_data_f_15__9_;
   wire proc_input_NIB_storage_data_f_15__10_;
   wire proc_input_NIB_storage_data_f_15__11_;
   wire proc_input_NIB_storage_data_f_15__12_;
   wire proc_input_NIB_storage_data_f_15__13_;
   wire proc_input_NIB_storage_data_f_15__14_;
   wire proc_input_NIB_storage_data_f_15__15_;
   wire proc_input_NIB_storage_data_f_15__16_;
   wire proc_input_NIB_storage_data_f_15__17_;
   wire proc_input_NIB_storage_data_f_15__18_;
   wire proc_input_NIB_storage_data_f_15__19_;
   wire proc_input_NIB_storage_data_f_15__20_;
   wire proc_input_NIB_storage_data_f_15__21_;
   wire proc_input_NIB_storage_data_f_15__22_;
   wire proc_input_NIB_storage_data_f_15__23_;
   wire proc_input_NIB_storage_data_f_15__24_;
   wire proc_input_NIB_storage_data_f_15__25_;
   wire proc_input_NIB_storage_data_f_15__26_;
   wire proc_input_NIB_storage_data_f_15__27_;
   wire proc_input_NIB_storage_data_f_15__28_;
   wire proc_input_NIB_storage_data_f_15__29_;
   wire proc_input_NIB_storage_data_f_15__30_;
   wire proc_input_NIB_storage_data_f_15__31_;
   wire proc_input_NIB_storage_data_f_15__32_;
   wire proc_input_NIB_storage_data_f_15__33_;
   wire proc_input_NIB_storage_data_f_15__34_;
   wire proc_input_NIB_storage_data_f_15__35_;
   wire proc_input_NIB_storage_data_f_15__36_;
   wire proc_input_NIB_storage_data_f_15__37_;
   wire proc_input_NIB_storage_data_f_15__38_;
   wire proc_input_NIB_storage_data_f_15__39_;
   wire proc_input_NIB_storage_data_f_15__40_;
   wire proc_input_NIB_storage_data_f_15__41_;
   wire proc_input_NIB_storage_data_f_15__42_;
   wire proc_input_NIB_storage_data_f_15__43_;
   wire proc_input_NIB_storage_data_f_15__44_;
   wire proc_input_NIB_storage_data_f_15__45_;
   wire proc_input_NIB_storage_data_f_15__46_;
   wire proc_input_NIB_storage_data_f_15__47_;
   wire proc_input_NIB_storage_data_f_15__48_;
   wire proc_input_NIB_storage_data_f_15__49_;
   wire proc_input_NIB_storage_data_f_15__50_;
   wire proc_input_NIB_storage_data_f_15__51_;
   wire proc_input_NIB_storage_data_f_15__52_;
   wire proc_input_NIB_storage_data_f_15__53_;
   wire proc_input_NIB_storage_data_f_15__54_;
   wire proc_input_NIB_storage_data_f_15__55_;
   wire proc_input_NIB_storage_data_f_15__56_;
   wire proc_input_NIB_storage_data_f_15__57_;
   wire proc_input_NIB_storage_data_f_15__58_;
   wire proc_input_NIB_storage_data_f_15__59_;
   wire proc_input_NIB_storage_data_f_15__60_;
   wire proc_input_NIB_storage_data_f_15__61_;
   wire proc_input_NIB_storage_data_f_15__62_;
   wire proc_input_NIB_storage_data_f_15__63_;
   wire proc_input_NIB_storage_data_f_14__0_;
   wire proc_input_NIB_storage_data_f_14__1_;
   wire proc_input_NIB_storage_data_f_14__2_;
   wire proc_input_NIB_storage_data_f_14__3_;
   wire proc_input_NIB_storage_data_f_14__4_;
   wire proc_input_NIB_storage_data_f_14__5_;
   wire proc_input_NIB_storage_data_f_14__6_;
   wire proc_input_NIB_storage_data_f_14__7_;
   wire proc_input_NIB_storage_data_f_14__8_;
   wire proc_input_NIB_storage_data_f_14__9_;
   wire proc_input_NIB_storage_data_f_14__10_;
   wire proc_input_NIB_storage_data_f_14__11_;
   wire proc_input_NIB_storage_data_f_14__12_;
   wire proc_input_NIB_storage_data_f_14__13_;
   wire proc_input_NIB_storage_data_f_14__14_;
   wire proc_input_NIB_storage_data_f_14__15_;
   wire proc_input_NIB_storage_data_f_14__16_;
   wire proc_input_NIB_storage_data_f_14__17_;
   wire proc_input_NIB_storage_data_f_14__18_;
   wire proc_input_NIB_storage_data_f_14__19_;
   wire proc_input_NIB_storage_data_f_14__20_;
   wire proc_input_NIB_storage_data_f_14__21_;
   wire proc_input_NIB_storage_data_f_14__22_;
   wire proc_input_NIB_storage_data_f_14__23_;
   wire proc_input_NIB_storage_data_f_14__24_;
   wire proc_input_NIB_storage_data_f_14__25_;
   wire proc_input_NIB_storage_data_f_14__26_;
   wire proc_input_NIB_storage_data_f_14__27_;
   wire proc_input_NIB_storage_data_f_14__28_;
   wire proc_input_NIB_storage_data_f_14__29_;
   wire proc_input_NIB_storage_data_f_14__30_;
   wire proc_input_NIB_storage_data_f_14__31_;
   wire proc_input_NIB_storage_data_f_14__32_;
   wire proc_input_NIB_storage_data_f_14__33_;
   wire proc_input_NIB_storage_data_f_14__34_;
   wire proc_input_NIB_storage_data_f_14__35_;
   wire proc_input_NIB_storage_data_f_14__36_;
   wire proc_input_NIB_storage_data_f_14__37_;
   wire proc_input_NIB_storage_data_f_14__38_;
   wire proc_input_NIB_storage_data_f_14__39_;
   wire proc_input_NIB_storage_data_f_14__40_;
   wire proc_input_NIB_storage_data_f_14__41_;
   wire proc_input_NIB_storage_data_f_14__42_;
   wire proc_input_NIB_storage_data_f_14__43_;
   wire proc_input_NIB_storage_data_f_14__44_;
   wire proc_input_NIB_storage_data_f_14__45_;
   wire proc_input_NIB_storage_data_f_14__46_;
   wire proc_input_NIB_storage_data_f_14__47_;
   wire proc_input_NIB_storage_data_f_14__48_;
   wire proc_input_NIB_storage_data_f_14__49_;
   wire proc_input_NIB_storage_data_f_14__50_;
   wire proc_input_NIB_storage_data_f_14__51_;
   wire proc_input_NIB_storage_data_f_14__52_;
   wire proc_input_NIB_storage_data_f_14__53_;
   wire proc_input_NIB_storage_data_f_14__54_;
   wire proc_input_NIB_storage_data_f_14__55_;
   wire proc_input_NIB_storage_data_f_14__56_;
   wire proc_input_NIB_storage_data_f_14__57_;
   wire proc_input_NIB_storage_data_f_14__58_;
   wire proc_input_NIB_storage_data_f_14__59_;
   wire proc_input_NIB_storage_data_f_14__60_;
   wire proc_input_NIB_storage_data_f_14__61_;
   wire proc_input_NIB_storage_data_f_14__62_;
   wire proc_input_NIB_storage_data_f_14__63_;
   wire proc_input_NIB_storage_data_f_13__0_;
   wire proc_input_NIB_storage_data_f_13__1_;
   wire proc_input_NIB_storage_data_f_13__2_;
   wire proc_input_NIB_storage_data_f_13__3_;
   wire proc_input_NIB_storage_data_f_13__4_;
   wire proc_input_NIB_storage_data_f_13__5_;
   wire proc_input_NIB_storage_data_f_13__6_;
   wire proc_input_NIB_storage_data_f_13__7_;
   wire proc_input_NIB_storage_data_f_13__8_;
   wire proc_input_NIB_storage_data_f_13__9_;
   wire proc_input_NIB_storage_data_f_13__10_;
   wire proc_input_NIB_storage_data_f_13__11_;
   wire proc_input_NIB_storage_data_f_13__12_;
   wire proc_input_NIB_storage_data_f_13__13_;
   wire proc_input_NIB_storage_data_f_13__14_;
   wire proc_input_NIB_storage_data_f_13__15_;
   wire proc_input_NIB_storage_data_f_13__16_;
   wire proc_input_NIB_storage_data_f_13__17_;
   wire proc_input_NIB_storage_data_f_13__18_;
   wire proc_input_NIB_storage_data_f_13__19_;
   wire proc_input_NIB_storage_data_f_13__20_;
   wire proc_input_NIB_storage_data_f_13__21_;
   wire proc_input_NIB_storage_data_f_13__22_;
   wire proc_input_NIB_storage_data_f_13__23_;
   wire proc_input_NIB_storage_data_f_13__24_;
   wire proc_input_NIB_storage_data_f_13__25_;
   wire proc_input_NIB_storage_data_f_13__26_;
   wire proc_input_NIB_storage_data_f_13__27_;
   wire proc_input_NIB_storage_data_f_13__28_;
   wire proc_input_NIB_storage_data_f_13__29_;
   wire proc_input_NIB_storage_data_f_13__30_;
   wire proc_input_NIB_storage_data_f_13__31_;
   wire proc_input_NIB_storage_data_f_13__32_;
   wire proc_input_NIB_storage_data_f_13__33_;
   wire proc_input_NIB_storage_data_f_13__34_;
   wire proc_input_NIB_storage_data_f_13__35_;
   wire proc_input_NIB_storage_data_f_13__36_;
   wire proc_input_NIB_storage_data_f_13__37_;
   wire proc_input_NIB_storage_data_f_13__38_;
   wire proc_input_NIB_storage_data_f_13__39_;
   wire proc_input_NIB_storage_data_f_13__40_;
   wire proc_input_NIB_storage_data_f_13__41_;
   wire proc_input_NIB_storage_data_f_13__42_;
   wire proc_input_NIB_storage_data_f_13__43_;
   wire proc_input_NIB_storage_data_f_13__44_;
   wire proc_input_NIB_storage_data_f_13__45_;
   wire proc_input_NIB_storage_data_f_13__46_;
   wire proc_input_NIB_storage_data_f_13__47_;
   wire proc_input_NIB_storage_data_f_13__48_;
   wire proc_input_NIB_storage_data_f_13__49_;
   wire proc_input_NIB_storage_data_f_13__50_;
   wire proc_input_NIB_storage_data_f_13__51_;
   wire proc_input_NIB_storage_data_f_13__52_;
   wire proc_input_NIB_storage_data_f_13__53_;
   wire proc_input_NIB_storage_data_f_13__54_;
   wire proc_input_NIB_storage_data_f_13__55_;
   wire proc_input_NIB_storage_data_f_13__56_;
   wire proc_input_NIB_storage_data_f_13__57_;
   wire proc_input_NIB_storage_data_f_13__58_;
   wire proc_input_NIB_storage_data_f_13__59_;
   wire proc_input_NIB_storage_data_f_13__60_;
   wire proc_input_NIB_storage_data_f_13__61_;
   wire proc_input_NIB_storage_data_f_13__62_;
   wire proc_input_NIB_storage_data_f_13__63_;
   wire proc_input_NIB_storage_data_f_12__0_;
   wire proc_input_NIB_storage_data_f_12__1_;
   wire proc_input_NIB_storage_data_f_12__2_;
   wire proc_input_NIB_storage_data_f_12__3_;
   wire proc_input_NIB_storage_data_f_12__4_;
   wire proc_input_NIB_storage_data_f_12__5_;
   wire proc_input_NIB_storage_data_f_12__6_;
   wire proc_input_NIB_storage_data_f_12__7_;
   wire proc_input_NIB_storage_data_f_12__8_;
   wire proc_input_NIB_storage_data_f_12__9_;
   wire proc_input_NIB_storage_data_f_12__10_;
   wire proc_input_NIB_storage_data_f_12__11_;
   wire proc_input_NIB_storage_data_f_12__12_;
   wire proc_input_NIB_storage_data_f_12__13_;
   wire proc_input_NIB_storage_data_f_12__14_;
   wire proc_input_NIB_storage_data_f_12__15_;
   wire proc_input_NIB_storage_data_f_12__16_;
   wire proc_input_NIB_storage_data_f_12__17_;
   wire proc_input_NIB_storage_data_f_12__18_;
   wire proc_input_NIB_storage_data_f_12__19_;
   wire proc_input_NIB_storage_data_f_12__20_;
   wire proc_input_NIB_storage_data_f_12__21_;
   wire proc_input_NIB_storage_data_f_12__22_;
   wire proc_input_NIB_storage_data_f_12__23_;
   wire proc_input_NIB_storage_data_f_12__24_;
   wire proc_input_NIB_storage_data_f_12__25_;
   wire proc_input_NIB_storage_data_f_12__26_;
   wire proc_input_NIB_storage_data_f_12__27_;
   wire proc_input_NIB_storage_data_f_12__28_;
   wire proc_input_NIB_storage_data_f_12__29_;
   wire proc_input_NIB_storage_data_f_12__30_;
   wire proc_input_NIB_storage_data_f_12__31_;
   wire proc_input_NIB_storage_data_f_12__32_;
   wire proc_input_NIB_storage_data_f_12__33_;
   wire proc_input_NIB_storage_data_f_12__34_;
   wire proc_input_NIB_storage_data_f_12__35_;
   wire proc_input_NIB_storage_data_f_12__36_;
   wire proc_input_NIB_storage_data_f_12__37_;
   wire proc_input_NIB_storage_data_f_12__38_;
   wire proc_input_NIB_storage_data_f_12__39_;
   wire proc_input_NIB_storage_data_f_12__40_;
   wire proc_input_NIB_storage_data_f_12__41_;
   wire proc_input_NIB_storage_data_f_12__42_;
   wire proc_input_NIB_storage_data_f_12__43_;
   wire proc_input_NIB_storage_data_f_12__44_;
   wire proc_input_NIB_storage_data_f_12__45_;
   wire proc_input_NIB_storage_data_f_12__46_;
   wire proc_input_NIB_storage_data_f_12__47_;
   wire proc_input_NIB_storage_data_f_12__48_;
   wire proc_input_NIB_storage_data_f_12__49_;
   wire proc_input_NIB_storage_data_f_12__50_;
   wire proc_input_NIB_storage_data_f_12__51_;
   wire proc_input_NIB_storage_data_f_12__52_;
   wire proc_input_NIB_storage_data_f_12__53_;
   wire proc_input_NIB_storage_data_f_12__54_;
   wire proc_input_NIB_storage_data_f_12__55_;
   wire proc_input_NIB_storage_data_f_12__56_;
   wire proc_input_NIB_storage_data_f_12__57_;
   wire proc_input_NIB_storage_data_f_12__58_;
   wire proc_input_NIB_storage_data_f_12__59_;
   wire proc_input_NIB_storage_data_f_12__60_;
   wire proc_input_NIB_storage_data_f_12__61_;
   wire proc_input_NIB_storage_data_f_12__62_;
   wire proc_input_NIB_storage_data_f_12__63_;
   wire proc_input_NIB_storage_data_f_11__0_;
   wire proc_input_NIB_storage_data_f_11__1_;
   wire proc_input_NIB_storage_data_f_11__2_;
   wire proc_input_NIB_storage_data_f_11__3_;
   wire proc_input_NIB_storage_data_f_11__4_;
   wire proc_input_NIB_storage_data_f_11__5_;
   wire proc_input_NIB_storage_data_f_11__6_;
   wire proc_input_NIB_storage_data_f_11__7_;
   wire proc_input_NIB_storage_data_f_11__8_;
   wire proc_input_NIB_storage_data_f_11__9_;
   wire proc_input_NIB_storage_data_f_11__10_;
   wire proc_input_NIB_storage_data_f_11__11_;
   wire proc_input_NIB_storage_data_f_11__12_;
   wire proc_input_NIB_storage_data_f_11__13_;
   wire proc_input_NIB_storage_data_f_11__14_;
   wire proc_input_NIB_storage_data_f_11__15_;
   wire proc_input_NIB_storage_data_f_11__16_;
   wire proc_input_NIB_storage_data_f_11__17_;
   wire proc_input_NIB_storage_data_f_11__18_;
   wire proc_input_NIB_storage_data_f_11__19_;
   wire proc_input_NIB_storage_data_f_11__20_;
   wire proc_input_NIB_storage_data_f_11__21_;
   wire proc_input_NIB_storage_data_f_11__22_;
   wire proc_input_NIB_storage_data_f_11__23_;
   wire proc_input_NIB_storage_data_f_11__24_;
   wire proc_input_NIB_storage_data_f_11__25_;
   wire proc_input_NIB_storage_data_f_11__26_;
   wire proc_input_NIB_storage_data_f_11__27_;
   wire proc_input_NIB_storage_data_f_11__28_;
   wire proc_input_NIB_storage_data_f_11__29_;
   wire proc_input_NIB_storage_data_f_11__30_;
   wire proc_input_NIB_storage_data_f_11__31_;
   wire proc_input_NIB_storage_data_f_11__32_;
   wire proc_input_NIB_storage_data_f_11__33_;
   wire proc_input_NIB_storage_data_f_11__34_;
   wire proc_input_NIB_storage_data_f_11__35_;
   wire proc_input_NIB_storage_data_f_11__36_;
   wire proc_input_NIB_storage_data_f_11__37_;
   wire proc_input_NIB_storage_data_f_11__38_;
   wire proc_input_NIB_storage_data_f_11__39_;
   wire proc_input_NIB_storage_data_f_11__40_;
   wire proc_input_NIB_storage_data_f_11__41_;
   wire proc_input_NIB_storage_data_f_11__42_;
   wire proc_input_NIB_storage_data_f_11__43_;
   wire proc_input_NIB_storage_data_f_11__44_;
   wire proc_input_NIB_storage_data_f_11__45_;
   wire proc_input_NIB_storage_data_f_11__46_;
   wire proc_input_NIB_storage_data_f_11__47_;
   wire proc_input_NIB_storage_data_f_11__48_;
   wire proc_input_NIB_storage_data_f_11__49_;
   wire proc_input_NIB_storage_data_f_11__50_;
   wire proc_input_NIB_storage_data_f_11__51_;
   wire proc_input_NIB_storage_data_f_11__52_;
   wire proc_input_NIB_storage_data_f_11__53_;
   wire proc_input_NIB_storage_data_f_11__54_;
   wire proc_input_NIB_storage_data_f_11__55_;
   wire proc_input_NIB_storage_data_f_11__56_;
   wire proc_input_NIB_storage_data_f_11__57_;
   wire proc_input_NIB_storage_data_f_11__58_;
   wire proc_input_NIB_storage_data_f_11__59_;
   wire proc_input_NIB_storage_data_f_11__60_;
   wire proc_input_NIB_storage_data_f_11__61_;
   wire proc_input_NIB_storage_data_f_11__62_;
   wire proc_input_NIB_storage_data_f_11__63_;
   wire proc_input_NIB_storage_data_f_10__0_;
   wire proc_input_NIB_storage_data_f_10__1_;
   wire proc_input_NIB_storage_data_f_10__2_;
   wire proc_input_NIB_storage_data_f_10__3_;
   wire proc_input_NIB_storage_data_f_10__4_;
   wire proc_input_NIB_storage_data_f_10__5_;
   wire proc_input_NIB_storage_data_f_10__6_;
   wire proc_input_NIB_storage_data_f_10__7_;
   wire proc_input_NIB_storage_data_f_10__8_;
   wire proc_input_NIB_storage_data_f_10__9_;
   wire proc_input_NIB_storage_data_f_10__10_;
   wire proc_input_NIB_storage_data_f_10__11_;
   wire proc_input_NIB_storage_data_f_10__12_;
   wire proc_input_NIB_storage_data_f_10__13_;
   wire proc_input_NIB_storage_data_f_10__14_;
   wire proc_input_NIB_storage_data_f_10__15_;
   wire proc_input_NIB_storage_data_f_10__16_;
   wire proc_input_NIB_storage_data_f_10__17_;
   wire proc_input_NIB_storage_data_f_10__18_;
   wire proc_input_NIB_storage_data_f_10__19_;
   wire proc_input_NIB_storage_data_f_10__20_;
   wire proc_input_NIB_storage_data_f_10__21_;
   wire proc_input_NIB_storage_data_f_10__22_;
   wire proc_input_NIB_storage_data_f_10__23_;
   wire proc_input_NIB_storage_data_f_10__24_;
   wire proc_input_NIB_storage_data_f_10__25_;
   wire proc_input_NIB_storage_data_f_10__26_;
   wire proc_input_NIB_storage_data_f_10__27_;
   wire proc_input_NIB_storage_data_f_10__28_;
   wire proc_input_NIB_storage_data_f_10__29_;
   wire proc_input_NIB_storage_data_f_10__30_;
   wire proc_input_NIB_storage_data_f_10__31_;
   wire proc_input_NIB_storage_data_f_10__32_;
   wire proc_input_NIB_storage_data_f_10__33_;
   wire proc_input_NIB_storage_data_f_10__34_;
   wire proc_input_NIB_storage_data_f_10__35_;
   wire proc_input_NIB_storage_data_f_10__36_;
   wire proc_input_NIB_storage_data_f_10__37_;
   wire proc_input_NIB_storage_data_f_10__38_;
   wire proc_input_NIB_storage_data_f_10__39_;
   wire proc_input_NIB_storage_data_f_10__40_;
   wire proc_input_NIB_storage_data_f_10__41_;
   wire proc_input_NIB_storage_data_f_10__42_;
   wire proc_input_NIB_storage_data_f_10__43_;
   wire proc_input_NIB_storage_data_f_10__44_;
   wire proc_input_NIB_storage_data_f_10__45_;
   wire proc_input_NIB_storage_data_f_10__46_;
   wire proc_input_NIB_storage_data_f_10__47_;
   wire proc_input_NIB_storage_data_f_10__48_;
   wire proc_input_NIB_storage_data_f_10__49_;
   wire proc_input_NIB_storage_data_f_10__50_;
   wire proc_input_NIB_storage_data_f_10__51_;
   wire proc_input_NIB_storage_data_f_10__52_;
   wire proc_input_NIB_storage_data_f_10__53_;
   wire proc_input_NIB_storage_data_f_10__54_;
   wire proc_input_NIB_storage_data_f_10__55_;
   wire proc_input_NIB_storage_data_f_10__56_;
   wire proc_input_NIB_storage_data_f_10__57_;
   wire proc_input_NIB_storage_data_f_10__58_;
   wire proc_input_NIB_storage_data_f_10__59_;
   wire proc_input_NIB_storage_data_f_10__60_;
   wire proc_input_NIB_storage_data_f_10__61_;
   wire proc_input_NIB_storage_data_f_10__62_;
   wire proc_input_NIB_storage_data_f_10__63_;
   wire proc_input_NIB_storage_data_f_9__0_;
   wire proc_input_NIB_storage_data_f_9__1_;
   wire proc_input_NIB_storage_data_f_9__2_;
   wire proc_input_NIB_storage_data_f_9__3_;
   wire proc_input_NIB_storage_data_f_9__4_;
   wire proc_input_NIB_storage_data_f_9__5_;
   wire proc_input_NIB_storage_data_f_9__6_;
   wire proc_input_NIB_storage_data_f_9__7_;
   wire proc_input_NIB_storage_data_f_9__8_;
   wire proc_input_NIB_storage_data_f_9__9_;
   wire proc_input_NIB_storage_data_f_9__10_;
   wire proc_input_NIB_storage_data_f_9__11_;
   wire proc_input_NIB_storage_data_f_9__12_;
   wire proc_input_NIB_storage_data_f_9__13_;
   wire proc_input_NIB_storage_data_f_9__14_;
   wire proc_input_NIB_storage_data_f_9__15_;
   wire proc_input_NIB_storage_data_f_9__16_;
   wire proc_input_NIB_storage_data_f_9__17_;
   wire proc_input_NIB_storage_data_f_9__18_;
   wire proc_input_NIB_storage_data_f_9__19_;
   wire proc_input_NIB_storage_data_f_9__20_;
   wire proc_input_NIB_storage_data_f_9__21_;
   wire proc_input_NIB_storage_data_f_9__22_;
   wire proc_input_NIB_storage_data_f_9__23_;
   wire proc_input_NIB_storage_data_f_9__24_;
   wire proc_input_NIB_storage_data_f_9__25_;
   wire proc_input_NIB_storage_data_f_9__26_;
   wire proc_input_NIB_storage_data_f_9__27_;
   wire proc_input_NIB_storage_data_f_9__28_;
   wire proc_input_NIB_storage_data_f_9__29_;
   wire proc_input_NIB_storage_data_f_9__30_;
   wire proc_input_NIB_storage_data_f_9__31_;
   wire proc_input_NIB_storage_data_f_9__32_;
   wire proc_input_NIB_storage_data_f_9__33_;
   wire proc_input_NIB_storage_data_f_9__34_;
   wire proc_input_NIB_storage_data_f_9__35_;
   wire proc_input_NIB_storage_data_f_9__36_;
   wire proc_input_NIB_storage_data_f_9__37_;
   wire proc_input_NIB_storage_data_f_9__38_;
   wire proc_input_NIB_storage_data_f_9__39_;
   wire proc_input_NIB_storage_data_f_9__40_;
   wire proc_input_NIB_storage_data_f_9__41_;
   wire proc_input_NIB_storage_data_f_9__42_;
   wire proc_input_NIB_storage_data_f_9__43_;
   wire proc_input_NIB_storage_data_f_9__44_;
   wire proc_input_NIB_storage_data_f_9__45_;
   wire proc_input_NIB_storage_data_f_9__46_;
   wire proc_input_NIB_storage_data_f_9__47_;
   wire proc_input_NIB_storage_data_f_9__48_;
   wire proc_input_NIB_storage_data_f_9__49_;
   wire proc_input_NIB_storage_data_f_9__50_;
   wire proc_input_NIB_storage_data_f_9__51_;
   wire proc_input_NIB_storage_data_f_9__52_;
   wire proc_input_NIB_storage_data_f_9__53_;
   wire proc_input_NIB_storage_data_f_9__54_;
   wire proc_input_NIB_storage_data_f_9__55_;
   wire proc_input_NIB_storage_data_f_9__56_;
   wire proc_input_NIB_storage_data_f_9__57_;
   wire proc_input_NIB_storage_data_f_9__58_;
   wire proc_input_NIB_storage_data_f_9__59_;
   wire proc_input_NIB_storage_data_f_9__60_;
   wire proc_input_NIB_storage_data_f_9__61_;
   wire proc_input_NIB_storage_data_f_9__62_;
   wire proc_input_NIB_storage_data_f_9__63_;
   wire proc_input_NIB_storage_data_f_8__0_;
   wire proc_input_NIB_storage_data_f_8__1_;
   wire proc_input_NIB_storage_data_f_8__2_;
   wire proc_input_NIB_storage_data_f_8__3_;
   wire proc_input_NIB_storage_data_f_8__4_;
   wire proc_input_NIB_storage_data_f_8__5_;
   wire proc_input_NIB_storage_data_f_8__6_;
   wire proc_input_NIB_storage_data_f_8__7_;
   wire proc_input_NIB_storage_data_f_8__8_;
   wire proc_input_NIB_storage_data_f_8__9_;
   wire proc_input_NIB_storage_data_f_8__10_;
   wire proc_input_NIB_storage_data_f_8__11_;
   wire proc_input_NIB_storage_data_f_8__12_;
   wire proc_input_NIB_storage_data_f_8__13_;
   wire proc_input_NIB_storage_data_f_8__14_;
   wire proc_input_NIB_storage_data_f_8__15_;
   wire proc_input_NIB_storage_data_f_8__16_;
   wire proc_input_NIB_storage_data_f_8__17_;
   wire proc_input_NIB_storage_data_f_8__18_;
   wire proc_input_NIB_storage_data_f_8__19_;
   wire proc_input_NIB_storage_data_f_8__20_;
   wire proc_input_NIB_storage_data_f_8__21_;
   wire proc_input_NIB_storage_data_f_8__22_;
   wire proc_input_NIB_storage_data_f_8__23_;
   wire proc_input_NIB_storage_data_f_8__24_;
   wire proc_input_NIB_storage_data_f_8__25_;
   wire proc_input_NIB_storage_data_f_8__26_;
   wire proc_input_NIB_storage_data_f_8__27_;
   wire proc_input_NIB_storage_data_f_8__28_;
   wire proc_input_NIB_storage_data_f_8__29_;
   wire proc_input_NIB_storage_data_f_8__30_;
   wire proc_input_NIB_storage_data_f_8__31_;
   wire proc_input_NIB_storage_data_f_8__32_;
   wire proc_input_NIB_storage_data_f_8__33_;
   wire proc_input_NIB_storage_data_f_8__34_;
   wire proc_input_NIB_storage_data_f_8__35_;
   wire proc_input_NIB_storage_data_f_8__36_;
   wire proc_input_NIB_storage_data_f_8__37_;
   wire proc_input_NIB_storage_data_f_8__38_;
   wire proc_input_NIB_storage_data_f_8__39_;
   wire proc_input_NIB_storage_data_f_8__40_;
   wire proc_input_NIB_storage_data_f_8__41_;
   wire proc_input_NIB_storage_data_f_8__42_;
   wire proc_input_NIB_storage_data_f_8__43_;
   wire proc_input_NIB_storage_data_f_8__44_;
   wire proc_input_NIB_storage_data_f_8__45_;
   wire proc_input_NIB_storage_data_f_8__46_;
   wire proc_input_NIB_storage_data_f_8__47_;
   wire proc_input_NIB_storage_data_f_8__48_;
   wire proc_input_NIB_storage_data_f_8__49_;
   wire proc_input_NIB_storage_data_f_8__50_;
   wire proc_input_NIB_storage_data_f_8__51_;
   wire proc_input_NIB_storage_data_f_8__52_;
   wire proc_input_NIB_storage_data_f_8__53_;
   wire proc_input_NIB_storage_data_f_8__54_;
   wire proc_input_NIB_storage_data_f_8__55_;
   wire proc_input_NIB_storage_data_f_8__56_;
   wire proc_input_NIB_storage_data_f_8__57_;
   wire proc_input_NIB_storage_data_f_8__58_;
   wire proc_input_NIB_storage_data_f_8__59_;
   wire proc_input_NIB_storage_data_f_8__60_;
   wire proc_input_NIB_storage_data_f_8__61_;
   wire proc_input_NIB_storage_data_f_8__62_;
   wire proc_input_NIB_storage_data_f_8__63_;
   wire proc_input_NIB_storage_data_f_7__0_;
   wire proc_input_NIB_storage_data_f_7__1_;
   wire proc_input_NIB_storage_data_f_7__2_;
   wire proc_input_NIB_storage_data_f_7__3_;
   wire proc_input_NIB_storage_data_f_7__4_;
   wire proc_input_NIB_storage_data_f_7__5_;
   wire proc_input_NIB_storage_data_f_7__6_;
   wire proc_input_NIB_storage_data_f_7__7_;
   wire proc_input_NIB_storage_data_f_7__8_;
   wire proc_input_NIB_storage_data_f_7__9_;
   wire proc_input_NIB_storage_data_f_7__10_;
   wire proc_input_NIB_storage_data_f_7__11_;
   wire proc_input_NIB_storage_data_f_7__12_;
   wire proc_input_NIB_storage_data_f_7__13_;
   wire proc_input_NIB_storage_data_f_7__14_;
   wire proc_input_NIB_storage_data_f_7__15_;
   wire proc_input_NIB_storage_data_f_7__16_;
   wire proc_input_NIB_storage_data_f_7__17_;
   wire proc_input_NIB_storage_data_f_7__18_;
   wire proc_input_NIB_storage_data_f_7__19_;
   wire proc_input_NIB_storage_data_f_7__20_;
   wire proc_input_NIB_storage_data_f_7__21_;
   wire proc_input_NIB_storage_data_f_7__22_;
   wire proc_input_NIB_storage_data_f_7__23_;
   wire proc_input_NIB_storage_data_f_7__24_;
   wire proc_input_NIB_storage_data_f_7__25_;
   wire proc_input_NIB_storage_data_f_7__26_;
   wire proc_input_NIB_storage_data_f_7__27_;
   wire proc_input_NIB_storage_data_f_7__28_;
   wire proc_input_NIB_storage_data_f_7__29_;
   wire proc_input_NIB_storage_data_f_7__30_;
   wire proc_input_NIB_storage_data_f_7__31_;
   wire proc_input_NIB_storage_data_f_7__32_;
   wire proc_input_NIB_storage_data_f_7__33_;
   wire proc_input_NIB_storage_data_f_7__34_;
   wire proc_input_NIB_storage_data_f_7__35_;
   wire proc_input_NIB_storage_data_f_7__36_;
   wire proc_input_NIB_storage_data_f_7__37_;
   wire proc_input_NIB_storage_data_f_7__38_;
   wire proc_input_NIB_storage_data_f_7__39_;
   wire proc_input_NIB_storage_data_f_7__40_;
   wire proc_input_NIB_storage_data_f_7__41_;
   wire proc_input_NIB_storage_data_f_7__42_;
   wire proc_input_NIB_storage_data_f_7__43_;
   wire proc_input_NIB_storage_data_f_7__44_;
   wire proc_input_NIB_storage_data_f_7__45_;
   wire proc_input_NIB_storage_data_f_7__46_;
   wire proc_input_NIB_storage_data_f_7__47_;
   wire proc_input_NIB_storage_data_f_7__48_;
   wire proc_input_NIB_storage_data_f_7__49_;
   wire proc_input_NIB_storage_data_f_7__50_;
   wire proc_input_NIB_storage_data_f_7__51_;
   wire proc_input_NIB_storage_data_f_7__52_;
   wire proc_input_NIB_storage_data_f_7__53_;
   wire proc_input_NIB_storage_data_f_7__54_;
   wire proc_input_NIB_storage_data_f_7__55_;
   wire proc_input_NIB_storage_data_f_7__56_;
   wire proc_input_NIB_storage_data_f_7__57_;
   wire proc_input_NIB_storage_data_f_7__58_;
   wire proc_input_NIB_storage_data_f_7__59_;
   wire proc_input_NIB_storage_data_f_7__60_;
   wire proc_input_NIB_storage_data_f_7__61_;
   wire proc_input_NIB_storage_data_f_7__62_;
   wire proc_input_NIB_storage_data_f_7__63_;
   wire proc_input_NIB_storage_data_f_6__0_;
   wire proc_input_NIB_storage_data_f_6__1_;
   wire proc_input_NIB_storage_data_f_6__2_;
   wire proc_input_NIB_storage_data_f_6__3_;
   wire proc_input_NIB_storage_data_f_6__4_;
   wire proc_input_NIB_storage_data_f_6__5_;
   wire proc_input_NIB_storage_data_f_6__6_;
   wire proc_input_NIB_storage_data_f_6__7_;
   wire proc_input_NIB_storage_data_f_6__8_;
   wire proc_input_NIB_storage_data_f_6__9_;
   wire proc_input_NIB_storage_data_f_6__10_;
   wire proc_input_NIB_storage_data_f_6__11_;
   wire proc_input_NIB_storage_data_f_6__12_;
   wire proc_input_NIB_storage_data_f_6__13_;
   wire proc_input_NIB_storage_data_f_6__14_;
   wire proc_input_NIB_storage_data_f_6__15_;
   wire proc_input_NIB_storage_data_f_6__16_;
   wire proc_input_NIB_storage_data_f_6__17_;
   wire proc_input_NIB_storage_data_f_6__18_;
   wire proc_input_NIB_storage_data_f_6__19_;
   wire proc_input_NIB_storage_data_f_6__20_;
   wire proc_input_NIB_storage_data_f_6__21_;
   wire proc_input_NIB_storage_data_f_6__22_;
   wire proc_input_NIB_storage_data_f_6__23_;
   wire proc_input_NIB_storage_data_f_6__24_;
   wire proc_input_NIB_storage_data_f_6__25_;
   wire proc_input_NIB_storage_data_f_6__26_;
   wire proc_input_NIB_storage_data_f_6__27_;
   wire proc_input_NIB_storage_data_f_6__28_;
   wire proc_input_NIB_storage_data_f_6__29_;
   wire proc_input_NIB_storage_data_f_6__30_;
   wire proc_input_NIB_storage_data_f_6__31_;
   wire proc_input_NIB_storage_data_f_6__32_;
   wire proc_input_NIB_storage_data_f_6__33_;
   wire proc_input_NIB_storage_data_f_6__34_;
   wire proc_input_NIB_storage_data_f_6__35_;
   wire proc_input_NIB_storage_data_f_6__36_;
   wire proc_input_NIB_storage_data_f_6__37_;
   wire proc_input_NIB_storage_data_f_6__38_;
   wire proc_input_NIB_storage_data_f_6__39_;
   wire proc_input_NIB_storage_data_f_6__40_;
   wire proc_input_NIB_storage_data_f_6__41_;
   wire proc_input_NIB_storage_data_f_6__42_;
   wire proc_input_NIB_storage_data_f_6__43_;
   wire proc_input_NIB_storage_data_f_6__44_;
   wire proc_input_NIB_storage_data_f_6__45_;
   wire proc_input_NIB_storage_data_f_6__46_;
   wire proc_input_NIB_storage_data_f_6__47_;
   wire proc_input_NIB_storage_data_f_6__48_;
   wire proc_input_NIB_storage_data_f_6__49_;
   wire proc_input_NIB_storage_data_f_6__50_;
   wire proc_input_NIB_storage_data_f_6__51_;
   wire proc_input_NIB_storage_data_f_6__52_;
   wire proc_input_NIB_storage_data_f_6__53_;
   wire proc_input_NIB_storage_data_f_6__54_;
   wire proc_input_NIB_storage_data_f_6__55_;
   wire proc_input_NIB_storage_data_f_6__56_;
   wire proc_input_NIB_storage_data_f_6__57_;
   wire proc_input_NIB_storage_data_f_6__58_;
   wire proc_input_NIB_storage_data_f_6__59_;
   wire proc_input_NIB_storage_data_f_6__60_;
   wire proc_input_NIB_storage_data_f_6__61_;
   wire proc_input_NIB_storage_data_f_6__62_;
   wire proc_input_NIB_storage_data_f_6__63_;
   wire proc_input_NIB_storage_data_f_5__0_;
   wire proc_input_NIB_storage_data_f_5__1_;
   wire proc_input_NIB_storage_data_f_5__2_;
   wire proc_input_NIB_storage_data_f_5__3_;
   wire proc_input_NIB_storage_data_f_5__4_;
   wire proc_input_NIB_storage_data_f_5__5_;
   wire proc_input_NIB_storage_data_f_5__6_;
   wire proc_input_NIB_storage_data_f_5__7_;
   wire proc_input_NIB_storage_data_f_5__8_;
   wire proc_input_NIB_storage_data_f_5__9_;
   wire proc_input_NIB_storage_data_f_5__10_;
   wire proc_input_NIB_storage_data_f_5__11_;
   wire proc_input_NIB_storage_data_f_5__12_;
   wire proc_input_NIB_storage_data_f_5__13_;
   wire proc_input_NIB_storage_data_f_5__14_;
   wire proc_input_NIB_storage_data_f_5__15_;
   wire proc_input_NIB_storage_data_f_5__16_;
   wire proc_input_NIB_storage_data_f_5__17_;
   wire proc_input_NIB_storage_data_f_5__18_;
   wire proc_input_NIB_storage_data_f_5__19_;
   wire proc_input_NIB_storage_data_f_5__20_;
   wire proc_input_NIB_storage_data_f_5__21_;
   wire proc_input_NIB_storage_data_f_5__22_;
   wire proc_input_NIB_storage_data_f_5__23_;
   wire proc_input_NIB_storage_data_f_5__24_;
   wire proc_input_NIB_storage_data_f_5__25_;
   wire proc_input_NIB_storage_data_f_5__26_;
   wire proc_input_NIB_storage_data_f_5__27_;
   wire proc_input_NIB_storage_data_f_5__28_;
   wire proc_input_NIB_storage_data_f_5__29_;
   wire proc_input_NIB_storage_data_f_5__30_;
   wire proc_input_NIB_storage_data_f_5__31_;
   wire proc_input_NIB_storage_data_f_5__32_;
   wire proc_input_NIB_storage_data_f_5__33_;
   wire proc_input_NIB_storage_data_f_5__34_;
   wire proc_input_NIB_storage_data_f_5__35_;
   wire proc_input_NIB_storage_data_f_5__36_;
   wire proc_input_NIB_storage_data_f_5__37_;
   wire proc_input_NIB_storage_data_f_5__38_;
   wire proc_input_NIB_storage_data_f_5__39_;
   wire proc_input_NIB_storage_data_f_5__40_;
   wire proc_input_NIB_storage_data_f_5__41_;
   wire proc_input_NIB_storage_data_f_5__42_;
   wire proc_input_NIB_storage_data_f_5__43_;
   wire proc_input_NIB_storage_data_f_5__44_;
   wire proc_input_NIB_storage_data_f_5__45_;
   wire proc_input_NIB_storage_data_f_5__46_;
   wire proc_input_NIB_storage_data_f_5__47_;
   wire proc_input_NIB_storage_data_f_5__48_;
   wire proc_input_NIB_storage_data_f_5__49_;
   wire proc_input_NIB_storage_data_f_5__50_;
   wire proc_input_NIB_storage_data_f_5__51_;
   wire proc_input_NIB_storage_data_f_5__52_;
   wire proc_input_NIB_storage_data_f_5__53_;
   wire proc_input_NIB_storage_data_f_5__54_;
   wire proc_input_NIB_storage_data_f_5__55_;
   wire proc_input_NIB_storage_data_f_5__56_;
   wire proc_input_NIB_storage_data_f_5__57_;
   wire proc_input_NIB_storage_data_f_5__58_;
   wire proc_input_NIB_storage_data_f_5__59_;
   wire proc_input_NIB_storage_data_f_5__60_;
   wire proc_input_NIB_storage_data_f_5__61_;
   wire proc_input_NIB_storage_data_f_5__62_;
   wire proc_input_NIB_storage_data_f_5__63_;
   wire proc_input_NIB_storage_data_f_4__0_;
   wire proc_input_NIB_storage_data_f_4__1_;
   wire proc_input_NIB_storage_data_f_4__2_;
   wire proc_input_NIB_storage_data_f_4__3_;
   wire proc_input_NIB_storage_data_f_4__4_;
   wire proc_input_NIB_storage_data_f_4__5_;
   wire proc_input_NIB_storage_data_f_4__6_;
   wire proc_input_NIB_storage_data_f_4__7_;
   wire proc_input_NIB_storage_data_f_4__8_;
   wire proc_input_NIB_storage_data_f_4__9_;
   wire proc_input_NIB_storage_data_f_4__10_;
   wire proc_input_NIB_storage_data_f_4__11_;
   wire proc_input_NIB_storage_data_f_4__12_;
   wire proc_input_NIB_storage_data_f_4__13_;
   wire proc_input_NIB_storage_data_f_4__14_;
   wire proc_input_NIB_storage_data_f_4__15_;
   wire proc_input_NIB_storage_data_f_4__16_;
   wire proc_input_NIB_storage_data_f_4__17_;
   wire proc_input_NIB_storage_data_f_4__18_;
   wire proc_input_NIB_storage_data_f_4__19_;
   wire proc_input_NIB_storage_data_f_4__20_;
   wire proc_input_NIB_storage_data_f_4__21_;
   wire proc_input_NIB_storage_data_f_4__22_;
   wire proc_input_NIB_storage_data_f_4__23_;
   wire proc_input_NIB_storage_data_f_4__24_;
   wire proc_input_NIB_storage_data_f_4__25_;
   wire proc_input_NIB_storage_data_f_4__26_;
   wire proc_input_NIB_storage_data_f_4__27_;
   wire proc_input_NIB_storage_data_f_4__28_;
   wire proc_input_NIB_storage_data_f_4__29_;
   wire proc_input_NIB_storage_data_f_4__30_;
   wire proc_input_NIB_storage_data_f_4__31_;
   wire proc_input_NIB_storage_data_f_4__32_;
   wire proc_input_NIB_storage_data_f_4__33_;
   wire proc_input_NIB_storage_data_f_4__34_;
   wire proc_input_NIB_storage_data_f_4__35_;
   wire proc_input_NIB_storage_data_f_4__36_;
   wire proc_input_NIB_storage_data_f_4__37_;
   wire proc_input_NIB_storage_data_f_4__38_;
   wire proc_input_NIB_storage_data_f_4__39_;
   wire proc_input_NIB_storage_data_f_4__40_;
   wire proc_input_NIB_storage_data_f_4__41_;
   wire proc_input_NIB_storage_data_f_4__42_;
   wire proc_input_NIB_storage_data_f_4__43_;
   wire proc_input_NIB_storage_data_f_4__44_;
   wire proc_input_NIB_storage_data_f_4__45_;
   wire proc_input_NIB_storage_data_f_4__46_;
   wire proc_input_NIB_storage_data_f_4__47_;
   wire proc_input_NIB_storage_data_f_4__48_;
   wire proc_input_NIB_storage_data_f_4__49_;
   wire proc_input_NIB_storage_data_f_4__50_;
   wire proc_input_NIB_storage_data_f_4__51_;
   wire proc_input_NIB_storage_data_f_4__52_;
   wire proc_input_NIB_storage_data_f_4__53_;
   wire proc_input_NIB_storage_data_f_4__54_;
   wire proc_input_NIB_storage_data_f_4__55_;
   wire proc_input_NIB_storage_data_f_4__56_;
   wire proc_input_NIB_storage_data_f_4__57_;
   wire proc_input_NIB_storage_data_f_4__58_;
   wire proc_input_NIB_storage_data_f_4__59_;
   wire proc_input_NIB_storage_data_f_4__60_;
   wire proc_input_NIB_storage_data_f_4__61_;
   wire proc_input_NIB_storage_data_f_4__62_;
   wire proc_input_NIB_storage_data_f_4__63_;
   wire proc_input_NIB_storage_data_f_3__0_;
   wire proc_input_NIB_storage_data_f_3__1_;
   wire proc_input_NIB_storage_data_f_3__2_;
   wire proc_input_NIB_storage_data_f_3__3_;
   wire proc_input_NIB_storage_data_f_3__4_;
   wire proc_input_NIB_storage_data_f_3__5_;
   wire proc_input_NIB_storage_data_f_3__6_;
   wire proc_input_NIB_storage_data_f_3__7_;
   wire proc_input_NIB_storage_data_f_3__8_;
   wire proc_input_NIB_storage_data_f_3__9_;
   wire proc_input_NIB_storage_data_f_3__10_;
   wire proc_input_NIB_storage_data_f_3__11_;
   wire proc_input_NIB_storage_data_f_3__12_;
   wire proc_input_NIB_storage_data_f_3__13_;
   wire proc_input_NIB_storage_data_f_3__14_;
   wire proc_input_NIB_storage_data_f_3__15_;
   wire proc_input_NIB_storage_data_f_3__16_;
   wire proc_input_NIB_storage_data_f_3__17_;
   wire proc_input_NIB_storage_data_f_3__18_;
   wire proc_input_NIB_storage_data_f_3__19_;
   wire proc_input_NIB_storage_data_f_3__20_;
   wire proc_input_NIB_storage_data_f_3__21_;
   wire proc_input_NIB_storage_data_f_3__22_;
   wire proc_input_NIB_storage_data_f_3__23_;
   wire proc_input_NIB_storage_data_f_3__24_;
   wire proc_input_NIB_storage_data_f_3__25_;
   wire proc_input_NIB_storage_data_f_3__26_;
   wire proc_input_NIB_storage_data_f_3__27_;
   wire proc_input_NIB_storage_data_f_3__28_;
   wire proc_input_NIB_storage_data_f_3__29_;
   wire proc_input_NIB_storage_data_f_3__30_;
   wire proc_input_NIB_storage_data_f_3__31_;
   wire proc_input_NIB_storage_data_f_3__32_;
   wire proc_input_NIB_storage_data_f_3__33_;
   wire proc_input_NIB_storage_data_f_3__34_;
   wire proc_input_NIB_storage_data_f_3__35_;
   wire proc_input_NIB_storage_data_f_3__36_;
   wire proc_input_NIB_storage_data_f_3__37_;
   wire proc_input_NIB_storage_data_f_3__38_;
   wire proc_input_NIB_storage_data_f_3__39_;
   wire proc_input_NIB_storage_data_f_3__40_;
   wire proc_input_NIB_storage_data_f_3__41_;
   wire proc_input_NIB_storage_data_f_3__42_;
   wire proc_input_NIB_storage_data_f_3__43_;
   wire proc_input_NIB_storage_data_f_3__44_;
   wire proc_input_NIB_storage_data_f_3__45_;
   wire proc_input_NIB_storage_data_f_3__46_;
   wire proc_input_NIB_storage_data_f_3__47_;
   wire proc_input_NIB_storage_data_f_3__48_;
   wire proc_input_NIB_storage_data_f_3__49_;
   wire proc_input_NIB_storage_data_f_3__50_;
   wire proc_input_NIB_storage_data_f_3__51_;
   wire proc_input_NIB_storage_data_f_3__52_;
   wire proc_input_NIB_storage_data_f_3__53_;
   wire proc_input_NIB_storage_data_f_3__54_;
   wire proc_input_NIB_storage_data_f_3__55_;
   wire proc_input_NIB_storage_data_f_3__56_;
   wire proc_input_NIB_storage_data_f_3__57_;
   wire proc_input_NIB_storage_data_f_3__58_;
   wire proc_input_NIB_storage_data_f_3__59_;
   wire proc_input_NIB_storage_data_f_3__60_;
   wire proc_input_NIB_storage_data_f_3__61_;
   wire proc_input_NIB_storage_data_f_3__62_;
   wire proc_input_NIB_storage_data_f_3__63_;
   wire proc_input_NIB_storage_data_f_2__0_;
   wire proc_input_NIB_storage_data_f_2__1_;
   wire proc_input_NIB_storage_data_f_2__2_;
   wire proc_input_NIB_storage_data_f_2__3_;
   wire proc_input_NIB_storage_data_f_2__4_;
   wire proc_input_NIB_storage_data_f_2__5_;
   wire proc_input_NIB_storage_data_f_2__6_;
   wire proc_input_NIB_storage_data_f_2__7_;
   wire proc_input_NIB_storage_data_f_2__8_;
   wire proc_input_NIB_storage_data_f_2__9_;
   wire proc_input_NIB_storage_data_f_2__10_;
   wire proc_input_NIB_storage_data_f_2__11_;
   wire proc_input_NIB_storage_data_f_2__12_;
   wire proc_input_NIB_storage_data_f_2__13_;
   wire proc_input_NIB_storage_data_f_2__14_;
   wire proc_input_NIB_storage_data_f_2__15_;
   wire proc_input_NIB_storage_data_f_2__16_;
   wire proc_input_NIB_storage_data_f_2__17_;
   wire proc_input_NIB_storage_data_f_2__18_;
   wire proc_input_NIB_storage_data_f_2__19_;
   wire proc_input_NIB_storage_data_f_2__20_;
   wire proc_input_NIB_storage_data_f_2__21_;
   wire proc_input_NIB_storage_data_f_2__22_;
   wire proc_input_NIB_storage_data_f_2__23_;
   wire proc_input_NIB_storage_data_f_2__24_;
   wire proc_input_NIB_storage_data_f_2__25_;
   wire proc_input_NIB_storage_data_f_2__26_;
   wire proc_input_NIB_storage_data_f_2__27_;
   wire proc_input_NIB_storage_data_f_2__28_;
   wire proc_input_NIB_storage_data_f_2__29_;
   wire proc_input_NIB_storage_data_f_2__30_;
   wire proc_input_NIB_storage_data_f_2__31_;
   wire proc_input_NIB_storage_data_f_2__32_;
   wire proc_input_NIB_storage_data_f_2__33_;
   wire proc_input_NIB_storage_data_f_2__34_;
   wire proc_input_NIB_storage_data_f_2__35_;
   wire proc_input_NIB_storage_data_f_2__36_;
   wire proc_input_NIB_storage_data_f_2__37_;
   wire proc_input_NIB_storage_data_f_2__38_;
   wire proc_input_NIB_storage_data_f_2__39_;
   wire proc_input_NIB_storage_data_f_2__40_;
   wire proc_input_NIB_storage_data_f_2__41_;
   wire proc_input_NIB_storage_data_f_2__42_;
   wire proc_input_NIB_storage_data_f_2__43_;
   wire proc_input_NIB_storage_data_f_2__44_;
   wire proc_input_NIB_storage_data_f_2__45_;
   wire proc_input_NIB_storage_data_f_2__46_;
   wire proc_input_NIB_storage_data_f_2__47_;
   wire proc_input_NIB_storage_data_f_2__48_;
   wire proc_input_NIB_storage_data_f_2__49_;
   wire proc_input_NIB_storage_data_f_2__50_;
   wire proc_input_NIB_storage_data_f_2__51_;
   wire proc_input_NIB_storage_data_f_2__52_;
   wire proc_input_NIB_storage_data_f_2__53_;
   wire proc_input_NIB_storage_data_f_2__54_;
   wire proc_input_NIB_storage_data_f_2__55_;
   wire proc_input_NIB_storage_data_f_2__56_;
   wire proc_input_NIB_storage_data_f_2__57_;
   wire proc_input_NIB_storage_data_f_2__58_;
   wire proc_input_NIB_storage_data_f_2__59_;
   wire proc_input_NIB_storage_data_f_2__60_;
   wire proc_input_NIB_storage_data_f_2__61_;
   wire proc_input_NIB_storage_data_f_2__62_;
   wire proc_input_NIB_storage_data_f_2__63_;
   wire proc_input_NIB_storage_data_f_1__0_;
   wire proc_input_NIB_storage_data_f_1__1_;
   wire proc_input_NIB_storage_data_f_1__2_;
   wire proc_input_NIB_storage_data_f_1__3_;
   wire proc_input_NIB_storage_data_f_1__4_;
   wire proc_input_NIB_storage_data_f_1__5_;
   wire proc_input_NIB_storage_data_f_1__6_;
   wire proc_input_NIB_storage_data_f_1__7_;
   wire proc_input_NIB_storage_data_f_1__8_;
   wire proc_input_NIB_storage_data_f_1__9_;
   wire proc_input_NIB_storage_data_f_1__10_;
   wire proc_input_NIB_storage_data_f_1__11_;
   wire proc_input_NIB_storage_data_f_1__12_;
   wire proc_input_NIB_storage_data_f_1__13_;
   wire proc_input_NIB_storage_data_f_1__14_;
   wire proc_input_NIB_storage_data_f_1__15_;
   wire proc_input_NIB_storage_data_f_1__16_;
   wire proc_input_NIB_storage_data_f_1__17_;
   wire proc_input_NIB_storage_data_f_1__18_;
   wire proc_input_NIB_storage_data_f_1__19_;
   wire proc_input_NIB_storage_data_f_1__20_;
   wire proc_input_NIB_storage_data_f_1__21_;
   wire proc_input_NIB_storage_data_f_1__22_;
   wire proc_input_NIB_storage_data_f_1__23_;
   wire proc_input_NIB_storage_data_f_1__24_;
   wire proc_input_NIB_storage_data_f_1__25_;
   wire proc_input_NIB_storage_data_f_1__26_;
   wire proc_input_NIB_storage_data_f_1__27_;
   wire proc_input_NIB_storage_data_f_1__28_;
   wire proc_input_NIB_storage_data_f_1__29_;
   wire proc_input_NIB_storage_data_f_1__30_;
   wire proc_input_NIB_storage_data_f_1__31_;
   wire proc_input_NIB_storage_data_f_1__32_;
   wire proc_input_NIB_storage_data_f_1__33_;
   wire proc_input_NIB_storage_data_f_1__34_;
   wire proc_input_NIB_storage_data_f_1__35_;
   wire proc_input_NIB_storage_data_f_1__36_;
   wire proc_input_NIB_storage_data_f_1__37_;
   wire proc_input_NIB_storage_data_f_1__38_;
   wire proc_input_NIB_storage_data_f_1__39_;
   wire proc_input_NIB_storage_data_f_1__40_;
   wire proc_input_NIB_storage_data_f_1__41_;
   wire proc_input_NIB_storage_data_f_1__42_;
   wire proc_input_NIB_storage_data_f_1__43_;
   wire proc_input_NIB_storage_data_f_1__44_;
   wire proc_input_NIB_storage_data_f_1__45_;
   wire proc_input_NIB_storage_data_f_1__46_;
   wire proc_input_NIB_storage_data_f_1__47_;
   wire proc_input_NIB_storage_data_f_1__48_;
   wire proc_input_NIB_storage_data_f_1__49_;
   wire proc_input_NIB_storage_data_f_1__50_;
   wire proc_input_NIB_storage_data_f_1__51_;
   wire proc_input_NIB_storage_data_f_1__52_;
   wire proc_input_NIB_storage_data_f_1__53_;
   wire proc_input_NIB_storage_data_f_1__54_;
   wire proc_input_NIB_storage_data_f_1__55_;
   wire proc_input_NIB_storage_data_f_1__56_;
   wire proc_input_NIB_storage_data_f_1__57_;
   wire proc_input_NIB_storage_data_f_1__58_;
   wire proc_input_NIB_storage_data_f_1__59_;
   wire proc_input_NIB_storage_data_f_1__60_;
   wire proc_input_NIB_storage_data_f_1__61_;
   wire proc_input_NIB_storage_data_f_1__62_;
   wire proc_input_NIB_storage_data_f_1__63_;
   wire proc_input_NIB_storage_data_f_0__0_;
   wire proc_input_NIB_storage_data_f_0__1_;
   wire proc_input_NIB_storage_data_f_0__2_;
   wire proc_input_NIB_storage_data_f_0__3_;
   wire proc_input_NIB_storage_data_f_0__4_;
   wire proc_input_NIB_storage_data_f_0__5_;
   wire proc_input_NIB_storage_data_f_0__6_;
   wire proc_input_NIB_storage_data_f_0__7_;
   wire proc_input_NIB_storage_data_f_0__8_;
   wire proc_input_NIB_storage_data_f_0__9_;
   wire proc_input_NIB_storage_data_f_0__10_;
   wire proc_input_NIB_storage_data_f_0__11_;
   wire proc_input_NIB_storage_data_f_0__12_;
   wire proc_input_NIB_storage_data_f_0__13_;
   wire proc_input_NIB_storage_data_f_0__14_;
   wire proc_input_NIB_storage_data_f_0__15_;
   wire proc_input_NIB_storage_data_f_0__16_;
   wire proc_input_NIB_storage_data_f_0__17_;
   wire proc_input_NIB_storage_data_f_0__18_;
   wire proc_input_NIB_storage_data_f_0__19_;
   wire proc_input_NIB_storage_data_f_0__20_;
   wire proc_input_NIB_storage_data_f_0__21_;
   wire proc_input_NIB_storage_data_f_0__22_;
   wire proc_input_NIB_storage_data_f_0__23_;
   wire proc_input_NIB_storage_data_f_0__24_;
   wire proc_input_NIB_storage_data_f_0__25_;
   wire proc_input_NIB_storage_data_f_0__26_;
   wire proc_input_NIB_storage_data_f_0__27_;
   wire proc_input_NIB_storage_data_f_0__28_;
   wire proc_input_NIB_storage_data_f_0__29_;
   wire proc_input_NIB_storage_data_f_0__30_;
   wire proc_input_NIB_storage_data_f_0__31_;
   wire proc_input_NIB_storage_data_f_0__32_;
   wire proc_input_NIB_storage_data_f_0__33_;
   wire proc_input_NIB_storage_data_f_0__34_;
   wire proc_input_NIB_storage_data_f_0__35_;
   wire proc_input_NIB_storage_data_f_0__36_;
   wire proc_input_NIB_storage_data_f_0__37_;
   wire proc_input_NIB_storage_data_f_0__38_;
   wire proc_input_NIB_storage_data_f_0__39_;
   wire proc_input_NIB_storage_data_f_0__40_;
   wire proc_input_NIB_storage_data_f_0__41_;
   wire proc_input_NIB_storage_data_f_0__42_;
   wire proc_input_NIB_storage_data_f_0__43_;
   wire proc_input_NIB_storage_data_f_0__44_;
   wire proc_input_NIB_storage_data_f_0__45_;
   wire proc_input_NIB_storage_data_f_0__46_;
   wire proc_input_NIB_storage_data_f_0__47_;
   wire proc_input_NIB_storage_data_f_0__48_;
   wire proc_input_NIB_storage_data_f_0__49_;
   wire proc_input_NIB_storage_data_f_0__50_;
   wire proc_input_NIB_storage_data_f_0__51_;
   wire proc_input_NIB_storage_data_f_0__52_;
   wire proc_input_NIB_storage_data_f_0__53_;
   wire proc_input_NIB_storage_data_f_0__54_;
   wire proc_input_NIB_storage_data_f_0__55_;
   wire proc_input_NIB_storage_data_f_0__56_;
   wire proc_input_NIB_storage_data_f_0__57_;
   wire proc_input_NIB_storage_data_f_0__58_;
   wire proc_input_NIB_storage_data_f_0__59_;
   wire proc_input_NIB_storage_data_f_0__60_;
   wire proc_input_NIB_storage_data_f_0__61_;
   wire proc_input_NIB_storage_data_f_0__62_;
   wire proc_input_NIB_storage_data_f_0__63_;
   wire proc_input_NIB_head_ptr_f_0_;
   wire proc_input_NIB_head_ptr_f_1_;
   wire proc_input_NIB_head_ptr_f_2_;
   wire proc_input_NIB_head_ptr_f_3_;
   wire north_input_control_N53;
   wire north_input_control_N52;
   wire north_input_control_N51;
   wire north_input_control_N49;
   wire north_input_control_N48;
   wire north_input_control_N47;
   wire north_input_control_N46;
   wire north_input_control_N45;
   wire north_input_control_N44;
   wire north_input_control_N43;
   wire north_input_control_N42;
   wire north_input_control_count_zero_f;
   wire north_input_control_header_last_f;
   wire north_input_control_count_one_f;
   wire north_input_control_tail_last_f;
   wire north_input_control_thanks_all_f;
   wire north_input_control_count_f_0_;
   wire north_input_control_count_f_1_;
   wire north_input_control_count_f_2_;
   wire north_input_control_count_f_3_;
   wire north_input_control_count_f_4_;
   wire north_input_control_count_f_5_;
   wire north_input_control_count_f_6_;
   wire north_input_control_count_f_7_;
   wire east_input_control_N53;
   wire east_input_control_N52;
   wire east_input_control_N51;
   wire east_input_control_N49;
   wire east_input_control_N48;
   wire east_input_control_N47;
   wire east_input_control_N46;
   wire east_input_control_N45;
   wire east_input_control_N44;
   wire east_input_control_N43;
   wire east_input_control_N42;
   wire east_input_control_N41;
   wire east_input_control_count_zero_f;
   wire east_input_control_header_last_f;
   wire east_input_control_count_one_f;
   wire east_input_control_tail_last_f;
   wire east_input_control_thanks_all_f;
   wire east_input_control_count_f_0_;
   wire east_input_control_count_f_1_;
   wire east_input_control_count_f_2_;
   wire east_input_control_count_f_3_;
   wire east_input_control_count_f_4_;
   wire east_input_control_count_f_5_;
   wire east_input_control_count_f_6_;
   wire east_input_control_count_f_7_;
   wire south_input_control_N53;
   wire south_input_control_N52;
   wire south_input_control_N51;
   wire south_input_control_N49;
   wire south_input_control_N48;
   wire south_input_control_N47;
   wire south_input_control_N46;
   wire south_input_control_N45;
   wire south_input_control_N44;
   wire south_input_control_N43;
   wire south_input_control_N42;
   wire south_input_control_count_zero_f;
   wire south_input_control_header_last_f;
   wire south_input_control_count_one_f;
   wire south_input_control_tail_last_f;
   wire south_input_control_thanks_all_f;
   wire south_input_control_count_f_0_;
   wire south_input_control_count_f_1_;
   wire south_input_control_count_f_2_;
   wire south_input_control_count_f_3_;
   wire south_input_control_count_f_4_;
   wire south_input_control_count_f_5_;
   wire south_input_control_count_f_6_;
   wire south_input_control_count_f_7_;
   wire west_input_control_N53;
   wire west_input_control_N52;
   wire west_input_control_N51;
   wire west_input_control_N49;
   wire west_input_control_N48;
   wire west_input_control_N47;
   wire west_input_control_N46;
   wire west_input_control_N45;
   wire west_input_control_N44;
   wire west_input_control_N43;
   wire west_input_control_N42;
   wire west_input_control_count_zero_f;
   wire west_input_control_header_last_f;
   wire west_input_control_count_one_f;
   wire west_input_control_tail_last_f;
   wire west_input_control_thanks_all_f;
   wire west_input_control_count_f_0_;
   wire west_input_control_count_f_1_;
   wire west_input_control_count_f_2_;
   wire west_input_control_count_f_3_;
   wire west_input_control_count_f_4_;
   wire west_input_control_count_f_5_;
   wire west_input_control_count_f_6_;
   wire west_input_control_count_f_7_;
   wire proc_input_control_N53;
   wire proc_input_control_N52;
   wire proc_input_control_N51;
   wire proc_input_control_N49;
   wire proc_input_control_N48;
   wire proc_input_control_N47;
   wire proc_input_control_N46;
   wire proc_input_control_N45;
   wire proc_input_control_N44;
   wire proc_input_control_N43;
   wire proc_input_control_N42;
   wire proc_input_control_N41;
   wire proc_input_control_count_zero_f;
   wire proc_input_control_header_last_f;
   wire proc_input_control_count_one_f;
   wire proc_input_control_tail_last_f;
   wire proc_input_control_thanks_all_f;
   wire proc_input_control_count_f_0_;
   wire proc_input_control_count_f_1_;
   wire proc_input_control_count_f_2_;
   wire proc_input_control_count_f_3_;
   wire proc_input_control_count_f_4_;
   wire proc_input_control_count_f_5_;
   wire proc_input_control_count_f_6_;
   wire proc_input_control_count_f_7_;
   wire north_output_current_route_connection_0_;
   wire north_output_current_route_connection_1_;
   wire north_output_current_route_connection_2_;
   wire east_output_current_route_connection_0_;
   wire east_output_current_route_connection_1_;
   wire east_output_current_route_connection_2_;
   wire south_output_current_route_connection_0_;
   wire south_output_current_route_connection_1_;
   wire south_output_current_route_connection_2_;
   wire west_output_current_route_connection_0_;
   wire west_output_current_route_connection_1_;
   wire west_output_current_route_connection_2_;
   wire proc_output_current_route_connection_0_;
   wire proc_output_current_route_connection_1_;
   wire proc_output_current_route_connection_2_;
   wire north_output_space_N48;
   wire north_output_space_N47;
   wire north_output_space_N46;
   wire north_output_space_N45;
   wire north_output_space_N44;
   wire north_output_space_N43;
   wire north_output_space_N42;
   wire north_output_space_valid_f;
   wire north_output_space_is_one_f;
   wire north_output_space_yummy_f;
   wire north_output_space_is_two_or_more_f;
   wire north_output_space_count_f_0_;
   wire north_output_space_count_f_1_;
   wire north_output_space_count_f_2_;
   wire east_output_space_N48;
   wire east_output_space_N47;
   wire east_output_space_N46;
   wire east_output_space_N45;
   wire east_output_space_N44;
   wire east_output_space_N43;
   wire east_output_space_N42;
   wire east_output_space_valid_f;
   wire east_output_space_is_one_f;
   wire east_output_space_yummy_f;
   wire east_output_space_is_two_or_more_f;
   wire east_output_space_count_f_0_;
   wire east_output_space_count_f_1_;
   wire east_output_space_count_f_2_;
   wire south_output_space_N48;
   wire south_output_space_N47;
   wire south_output_space_N46;
   wire south_output_space_N45;
   wire south_output_space_N44;
   wire south_output_space_N43;
   wire south_output_space_N42;
   wire south_output_space_valid_f;
   wire south_output_space_is_one_f;
   wire south_output_space_yummy_f;
   wire south_output_space_is_two_or_more_f;
   wire south_output_space_count_f_0_;
   wire south_output_space_count_f_1_;
   wire south_output_space_count_f_2_;
   wire west_output_space_N48;
   wire west_output_space_N47;
   wire west_output_space_N46;
   wire west_output_space_N45;
   wire west_output_space_N44;
   wire west_output_space_N43;
   wire west_output_space_N42;
   wire west_output_space_valid_f;
   wire west_output_space_is_one_f;
   wire west_output_space_yummy_f;
   wire west_output_space_is_two_or_more_f;
   wire west_output_space_count_f_0_;
   wire west_output_space_count_f_1_;
   wire west_output_space_count_f_2_;
   wire proc_output_space_N48;
   wire proc_output_space_N47;
   wire proc_output_space_N46;
   wire proc_output_space_N45;
   wire proc_output_space_N44;
   wire proc_output_space_N43;
   wire proc_output_space_N42;
   wire proc_output_space_valid_f;
   wire proc_output_space_is_one_f;
   wire proc_output_space_yummy_f;
   wire proc_output_space_is_two_or_more_f;
   wire proc_output_space_count_f_0_;
   wire proc_output_space_count_f_1_;
   wire proc_output_space_count_f_2_;
   wire north_output_control_N470;
   wire north_output_control_N469;
   wire north_output_control_N468;
   wire north_output_control_N467;
   wire north_output_control_N72;
   wire north_output_control_planned_f;
   wire east_output_control_N469;
   wire east_output_control_N468;
   wire east_output_control_N72;
   wire east_output_control_planned_f;
   wire south_output_control_N470;
   wire south_output_control_N469;
   wire south_output_control_N468;
   wire south_output_control_N467;
   wire south_output_control_N72;
   wire south_output_control_planned_f;
   wire west_output_control_N470;
   wire west_output_control_N469;
   wire west_output_control_N468;
   wire west_output_control_N467;
   wire west_output_control_N72;
   wire west_output_control_planned_f;
   wire proc_output_control_N470;
   wire proc_output_control_N469;
   wire proc_output_control_N468;
   wire proc_output_control_N467;
   wire proc_output_control_N72;
   wire proc_output_control_planned_f;
   wire n2418;
   wire n2423;
   wire n2433;
   wire n2438;
   wire n2443;
   wire n2558;
   wire n2563;
   wire n2573;
   wire n2578;
   wire n2583;
   wire n2688;
   wire n2693;
   wire n2703;
   wire n2833;
   wire n2838;
   wire n2843;
   wire n2848;
   wire n2853;
   wire n2858;
   wire n2863;
   wire n2868;
   wire n2873;
   wire n2988;
   wire n2993;
   wire n3003;
   wire n3093;
   wire n3098;
   wire n3103;
   wire n3108;
   wire n3113;
   wire n3118;
   wire n3123;
   wire n3128;
   wire n3133;
   wire n3138;
   wire n3143;
   wire n3148;
   wire n3153;
   wire n3158;
   wire n3163;
   wire n3168;
   wire n3173;
   wire n3178;
   wire n3183;
   wire n3188;
   wire n3193;
   wire n3198;
   wire n3203;
   wire n3208;
   wire n3213;
   wire n3218;
   wire n3223;
   wire n3228;
   wire n3233;
   wire n3238;
   wire n3243;
   wire n3248;
   wire n3253;
   wire n3258;
   wire n3263;
   wire n3268;
   wire n3273;
   wire n3278;
   wire n3283;
   wire n3288;
   wire n3293;
   wire n3298;
   wire n3303;
   wire n3308;
   wire n3313;
   wire n3318;
   wire n3323;
   wire n3328;
   wire n3333;
   wire n3338;
   wire n3343;
   wire n3348;
   wire n3353;
   wire n3358;
   wire n3363;
   wire n3368;
   wire n3373;
   wire n3378;
   wire n3383;
   wire n3388;
   wire n3393;
   wire n3398;
   wire n3403;
   wire n3408;
   wire n3413;
   wire n3418;
   wire n3423;
   wire n3428;
   wire n3433;
   wire n3438;
   wire n3443;
   wire n3448;
   wire n3453;
   wire n3458;
   wire n3463;
   wire n3468;
   wire n3473;
   wire n3478;
   wire n3483;
   wire n3488;
   wire n3493;
   wire n3498;
   wire n3503;
   wire n3508;
   wire n3513;
   wire n3518;
   wire n3523;
   wire n3528;
   wire n3533;
   wire n3538;
   wire n3543;
   wire n3548;
   wire n3553;
   wire n3558;
   wire n3563;
   wire n3568;
   wire n3573;
   wire n3578;
   wire n3583;
   wire n3588;
   wire n3593;
   wire n3598;
   wire n3603;
   wire n3608;
   wire n3613;
   wire n3618;
   wire n3623;
   wire n3628;
   wire n3633;
   wire n3638;
   wire n3643;
   wire n3648;
   wire n3653;
   wire n3658;
   wire n3663;
   wire n3668;
   wire n3673;
   wire n3678;
   wire n3683;
   wire n3688;
   wire n3693;
   wire n3698;
   wire n3703;
   wire n3708;
   wire n3713;
   wire n3718;
   wire n3723;
   wire n3728;
   wire n3733;
   wire n3738;
   wire n3743;
   wire n3748;
   wire n3753;
   wire n3758;
   wire n3763;
   wire n3768;
   wire n3773;
   wire n3778;
   wire n3783;
   wire n3788;
   wire n3793;
   wire n3798;
   wire n3803;
   wire n3808;
   wire n3813;
   wire n3818;
   wire n3823;
   wire n3828;
   wire n3833;
   wire n3838;
   wire n3843;
   wire n3848;
   wire n3853;
   wire n3858;
   wire n3863;
   wire n3868;
   wire n3873;
   wire n3878;
   wire n3883;
   wire n3888;
   wire n3893;
   wire n3898;
   wire n3903;
   wire n3908;
   wire n3913;
   wire n3918;
   wire n3923;
   wire n3928;
   wire n3933;
   wire n3938;
   wire n3943;
   wire n3948;
   wire n3953;
   wire n3958;
   wire n3963;
   wire n3968;
   wire n3973;
   wire n3978;
   wire n3983;
   wire n3988;
   wire n3993;
   wire n3998;
   wire n4003;
   wire n4008;
   wire n4013;
   wire n4018;
   wire n4023;
   wire n4028;
   wire n4033;
   wire n4038;
   wire n4043;
   wire n4048;
   wire n4053;
   wire n4058;
   wire n4063;
   wire n4068;
   wire n4073;
   wire n4078;
   wire n4083;
   wire n4088;
   wire n4093;
   wire n4098;
   wire n4103;
   wire n4108;
   wire n4113;
   wire n4118;
   wire n4123;
   wire n4128;
   wire n4133;
   wire n4138;
   wire n4143;
   wire n4148;
   wire n4153;
   wire n4158;
   wire n4163;
   wire n4168;
   wire n4173;
   wire n4178;
   wire n4183;
   wire n4188;
   wire n4193;
   wire n4198;
   wire n4203;
   wire n4208;
   wire n4213;
   wire n4218;
   wire n4223;
   wire n4228;
   wire n4233;
   wire n4238;
   wire n4243;
   wire n4248;
   wire n4253;
   wire n4258;
   wire n4263;
   wire n4268;
   wire n4273;
   wire n4278;
   wire n4283;
   wire n4288;
   wire n4293;
   wire n4298;
   wire n4303;
   wire n4308;
   wire n4313;
   wire n4318;
   wire n4323;
   wire n4328;
   wire n4333;
   wire n4338;
   wire n4343;
   wire n4348;
   wire n4353;
   wire n4358;
   wire n4363;
   wire n4368;
   wire n4373;
   wire n4378;
   wire n4383;
   wire n4388;
   wire n4393;
   wire n4398;
   wire n4403;
   wire n4408;
   wire n4413;
   wire n4418;
   wire n4423;
   wire n4428;
   wire n4433;
   wire n4438;
   wire n4443;
   wire n4448;
   wire n4453;
   wire n4458;
   wire n4463;
   wire n4468;
   wire n4473;
   wire n4478;
   wire n4483;
   wire n4488;
   wire n4493;
   wire n4498;
   wire n4503;
   wire n4508;
   wire n4513;
   wire n4518;
   wire n4523;
   wire n4528;
   wire n4533;
   wire n4538;
   wire n4543;
   wire n4548;
   wire n4553;
   wire n4558;
   wire n4563;
   wire n4568;
   wire n4573;
   wire n4578;
   wire n4583;
   wire n4588;
   wire n4593;
   wire n4598;
   wire n4603;
   wire n4608;
   wire n4613;
   wire n4618;
   wire n4623;
   wire n4628;
   wire n4633;
   wire n4638;
   wire n4643;
   wire n4648;
   wire n4653;
   wire n4658;
   wire n4663;
   wire n4668;
   wire n4673;
   wire n4678;
   wire n4683;
   wire n4688;
   wire n4693;
   wire n4698;
   wire n4703;
   wire n4708;
   wire n4713;
   wire n4718;
   wire n4723;
   wire n4728;
   wire n4733;
   wire n4738;
   wire n4743;
   wire n4748;
   wire n4753;
   wire n4758;
   wire n4763;
   wire n4768;
   wire n4773;
   wire n4778;
   wire n4783;
   wire n4788;
   wire n4793;
   wire n4798;
   wire n4803;
   wire n4808;
   wire n4813;
   wire n4818;
   wire n4823;
   wire n4828;
   wire n4833;
   wire n4838;
   wire n4843;
   wire n4848;
   wire n4853;
   wire n4858;
   wire n4863;
   wire n4868;
   wire n4873;
   wire n4878;
   wire n4883;
   wire n4888;
   wire n4893;
   wire n4898;
   wire n4903;
   wire n4908;
   wire n4913;
   wire n4918;
   wire n4923;
   wire n4928;
   wire n4933;
   wire n4938;
   wire n4943;
   wire n4948;
   wire n4953;
   wire n4958;
   wire n4963;
   wire n4968;
   wire n4973;
   wire n4978;
   wire n4983;
   wire n4988;
   wire n4993;
   wire n4998;
   wire n5003;
   wire n5008;
   wire n5013;
   wire n5018;
   wire n5023;
   wire n5028;
   wire n5033;
   wire n5038;
   wire n5043;
   wire n5048;
   wire n5053;
   wire n5058;
   wire n5063;
   wire n5068;
   wire n5073;
   wire n5078;
   wire n5083;
   wire n5088;
   wire n5093;
   wire n5098;
   wire n5103;
   wire n5108;
   wire n5113;
   wire n5118;
   wire n5123;
   wire n5128;
   wire n5133;
   wire n5138;
   wire n5143;
   wire n5148;
   wire n5153;
   wire n5158;
   wire n5163;
   wire n5168;
   wire n5173;
   wire n5178;
   wire n5183;
   wire n5188;
   wire n5193;
   wire n5198;
   wire n5203;
   wire n5208;
   wire n5213;
   wire n5218;
   wire n5223;
   wire n5228;
   wire n5233;
   wire n5238;
   wire n5243;
   wire n5248;
   wire n5253;
   wire n5258;
   wire n5263;
   wire n5268;
   wire n5273;
   wire n5278;
   wire n5283;
   wire n5288;
   wire n5293;
   wire n5298;
   wire n5303;
   wire n5308;
   wire n5313;
   wire n5318;
   wire n5323;
   wire n5328;
   wire n5333;
   wire n5338;
   wire n5343;
   wire n5348;
   wire n5353;
   wire n5358;
   wire n5363;
   wire n5368;
   wire n5373;
   wire n5378;
   wire n5383;
   wire n5388;
   wire n5393;
   wire n5398;
   wire n5403;
   wire n5408;
   wire n5413;
   wire n5418;
   wire n5423;
   wire n5428;
   wire n5433;
   wire n5438;
   wire n5443;
   wire n5448;
   wire n5453;
   wire n5458;
   wire n5463;
   wire n5468;
   wire n5473;
   wire n5478;
   wire n5483;
   wire n5488;
   wire n5493;
   wire n5498;
   wire n5503;
   wire n5508;
   wire n5513;
   wire n5518;
   wire n5523;
   wire n5528;
   wire n5533;
   wire n5538;
   wire n5543;
   wire n5548;
   wire n5553;
   wire n5558;
   wire n5563;
   wire n5568;
   wire n5573;
   wire n5578;
   wire n5583;
   wire n5588;
   wire n5593;
   wire n5598;
   wire n5603;
   wire n5608;
   wire n5613;
   wire n5618;
   wire n5623;
   wire n5628;
   wire n5633;
   wire n5638;
   wire n5643;
   wire n5648;
   wire n5653;
   wire n5658;
   wire n5663;
   wire n5668;
   wire n5673;
   wire n5678;
   wire n5683;
   wire n5688;
   wire n5693;
   wire n5698;
   wire n5703;
   wire n5708;
   wire n5713;
   wire n5718;
   wire n5723;
   wire n5728;
   wire n5733;
   wire n5738;
   wire n5743;
   wire n5748;
   wire n5753;
   wire n5758;
   wire n5763;
   wire n5768;
   wire n5773;
   wire n5778;
   wire n5783;
   wire n5788;
   wire n5793;
   wire n5798;
   wire n5803;
   wire n5808;
   wire n5813;
   wire n5818;
   wire n5823;
   wire n5828;
   wire n5833;
   wire n5838;
   wire n5843;
   wire n5848;
   wire n5853;
   wire n5858;
   wire n5863;
   wire n5868;
   wire n5873;
   wire n5878;
   wire n5883;
   wire n5888;
   wire n5893;
   wire n5898;
   wire n5903;
   wire n5908;
   wire n5913;
   wire n5918;
   wire n5923;
   wire n5928;
   wire n5933;
   wire n5938;
   wire n5943;
   wire n5948;
   wire n5953;
   wire n5958;
   wire n5963;
   wire n5968;
   wire n5973;
   wire n5978;
   wire n5983;
   wire n5988;
   wire n5993;
   wire n5998;
   wire n6003;
   wire n6008;
   wire n6013;
   wire n6018;
   wire n6023;
   wire n6028;
   wire n6033;
   wire n6038;
   wire n6043;
   wire n6048;
   wire n6053;
   wire n6058;
   wire n6063;
   wire n6068;
   wire n6073;
   wire n6078;
   wire n6083;
   wire n6088;
   wire n6093;
   wire n6098;
   wire n6103;
   wire n6108;
   wire n6113;
   wire n6118;
   wire n6123;
   wire n6128;
   wire n6133;
   wire n6138;
   wire n6143;
   wire n6148;
   wire n6153;
   wire n6158;
   wire n6163;
   wire n6168;
   wire n6173;
   wire n6178;
   wire n6183;
   wire n6188;
   wire n6193;
   wire n6198;
   wire n6203;
   wire n6208;
   wire n6213;
   wire n6218;
   wire n6223;
   wire n6228;
   wire n6233;
   wire n6238;
   wire n6243;
   wire n6248;
   wire n6253;
   wire n6258;
   wire n6263;
   wire n6268;
   wire n6273;
   wire n6278;
   wire n6283;
   wire n6288;
   wire n6293;
   wire n6298;
   wire n6303;
   wire n6308;
   wire n6313;
   wire n6318;
   wire n6323;
   wire n6328;
   wire n6333;
   wire n6338;
   wire n6343;
   wire n6348;
   wire n6353;
   wire n6358;
   wire n6363;
   wire n6368;
   wire n6373;
   wire n6378;
   wire n6383;
   wire n6388;
   wire n6393;
   wire n6398;
   wire n6403;
   wire n6408;
   wire n6413;
   wire n6418;
   wire n6423;
   wire n6428;
   wire n6433;
   wire n6438;
   wire n6443;
   wire n6448;
   wire n6453;
   wire n6458;
   wire n6463;
   wire n6468;
   wire n6473;
   wire n6478;
   wire n6483;
   wire n6488;
   wire n6493;
   wire n6498;
   wire n6503;
   wire n6508;
   wire n6513;
   wire n6518;
   wire n6523;
   wire n6528;
   wire n6533;
   wire n6538;
   wire n6543;
   wire n6548;
   wire n6553;
   wire n6558;
   wire n6563;
   wire n6568;
   wire n6573;
   wire n6578;
   wire n6583;
   wire n6588;
   wire n6593;
   wire n6598;
   wire n6603;
   wire n6608;
   wire n6613;
   wire n6618;
   wire n6623;
   wire n6628;
   wire n6633;
   wire n6638;
   wire n6643;
   wire n6648;
   wire n6653;
   wire n6658;
   wire n6663;
   wire n6668;
   wire n6673;
   wire n6678;
   wire n6683;
   wire n6688;
   wire n6693;
   wire n6698;
   wire n6703;
   wire n6708;
   wire n6713;
   wire n6718;
   wire n6723;
   wire n6728;
   wire n6733;
   wire n6738;
   wire n6743;
   wire n6748;
   wire n6753;
   wire n6758;
   wire n6763;
   wire n6768;
   wire n6773;
   wire n6778;
   wire n6783;
   wire n6788;
   wire n6793;
   wire n6798;
   wire n6803;
   wire n6808;
   wire n6813;
   wire n6818;
   wire n6823;
   wire n6828;
   wire n6833;
   wire n6838;
   wire n6843;
   wire n6848;
   wire n6853;
   wire n6858;
   wire n6863;
   wire n6868;
   wire n6873;
   wire n6878;
   wire n6883;
   wire n6888;
   wire n6893;
   wire n6898;
   wire n6903;
   wire n6908;
   wire n6913;
   wire n6918;
   wire n6923;
   wire n6928;
   wire n6933;
   wire n6938;
   wire n6943;
   wire n6948;
   wire n6953;
   wire n6958;
   wire n6963;
   wire n6968;
   wire n6973;
   wire n6978;
   wire n6983;
   wire n6988;
   wire n6993;
   wire n6998;
   wire n7003;
   wire n7008;
   wire n7013;
   wire n7018;
   wire n7023;
   wire n7028;
   wire n7033;
   wire n7038;
   wire n7043;
   wire n7048;
   wire n7053;
   wire n7058;
   wire n7063;
   wire n7068;
   wire n7073;
   wire n7078;
   wire n7083;
   wire n7088;
   wire n7093;
   wire n7098;
   wire n7103;
   wire n7108;
   wire n7113;
   wire n7118;
   wire n7123;
   wire n7128;
   wire n7133;
   wire n7138;
   wire n7143;
   wire n7148;
   wire n7153;
   wire n7158;
   wire n7163;
   wire n7168;
   wire n7173;
   wire n7178;
   wire n7183;
   wire n7188;
   wire n7193;
   wire n7198;
   wire n7203;
   wire n7208;
   wire n7213;
   wire n7218;
   wire n7223;
   wire n7228;
   wire n7233;
   wire n7238;
   wire n7243;
   wire n7248;
   wire n7253;
   wire n7258;
   wire n7263;
   wire n7268;
   wire n7273;
   wire n7278;
   wire n7283;
   wire n7288;
   wire n7293;
   wire n7298;
   wire n7303;
   wire n7308;
   wire n7313;
   wire n7318;
   wire n7323;
   wire n7328;
   wire n7333;
   wire n7338;
   wire n7343;
   wire n7348;
   wire n7353;
   wire n7358;
   wire n7363;
   wire n7368;
   wire n7373;
   wire n7378;
   wire n7383;
   wire n7388;
   wire n7393;
   wire n7398;
   wire n7403;
   wire n7408;
   wire n7413;
   wire n7418;
   wire n7423;
   wire n7428;
   wire n7433;
   wire n7438;
   wire n7443;
   wire n7448;
   wire n7453;
   wire n7458;
   wire n7463;
   wire n7468;
   wire n7473;
   wire n7478;
   wire n7483;
   wire n7488;
   wire n7493;
   wire n7498;
   wire n7503;
   wire n7508;
   wire n7513;
   wire n7518;
   wire n7523;
   wire n7528;
   wire n7533;
   wire n7538;
   wire n7543;
   wire n7548;
   wire n7553;
   wire n7558;
   wire n7563;
   wire n7568;
   wire n7573;
   wire n7578;
   wire n7583;
   wire n7588;
   wire n7593;
   wire n7598;
   wire n7603;
   wire n7608;
   wire n7613;
   wire n7618;
   wire n7623;
   wire n7628;
   wire n7633;
   wire n7638;
   wire n7643;
   wire n7648;
   wire n7653;
   wire n7658;
   wire n7663;
   wire n7668;
   wire n7673;
   wire n7678;
   wire n7683;
   wire n7688;
   wire n7693;
   wire n7698;
   wire n7703;
   wire n7708;
   wire n7713;
   wire n7718;
   wire n7723;
   wire n7728;
   wire n7733;
   wire n7738;
   wire n7743;
   wire n7748;
   wire n7753;
   wire n7758;
   wire n7763;
   wire n7768;
   wire n7773;
   wire n7778;
   wire n7783;
   wire n7788;
   wire n7793;
   wire n7798;
   wire n7803;
   wire n7808;
   wire n7813;
   wire n7818;
   wire n7823;
   wire n7828;
   wire n7833;
   wire n7838;
   wire n7843;
   wire n7848;
   wire n7853;
   wire n7858;
   wire n7863;
   wire n7868;
   wire n7873;
   wire n7878;
   wire n7883;
   wire n7888;
   wire n7893;
   wire n7898;
   wire n7903;
   wire n7908;
   wire n7913;
   wire n7918;
   wire n7923;
   wire n7928;
   wire n7933;
   wire n7938;
   wire n7943;
   wire n7948;
   wire n7953;
   wire n7958;
   wire n7963;
   wire n7968;
   wire n7973;
   wire n7978;
   wire n7983;
   wire n7988;
   wire n7993;
   wire n7998;
   wire n8003;
   wire n8008;
   wire n8013;
   wire n8018;
   wire n8023;
   wire n8028;
   wire n8033;
   wire n8038;
   wire n8043;
   wire n8048;
   wire n8053;
   wire n8058;
   wire n8063;
   wire n8068;
   wire n8073;
   wire n8078;
   wire n8083;
   wire n8088;
   wire n8093;
   wire n8098;
   wire n8103;
   wire n8108;
   wire n8113;
   wire n8118;
   wire n8123;
   wire n8128;
   wire n8133;
   wire n8138;
   wire n8143;
   wire n8148;
   wire n8153;
   wire n8158;
   wire n8163;
   wire n8168;
   wire n8173;
   wire n8178;
   wire n8183;
   wire n8188;
   wire n8193;
   wire n8198;
   wire n8203;
   wire n8208;
   wire n8213;
   wire n8218;
   wire n8223;
   wire n8228;
   wire n8233;
   wire n8238;
   wire n8243;
   wire n8248;
   wire n8253;
   wire n8258;
   wire n8263;
   wire n8268;
   wire n8273;
   wire n8278;
   wire n8283;
   wire n8288;
   wire n8293;
   wire n8298;
   wire n8303;
   wire n8308;
   wire n8313;
   wire n8318;
   wire n8323;
   wire n8328;
   wire n8333;
   wire n8338;
   wire n8343;
   wire n8348;
   wire n8353;
   wire n8358;
   wire n8363;
   wire n8368;
   wire n8373;
   wire n8378;
   wire n8383;
   wire n8388;
   wire n8393;
   wire n8398;
   wire n8403;
   wire n8408;
   wire n8413;
   wire n8418;
   wire n8423;
   wire n8428;
   wire n8433;
   wire n8438;
   wire n8443;
   wire n8448;
   wire n8453;
   wire n8458;
   wire n8463;
   wire n8468;
   wire n8473;
   wire n8478;
   wire n8483;
   wire n8488;
   wire n8493;
   wire n8498;
   wire n8503;
   wire n8508;
   wire n8513;
   wire n8518;
   wire n8523;
   wire n8528;
   wire n8533;
   wire n8538;
   wire n8543;
   wire n8548;
   wire n8553;
   wire n8558;
   wire n8563;
   wire n8568;
   wire n8573;
   wire n8578;
   wire n8583;
   wire n8588;
   wire n8593;
   wire n8598;
   wire n8603;
   wire n8608;
   wire n8613;
   wire n8618;
   wire n8623;
   wire n8628;
   wire n8633;
   wire n8638;
   wire n8643;
   wire n8648;
   wire n8653;
   wire n8658;
   wire n8663;
   wire n8668;
   wire n8673;
   wire n8678;
   wire n8683;
   wire n8688;
   wire n8693;
   wire n8698;
   wire n8703;
   wire n8708;
   wire n8713;
   wire n8718;
   wire n8723;
   wire n8728;
   wire n8733;
   wire n8738;
   wire n8743;
   wire n8748;
   wire n8753;
   wire n8758;
   wire n8763;
   wire n8768;
   wire n8773;
   wire n8778;
   wire n8783;
   wire n8788;
   wire n8793;
   wire n8798;
   wire n8803;
   wire n8808;
   wire n8813;
   wire n8818;
   wire n8823;
   wire n8828;
   wire n8833;
   wire n8838;
   wire n8843;
   wire n8848;
   wire n8853;
   wire n8858;
   wire n8863;
   wire n8868;
   wire n8873;
   wire n8878;
   wire n8883;
   wire n8888;
   wire n8893;
   wire n8898;
   wire n8903;
   wire n8908;
   wire n8913;
   wire n8918;
   wire n8923;
   wire n8928;
   wire n8933;
   wire n8938;
   wire n8943;
   wire n8948;
   wire n8953;
   wire n8958;
   wire n8963;
   wire n8968;
   wire n8973;
   wire n8978;
   wire n8983;
   wire n8988;
   wire n8993;
   wire n8998;
   wire n9003;
   wire n9008;
   wire n9013;
   wire n9018;
   wire n9023;
   wire n9028;
   wire n9033;
   wire n9038;
   wire n9043;
   wire n9048;
   wire n9053;
   wire n9058;
   wire n9063;
   wire n9068;
   wire n9073;
   wire n9078;
   wire n9083;
   wire n9088;
   wire n9093;
   wire n9098;
   wire n9103;
   wire n9108;
   wire n9113;
   wire n9118;
   wire n9123;
   wire n9128;
   wire n9133;
   wire n9138;
   wire n9143;
   wire n9148;
   wire n9153;
   wire n9158;
   wire n9163;
   wire n9168;
   wire n9173;
   wire n9178;
   wire n9183;
   wire n9188;
   wire n9193;
   wire n9198;
   wire n9203;
   wire n9208;
   wire n9213;
   wire n9218;
   wire n9223;
   wire n9228;
   wire n9233;
   wire n9238;
   wire n9243;
   wire n9248;
   wire n9253;
   wire n9258;
   wire n9263;
   wire n9268;
   wire n9273;
   wire n9278;
   wire n9283;
   wire n9288;
   wire n9293;
   wire n9298;
   wire n9303;
   wire n9308;
   wire n9313;
   wire n9318;
   wire n9323;
   wire n9328;
   wire n9333;
   wire n9338;
   wire n9343;
   wire n9348;
   wire n9353;
   wire n9358;
   wire n9363;
   wire n9368;
   wire n9373;
   wire n9378;
   wire n9383;
   wire n9388;
   wire n9393;
   wire n9398;
   wire n9403;
   wire n9408;
   wire n9413;
   wire n9418;
   wire n9423;
   wire n9428;
   wire n9433;
   wire n9438;
   wire n9443;
   wire n9448;
   wire n9453;
   wire n9458;
   wire n9463;
   wire n9468;
   wire n9473;
   wire n9478;
   wire n9483;
   wire n9488;
   wire n9493;
   wire n9498;
   wire n9503;
   wire n9508;
   wire n9513;
   wire n9518;
   wire n9523;
   wire n9528;
   wire n9533;
   wire n9538;
   wire n9543;
   wire n9548;
   wire n9553;
   wire n9558;
   wire n9563;
   wire n9568;
   wire n9573;
   wire n9578;
   wire n9583;
   wire n9588;
   wire n9593;
   wire n9598;
   wire n9603;
   wire n9608;
   wire n9613;
   wire n9618;
   wire n9623;
   wire n9628;
   wire n9633;
   wire n9638;
   wire n9643;
   wire n9648;
   wire n9653;
   wire n9658;
   wire n9663;
   wire n9668;
   wire n9673;
   wire n9678;
   wire n9683;
   wire n9688;
   wire n9693;
   wire n9698;
   wire n9703;
   wire n9708;
   wire n9713;
   wire n9718;
   wire n9723;
   wire n9728;
   wire n9733;
   wire n9738;
   wire n9743;
   wire n9748;
   wire n9753;
   wire n9758;
   wire n9763;
   wire n9768;
   wire n9773;
   wire n9778;
   wire n9783;
   wire n9788;
   wire n9793;
   wire n9798;
   wire n9803;
   wire n9808;
   wire n9813;
   wire n9818;
   wire n9823;
   wire n9828;
   wire n9833;
   wire n9838;
   wire n9843;
   wire n9848;
   wire n9853;
   wire n9858;
   wire n9863;
   wire n9868;
   wire n9873;
   wire n9878;
   wire n9883;
   wire n9888;
   wire n9893;
   wire n9898;
   wire n9903;
   wire n9908;
   wire n9913;
   wire n9918;
   wire n9923;
   wire n9928;
   wire n9933;
   wire n9938;
   wire n9943;
   wire n9948;
   wire n9953;
   wire n9958;
   wire n9963;
   wire n9968;
   wire n9973;
   wire n9978;
   wire n9983;
   wire n9988;
   wire n9993;
   wire n9998;
   wire n10003;
   wire n10008;
   wire n10013;
   wire n10018;
   wire n10023;
   wire n10028;
   wire n10033;
   wire n10038;
   wire n10043;
   wire n10048;
   wire n10053;
   wire n10058;
   wire n10063;
   wire n10068;
   wire n10073;
   wire n10078;
   wire n10083;
   wire n10088;
   wire n10093;
   wire n10098;
   wire n10103;
   wire n10108;
   wire n10113;
   wire n10118;
   wire n10123;
   wire n10128;
   wire n10133;
   wire n10138;
   wire n10143;
   wire n10148;
   wire n10153;
   wire n10158;
   wire n10163;
   wire n10168;
   wire n10173;
   wire n10178;
   wire n10183;
   wire n10188;
   wire n10193;
   wire n10198;
   wire n10203;
   wire n10208;
   wire n10213;
   wire n10218;
   wire n10223;
   wire n10228;
   wire n10233;
   wire n10238;
   wire n10243;
   wire n10248;
   wire n10253;
   wire n10258;
   wire n10263;
   wire n10268;
   wire n10273;
   wire n10278;
   wire n10283;
   wire n10288;
   wire n10293;
   wire n10298;
   wire n10303;
   wire n10308;
   wire n10313;
   wire n10318;
   wire n10323;
   wire n10328;
   wire n10333;
   wire n10338;
   wire n10343;
   wire n10348;
   wire n10353;
   wire n10358;
   wire n10363;
   wire n10368;
   wire n10373;
   wire n10378;
   wire n10383;
   wire n10388;
   wire n10393;
   wire n10398;
   wire n10403;
   wire n10408;
   wire n10413;
   wire n10418;
   wire n10423;
   wire n10428;
   wire n10433;
   wire n10438;
   wire n10443;
   wire n10448;
   wire n10453;
   wire n10458;
   wire n10463;
   wire n10468;
   wire n10473;
   wire n10478;
   wire n10483;
   wire n10488;
   wire n10493;
   wire n10498;
   wire n10503;
   wire n10508;
   wire n10513;
   wire n10518;
   wire n10523;
   wire n10528;
   wire n10533;
   wire n10538;
   wire n10543;
   wire n10548;
   wire n10553;
   wire n10558;
   wire n10563;
   wire n10568;
   wire n10573;
   wire n10578;
   wire n10583;
   wire n10588;
   wire n10593;
   wire n10598;
   wire n10603;
   wire n10608;
   wire n10613;
   wire n10618;
   wire n10623;
   wire n10628;
   wire n10633;
   wire n10638;
   wire n10643;
   wire n10648;
   wire n10653;
   wire n10658;
   wire n10663;
   wire n10668;
   wire n10673;
   wire n10678;
   wire n10683;
   wire n10688;
   wire n10693;
   wire n10698;
   wire n10703;
   wire n10708;
   wire n10713;
   wire n10718;
   wire n10723;
   wire n10728;
   wire n10733;
   wire n10738;
   wire n10743;
   wire n10748;
   wire n10753;
   wire n10758;
   wire n10763;
   wire n10768;
   wire n10773;
   wire n10778;
   wire n10783;
   wire n10788;
   wire n10793;
   wire n10798;
   wire n10803;
   wire n10808;
   wire n10813;
   wire n10818;
   wire n10823;
   wire n10828;
   wire n10833;
   wire n10838;
   wire n10843;
   wire n10848;
   wire n10853;
   wire n10858;
   wire n10863;
   wire n10868;
   wire n10873;
   wire n10878;
   wire n10883;
   wire n10888;
   wire n10893;
   wire n10898;
   wire n10903;
   wire n10908;
   wire n10913;
   wire n10918;
   wire n10923;
   wire n10928;
   wire n10933;
   wire n10938;
   wire n10943;
   wire n10948;
   wire n10953;
   wire n10958;
   wire n10963;
   wire n10968;
   wire n10973;
   wire n10978;
   wire n10983;
   wire n10988;
   wire n10993;
   wire n10998;
   wire n11003;
   wire n11008;
   wire n11013;
   wire n11018;
   wire n11023;
   wire n11028;
   wire n11033;
   wire n11038;
   wire n11043;
   wire n11048;
   wire n11053;
   wire n11058;
   wire n11063;
   wire n11068;
   wire n11073;
   wire n11078;
   wire n11083;
   wire n11088;
   wire n11093;
   wire n11098;
   wire n11103;
   wire n11108;
   wire n11113;
   wire n11118;
   wire n11123;
   wire n11128;
   wire n11133;
   wire n11138;
   wire n11143;
   wire n11148;
   wire n11153;
   wire n11158;
   wire n11163;
   wire n11168;
   wire n11173;
   wire n11178;
   wire n11183;
   wire n11188;
   wire n11193;
   wire n11198;
   wire n11203;
   wire n11208;
   wire n11213;
   wire n11218;
   wire n11223;
   wire n11228;
   wire n11233;
   wire n11238;
   wire n11243;
   wire n11248;
   wire n11253;
   wire n11258;
   wire n11263;
   wire n11268;
   wire n11273;
   wire n11278;
   wire n11283;
   wire n11288;
   wire n11293;
   wire n11298;
   wire n11303;
   wire n11308;
   wire n11313;
   wire n11318;
   wire n11323;
   wire n11328;
   wire n11333;
   wire n11338;
   wire n11343;
   wire n11348;
   wire n11353;
   wire n11358;
   wire n11363;
   wire n11368;
   wire n11373;
   wire n11378;
   wire n11383;
   wire n11388;
   wire n11393;
   wire n11398;
   wire n11403;
   wire n11408;
   wire n11413;
   wire n11418;
   wire n11423;
   wire n11428;
   wire n11433;
   wire n11438;
   wire n11443;
   wire n11448;
   wire n11453;
   wire n11458;
   wire n11463;
   wire n11468;
   wire n11473;
   wire n11478;
   wire n11483;
   wire n11488;
   wire n11493;
   wire n11498;
   wire n11503;
   wire n11508;
   wire n11513;
   wire n11518;
   wire n11523;
   wire n11528;
   wire n11533;
   wire n11538;
   wire n11543;
   wire n11548;
   wire n11553;
   wire n11558;
   wire n11563;
   wire n11568;
   wire n11573;
   wire n11578;
   wire n11583;
   wire n11588;
   wire n11593;
   wire n11598;
   wire n11603;
   wire n11608;
   wire n11613;
   wire n11618;
   wire n11623;
   wire n11628;
   wire n11633;
   wire n11638;
   wire n11643;
   wire n11648;
   wire n11653;
   wire n11658;
   wire n11663;
   wire n11668;
   wire n11673;
   wire n11678;
   wire n11683;
   wire n11688;
   wire n11693;
   wire n11698;
   wire n11703;
   wire n11708;
   wire n11713;
   wire n11718;
   wire n11723;
   wire n11728;
   wire n11733;
   wire n11738;
   wire n11743;
   wire n11748;
   wire n11753;
   wire n11758;
   wire n11763;
   wire n11768;
   wire n11773;
   wire n11778;
   wire n11783;
   wire n11788;
   wire n11793;
   wire n11798;
   wire n11803;
   wire n11808;
   wire n11813;
   wire n11818;
   wire n11823;
   wire n11828;
   wire n11833;
   wire n11838;
   wire n11843;
   wire n11848;
   wire n11853;
   wire n11858;
   wire n11863;
   wire n11868;
   wire n11873;
   wire n11878;
   wire n11883;
   wire n11888;
   wire n11893;
   wire n11898;
   wire n11903;
   wire n11908;
   wire n11913;
   wire n11918;
   wire n11923;
   wire n11928;
   wire n11933;
   wire n11938;
   wire n11943;
   wire n11948;
   wire n11953;
   wire n11958;
   wire n11963;
   wire n11968;
   wire n11973;
   wire n11978;
   wire n11983;
   wire n11988;
   wire n11993;
   wire n11998;
   wire n12003;
   wire n12008;
   wire n12013;
   wire n12018;
   wire n12023;
   wire n12028;
   wire n12033;
   wire n12038;
   wire n12043;
   wire n12048;
   wire n12053;
   wire n12058;
   wire n12063;
   wire n12068;
   wire n12073;
   wire n12078;
   wire n12083;
   wire n12088;
   wire n12093;
   wire n12098;
   wire n12103;
   wire n12108;
   wire n12113;
   wire n12118;
   wire n12123;
   wire n12128;
   wire n12133;
   wire n12138;
   wire n12143;
   wire n12148;
   wire n12153;
   wire n12158;
   wire n12163;
   wire n12168;
   wire n12173;
   wire n12178;
   wire n12183;
   wire n12188;
   wire n12193;
   wire n12198;
   wire n12203;
   wire n12208;
   wire n12213;
   wire n12218;
   wire n12223;
   wire n12228;
   wire n12233;
   wire n12238;
   wire n12243;
   wire n12248;
   wire n12253;
   wire n12258;
   wire n12263;
   wire n12268;
   wire n12273;
   wire n12278;
   wire n12283;
   wire n12288;
   wire n12293;
   wire n12298;
   wire n12303;
   wire n12308;
   wire n12313;
   wire n12318;
   wire n12323;
   wire n12328;
   wire n12333;
   wire n12338;
   wire n12343;
   wire n12348;
   wire n12353;
   wire n12358;
   wire n12363;
   wire n12368;
   wire n12373;
   wire n12378;
   wire n12383;
   wire n12388;
   wire n12393;
   wire n12398;
   wire n12403;
   wire n12408;
   wire n12413;
   wire n12418;
   wire n12423;
   wire n12428;
   wire n12433;
   wire n12438;
   wire n12443;
   wire n12448;
   wire n12453;
   wire n12458;
   wire n12463;
   wire n12468;
   wire n12473;
   wire n12478;
   wire n12483;
   wire n12488;
   wire n12493;
   wire n12498;
   wire n12503;
   wire n12508;
   wire n12513;
   wire n12518;
   wire n12523;
   wire n12528;
   wire n12533;
   wire n12538;
   wire n12543;
   wire n12548;
   wire n12553;
   wire n12558;
   wire n12563;
   wire n12568;
   wire n12573;
   wire n12578;
   wire n12583;
   wire n12588;
   wire n12593;
   wire n12598;
   wire n12603;
   wire n12608;
   wire n12613;
   wire n12618;
   wire n12623;
   wire n12628;
   wire n12633;
   wire n12638;
   wire n12643;
   wire n12648;
   wire n12653;
   wire n12658;
   wire n12663;
   wire n12668;
   wire n12673;
   wire n12678;
   wire n12683;
   wire n12688;
   wire n12693;
   wire n12698;
   wire n12703;
   wire n12708;
   wire n12713;
   wire n12718;
   wire n12723;
   wire n12728;
   wire n12733;
   wire n12738;
   wire n12743;
   wire n12748;
   wire n12753;
   wire n12758;
   wire n12763;
   wire n12768;
   wire n12773;
   wire n12778;
   wire n12783;
   wire n12788;
   wire n12793;
   wire n12798;
   wire n12803;
   wire n12808;
   wire n12813;
   wire n12818;
   wire n12823;
   wire n12828;
   wire n12833;
   wire n12838;
   wire n12843;
   wire n12848;
   wire n12853;
   wire n12858;
   wire n12863;
   wire n12868;
   wire n12873;
   wire n12878;
   wire n12883;
   wire n12888;
   wire n12893;
   wire n12898;
   wire n12903;
   wire n12908;
   wire n12913;
   wire n12918;
   wire n12923;
   wire n12928;
   wire n12933;
   wire n12938;
   wire n12943;
   wire n12948;
   wire n12953;
   wire n12958;
   wire n12963;
   wire n12968;
   wire n12973;
   wire n12978;
   wire n12983;
   wire n12988;
   wire n12993;
   wire n12998;
   wire n13003;
   wire n13008;
   wire n13013;
   wire n13018;
   wire n13023;
   wire n13028;
   wire n13033;
   wire n13038;
   wire n13043;
   wire n13048;
   wire n13053;
   wire n13058;
   wire n13063;
   wire n13068;
   wire n13073;
   wire n13078;
   wire n13083;
   wire n13088;
   wire n13093;
   wire n13098;
   wire n13103;
   wire n13108;
   wire n13113;
   wire n13118;
   wire n13123;
   wire n13128;
   wire n13133;
   wire n13138;
   wire n13143;
   wire n13148;
   wire n13153;
   wire n13158;
   wire n13163;
   wire n13168;
   wire n13173;
   wire n13178;
   wire n13183;
   wire n13188;
   wire n13193;
   wire n13198;
   wire n13203;
   wire n13208;
   wire n13213;
   wire n13218;
   wire n13223;
   wire n13228;
   wire n13233;
   wire n13238;
   wire n13243;
   wire n13248;
   wire n13253;
   wire n13258;
   wire n13263;
   wire n13268;
   wire n13273;
   wire n13278;
   wire n13283;
   wire n13288;
   wire n13293;
   wire n13298;
   wire n13303;
   wire n13308;
   wire n13313;
   wire n13318;
   wire n13323;
   wire n13328;
   wire n13333;
   wire n13338;
   wire n13343;
   wire n13348;
   wire n13353;
   wire n13358;
   wire n13363;
   wire n13368;
   wire n13373;
   wire n13378;
   wire n13383;
   wire n13388;
   wire n17736;
   wire n17737;
   wire n17738;
   wire n17739;
   wire n17740;
   wire n17741;
   wire n17742;
   wire n17743;
   wire n17744;
   wire n17747;
   wire n17749;
   wire n17751;
   wire n17753;
   wire n17754;
   wire n17755;
   wire n17756;
   wire n17757;
   wire n17758;
   wire n17759;
   wire n17760;
   wire n17761;
   wire n17762;
   wire n17763;
   wire n17764;
   wire n17765;
   wire n17766;
   wire n17767;
   wire n17768;
   wire n17769;
   wire n17770;
   wire n17771;
   wire n17772;
   wire n17773;
   wire n17774;
   wire n17777;
   wire n17779;
   wire n17780;
   wire n17782;
   wire n17783;
   wire n17784;
   wire n17785;
   wire n17786;
   wire n17787;
   wire n17788;
   wire n17789;
   wire n17792;
   wire n17793;
   wire n17794;
   wire n17795;
   wire n17796;
   wire n17797;
   wire n17798;
   wire n17799;
   wire n17800;
   wire n17801;
   wire n17802;
   wire n17803;
   wire n17804;
   wire n17805;
   wire n17806;
   wire n17807;
   wire n17808;
   wire n17809;
   wire n17810;
   wire n17811;
   wire n17812;
   wire n17813;
   wire n17814;
   wire n17815;
   wire n17816;
   wire n17817;
   wire n17818;
   wire n17819;
   wire n17820;
   wire n17821;
   wire n17822;
   wire n17823;
   wire n17824;
   wire n17825;
   wire n17826;
   wire n17827;
   wire n17828;
   wire n17829;
   wire n17830;
   wire n17831;
   wire n17832;
   wire n17833;
   wire n17834;
   wire n17835;
   wire n17836;
   wire n17837;
   wire n17838;
   wire n17839;
   wire n17840;
   wire n17841;
   wire n17842;
   wire n17843;
   wire n17844;
   wire n17845;
   wire n17846;
   wire n17847;
   wire n17848;
   wire n17849;
   wire n17850;
   wire n17851;
   wire n17852;
   wire n17853;
   wire n17854;
   wire n17855;
   wire n17856;
   wire n17857;
   wire n17858;
   wire n17859;
   wire n17860;
   wire n17861;
   wire n17862;
   wire n17863;
   wire n17864;
   wire n17865;
   wire n17866;
   wire n17867;
   wire n17868;
   wire n17869;
   wire n17870;
   wire n17871;
   wire n17872;
   wire n17873;
   wire n17874;
   wire n17875;
   wire n17876;
   wire n17877;
   wire n17878;
   wire n17879;
   wire n17880;
   wire n17881;
   wire n17882;
   wire n17883;
   wire n17884;
   wire n17885;
   wire n17886;
   wire n17887;
   wire n17888;
   wire n17889;
   wire n17890;
   wire n17891;
   wire n17892;
   wire n17893;
   wire n17894;
   wire n17895;
   wire n17896;
   wire n17897;
   wire n17898;
   wire n17899;
   wire n17900;
   wire n17901;
   wire n17902;
   wire n17903;
   wire n17904;
   wire n17905;
   wire n17906;
   wire n17907;
   wire n17908;
   wire n17909;
   wire n17910;
   wire n17911;
   wire n17912;
   wire n17913;
   wire n17914;
   wire n17915;
   wire n17916;
   wire n17917;
   wire n17918;
   wire n17919;
   wire n17920;
   wire n17921;
   wire n17922;
   wire n17923;
   wire n17924;
   wire n17925;
   wire n17926;
   wire n17927;
   wire n17928;
   wire n17929;
   wire n17930;
   wire n17931;
   wire n17932;
   wire n17933;
   wire n17934;
   wire n17935;
   wire n17936;
   wire n17937;
   wire n17938;
   wire n17939;
   wire n17940;
   wire n17941;
   wire n17942;
   wire n17943;
   wire n17944;
   wire n17947;
   wire n17948;
   wire n17949;
   wire n17950;
   wire n17951;
   wire n17952;
   wire n17953;
   wire n17954;
   wire n17955;
   wire n17956;
   wire n17957;
   wire n17958;
   wire n17959;
   wire n17960;
   wire n17961;
   wire n17962;
   wire n17963;
   wire n17964;
   wire n17965;
   wire n17966;
   wire n17967;
   wire n17968;
   wire n17969;
   wire n17970;
   wire n17971;
   wire n17972;
   wire n17973;
   wire n17974;
   wire n17975;
   wire n17976;
   wire n17977;
   wire n17978;
   wire n17979;
   wire n17980;
   wire n17981;
   wire n17982;
   wire n17983;
   wire n17984;
   wire n17985;
   wire n17986;
   wire n17987;
   wire n17988;
   wire n17989;
   wire n17990;
   wire n17991;
   wire n17992;
   wire n17993;
   wire n17994;
   wire n17995;
   wire n17996;
   wire n17997;
   wire n17998;
   wire n17999;
   wire n18000;
   wire n18002;
   wire n18003;
   wire n18004;
   wire n18005;
   wire n18006;
   wire n18007;
   wire n18008;
   wire n18009;
   wire n18010;
   wire n18011;
   wire n18012;
   wire n18013;
   wire n18014;
   wire n18015;
   wire n18016;
   wire n18017;
   wire n18018;
   wire n18019;
   wire n18020;
   wire n18021;
   wire n18022;
   wire n18023;
   wire n18024;
   wire n18025;
   wire n18026;
   wire n18027;
   wire n18028;
   wire n18029;
   wire n18030;
   wire n18031;
   wire n18032;
   wire n18033;
   wire n18034;
   wire n18035;
   wire n18036;
   wire n18037;
   wire n18038;
   wire n18039;
   wire n18051;
   wire n18057;
   wire n18058;
   wire n18059;
   wire n18060;
   wire n18061;
   wire n18064;
   wire n18065;
   wire n18066;
   wire n18067;
   wire n18068;
   wire n18069;
   wire n18070;
   wire n18071;
   wire n18072;
   wire n18074;
   wire n18075;
   wire n18076;
   wire n18077;
   wire n18078;
   wire n18079;
   wire n18080;
   wire n18081;
   wire n18082;
   wire n18083;
   wire n18084;
   wire n18085;
   wire n18086;
   wire n18087;
   wire n18088;
   wire n18089;
   wire n18090;
   wire n18091;
   wire n18092;
   wire n18093;
   wire n18094;
   wire n18095;
   wire n18096;
   wire n18097;
   wire n18098;
   wire n18099;
   wire n18100;
   wire n18101;
   wire n18102;
   wire n18103;
   wire n18104;
   wire n18105;
   wire n18106;
   wire n18107;
   wire n18108;
   wire n18109;
   wire n18112;
   wire n18113;
   wire n18114;
   wire n18115;
   wire n18116;
   wire n18117;
   wire n18118;
   wire n18119;
   wire n18120;
   wire n18121;
   wire n18122;
   wire n18123;
   wire n18124;
   wire n18125;
   wire n18126;
   wire n18127;
   wire n18128;
   wire n18129;
   wire n18130;
   wire n18131;
   wire n18132;
   wire n18133;
   wire n18134;
   wire n18136;
   wire n18137;
   wire n18138;
   wire n18139;
   wire n18140;
   wire n18141;
   wire n18142;
   wire n18143;
   wire n18145;
   wire n18146;
   wire n18147;
   wire n18148;
   wire n18149;
   wire n18150;
   wire n18151;
   wire n18152;
   wire n18153;
   wire n18154;
   wire n18155;
   wire n18156;
   wire n18157;
   wire n18158;
   wire n18159;
   wire n18160;
   wire n18161;
   wire n18162;
   wire n18163;
   wire n18164;
   wire n18165;
   wire n18166;
   wire n18167;
   wire n18168;
   wire n18169;
   wire n18170;
   wire n18171;
   wire n18172;
   wire n18173;
   wire n18174;
   wire n18175;
   wire n18176;
   wire n18177;
   wire n18178;
   wire n18179;
   wire n18180;
   wire n18181;
   wire n18182;
   wire n18183;
   wire n18184;
   wire n18185;
   wire n18186;
   wire n18187;
   wire n18188;
   wire n18189;
   wire n18190;
   wire n18191;
   wire n18192;
   wire n18193;
   wire n18194;
   wire n18195;
   wire n18196;
   wire n18197;
   wire n18198;
   wire n18199;
   wire n18200;
   wire n18201;
   wire n18202;
   wire n18203;
   wire n18204;
   wire n18205;
   wire n18206;
   wire n18207;
   wire n18208;
   wire n18209;
   wire n18210;
   wire n18211;
   wire n18212;
   wire n18213;
   wire n18214;
   wire n18215;
   wire n18216;
   wire n18217;
   wire n18218;
   wire n18219;
   wire n18220;
   wire n18221;
   wire n18223;
   wire n18224;
   wire n18225;
   wire n18226;
   wire n18227;
   wire n18228;
   wire n18229;
   wire n18230;
   wire n18231;
   wire n18232;
   wire n18233;
   wire n18234;
   wire n18235;
   wire n18236;
   wire n18237;
   wire n18238;
   wire n18239;
   wire n18240;
   wire n18241;
   wire n18242;
   wire n18243;
   wire n18244;
   wire n18245;
   wire n18246;
   wire n18247;
   wire n18248;
   wire n18249;
   wire n18250;
   wire n18251;
   wire n18252;
   wire n18253;
   wire n18254;
   wire n18255;
   wire n18256;
   wire n18257;
   wire n18258;
   wire n18259;
   wire n18260;
   wire n18261;
   wire n18262;
   wire n18263;
   wire n18264;
   wire n18265;
   wire n18266;
   wire n18267;
   wire n18268;
   wire n18269;
   wire n18270;
   wire n18271;
   wire n18272;
   wire n18273;
   wire n18274;
   wire n18275;
   wire n18276;
   wire n18277;
   wire n18278;
   wire n18279;
   wire n18280;
   wire n18281;
   wire n18282;
   wire n18283;
   wire n18284;
   wire n18285;
   wire n18286;
   wire n18287;
   wire n18288;
   wire n18289;
   wire n18290;
   wire n18291;
   wire n18292;
   wire n18293;
   wire n18294;
   wire n18295;
   wire n18296;
   wire n18297;
   wire n18298;
   wire n18299;
   wire n18300;
   wire n18301;
   wire n18302;
   wire n18303;
   wire n18304;
   wire n18305;
   wire n18306;
   wire n18307;
   wire n18308;
   wire n18309;
   wire n18310;
   wire n18311;
   wire n18312;
   wire n18313;
   wire n18314;
   wire n18315;
   wire n18316;
   wire n18317;
   wire n18318;
   wire n18319;
   wire n18320;
   wire n18321;
   wire n18322;
   wire n18323;
   wire n18324;
   wire n18325;
   wire n18326;
   wire n18327;
   wire n18328;
   wire n18331;
   wire n18332;
   wire n18333;
   wire n18334;
   wire n18335;
   wire n18336;
   wire n18337;
   wire n18338;
   wire n18339;
   wire n18340;
   wire n18341;
   wire n18342;
   wire n18343;
   wire n18344;
   wire n18345;
   wire n18346;
   wire n18347;
   wire n18348;
   wire n18349;
   wire n18350;
   wire n18351;
   wire n18352;
   wire n18353;
   wire n18354;
   wire n18355;
   wire n18356;
   wire n18357;
   wire n18358;
   wire n18359;
   wire n18360;
   wire n18361;
   wire n18362;
   wire n18363;
   wire n18364;
   wire n18365;
   wire n18366;
   wire n18367;
   wire n18368;
   wire n18369;
   wire n18370;
   wire n18371;
   wire n18372;
   wire n18373;
   wire n18374;
   wire n18375;
   wire n18376;
   wire n18377;
   wire n18378;
   wire n18379;
   wire n18380;
   wire n18381;
   wire n18382;
   wire n18383;
   wire n18384;
   wire n18385;
   wire n18386;
   wire n18387;
   wire n18388;
   wire n18389;
   wire n18390;
   wire n18391;
   wire n18392;
   wire n18393;
   wire n18394;
   wire n18395;
   wire n18396;
   wire n18397;
   wire n18398;
   wire n18399;
   wire n18400;
   wire n18401;
   wire n18402;
   wire n18403;
   wire n18404;
   wire n18405;
   wire n18406;
   wire n18407;
   wire n18408;
   wire n18409;
   wire n18410;
   wire n18411;
   wire n18412;
   wire n18413;
   wire n18414;
   wire n18415;
   wire n18416;
   wire n18417;
   wire n18418;
   wire n18419;
   wire n18420;
   wire n18422;
   wire n18423;
   wire n18424;
   wire n18425;
   wire n18426;
   wire n18427;
   wire n18428;
   wire n18429;
   wire n18430;
   wire n18431;
   wire n18432;
   wire n18433;
   wire n18434;
   wire n18435;
   wire n18436;
   wire n18437;
   wire n18438;
   wire n18439;
   wire n18440;
   wire n18441;
   wire n18442;
   wire n18443;
   wire n18444;
   wire n18445;
   wire n18446;
   wire n18447;
   wire n18448;
   wire n18449;
   wire n18450;
   wire n18451;
   wire n18452;
   wire n18453;
   wire n18454;
   wire n18455;
   wire n18456;
   wire n18457;
   wire n18458;
   wire n18459;
   wire n18460;
   wire n18461;
   wire n18462;
   wire n18463;
   wire n18464;
   wire n18465;
   wire n18466;
   wire n18467;
   wire n18468;
   wire n18469;
   wire n18470;
   wire n18471;
   wire n18472;
   wire n18473;
   wire n18474;
   wire n18475;
   wire n18476;
   wire n18477;
   wire n18478;
   wire n18479;
   wire n18480;
   wire n18481;
   wire n18482;
   wire n18483;
   wire n18484;
   wire n18485;
   wire n18486;
   wire n18487;
   wire n18488;
   wire n18489;
   wire n18490;
   wire n18491;
   wire n18492;
   wire n18493;
   wire n18494;
   wire n18495;
   wire n18496;
   wire n18497;
   wire n18498;
   wire n18499;
   wire n18500;
   wire n18501;
   wire n18502;
   wire n18503;
   wire n18504;
   wire n18505;
   wire n18506;
   wire n18507;
   wire n18508;
   wire n18509;
   wire n18510;
   wire n18511;
   wire n18512;
   wire n18513;
   wire n18514;
   wire n18515;
   wire n18516;
   wire n18517;
   wire n18518;
   wire n18519;
   wire n18520;
   wire n18521;
   wire n18522;
   wire n18523;
   wire n18524;
   wire n18525;
   wire n18526;
   wire n18527;
   wire n18528;
   wire n18529;
   wire n18530;
   wire n18531;
   wire n18532;
   wire n18533;
   wire n18534;
   wire n18535;
   wire n18536;
   wire n18537;
   wire n18538;
   wire n18539;
   wire n18540;
   wire n18541;
   wire n18542;
   wire n18543;
   wire n18544;
   wire n18545;
   wire n18546;
   wire n18547;
   wire n18548;
   wire n18549;
   wire n18550;
   wire n18551;
   wire n18552;
   wire n18553;
   wire n18554;
   wire n18555;
   wire n18556;
   wire n18557;
   wire n18558;
   wire n18559;
   wire n18560;
   wire n18561;
   wire n18562;
   wire n18563;
   wire n18564;
   wire n18565;
   wire n18566;
   wire n18567;
   wire n18568;
   wire n18569;
   wire n18570;
   wire n18571;
   wire n18572;
   wire n18573;
   wire n18574;
   wire n18575;
   wire n18576;
   wire n18577;
   wire n18578;
   wire n18579;
   wire n18580;
   wire n18581;
   wire n18582;
   wire n18583;
   wire n18584;
   wire n18585;
   wire n18586;
   wire n18587;
   wire n18588;
   wire n18589;
   wire n18591;
   wire n18592;
   wire n18593;
   wire n18594;
   wire n18595;
   wire n18596;
   wire n18597;
   wire n18598;
   wire n18599;
   wire n18600;
   wire n18601;
   wire n18602;
   wire n18603;
   wire n18604;
   wire n18605;
   wire n18606;
   wire n18607;
   wire n18608;
   wire n18609;
   wire n18610;
   wire n18611;
   wire n18612;
   wire n18613;
   wire n18614;
   wire n18615;
   wire n18616;
   wire n18617;
   wire n18618;
   wire n18619;
   wire n18620;
   wire n18621;
   wire n18622;
   wire n18623;
   wire n18624;
   wire n18625;
   wire n18626;
   wire n18627;
   wire n18628;
   wire n18629;
   wire n18630;
   wire n18631;
   wire n18632;
   wire n18633;
   wire n18634;
   wire n18635;
   wire n18636;
   wire n18637;
   wire n18638;
   wire n18639;
   wire n18640;
   wire n18641;
   wire n18642;
   wire n18643;
   wire n18644;
   wire n18645;
   wire n18646;
   wire n18647;
   wire n18648;
   wire n18649;
   wire n18650;
   wire n18651;
   wire n18652;
   wire n18653;
   wire n18654;
   wire n18655;
   wire n18656;
   wire n18657;
   wire n18658;
   wire n18659;
   wire n18660;
   wire n18661;
   wire n18662;
   wire n18663;
   wire n18664;
   wire n18665;
   wire n18666;
   wire n18667;
   wire n18668;
   wire n18669;
   wire n18670;
   wire n18671;
   wire n18672;
   wire n18673;
   wire n18674;
   wire n18675;
   wire n18676;
   wire n18677;
   wire n18678;
   wire n18679;
   wire n18680;
   wire n18681;
   wire n18682;
   wire n18683;
   wire n18684;
   wire n18685;
   wire n18686;
   wire n18687;
   wire n18688;
   wire n18689;
   wire n18690;
   wire n18691;
   wire n18692;
   wire n18693;
   wire n18694;
   wire n18695;
   wire n18696;
   wire n18697;
   wire n18698;
   wire n18699;
   wire n18700;
   wire n18701;
   wire n18702;
   wire n18703;
   wire n18704;
   wire n18705;
   wire n18706;
   wire n18707;
   wire n18708;
   wire n18709;
   wire n18710;
   wire n18711;
   wire n18712;
   wire n18713;
   wire n18714;
   wire n18715;
   wire n18716;
   wire n18717;
   wire n18718;
   wire n18719;
   wire n18720;
   wire n18721;
   wire n18722;
   wire n18723;
   wire n18724;
   wire n18725;
   wire n18726;
   wire n18727;
   wire n18728;
   wire n18729;
   wire n18730;
   wire n18731;
   wire n18732;
   wire n18733;
   wire n18734;
   wire n18735;
   wire n18736;
   wire n18737;
   wire n18738;
   wire n18739;
   wire n18740;
   wire n18741;
   wire n18742;
   wire n18743;
   wire n18744;
   wire n18745;
   wire n18746;
   wire n18747;
   wire n18748;
   wire n18749;
   wire n18750;
   wire n18751;
   wire n18752;
   wire n18753;
   wire n18754;
   wire n18755;
   wire n18756;
   wire n18757;
   wire n18758;
   wire n18759;
   wire n18760;
   wire n18761;
   wire n18762;
   wire n18763;
   wire n18764;
   wire n18765;
   wire n18766;
   wire n18767;
   wire n18768;
   wire n18769;
   wire n18770;
   wire n18771;
   wire n18772;
   wire n18773;
   wire n18774;
   wire n18775;
   wire n18776;
   wire n18777;
   wire n18778;
   wire n18779;
   wire n18780;
   wire n18781;
   wire n18782;
   wire n18783;
   wire n18784;
   wire n18785;
   wire n18786;
   wire n18787;
   wire n18788;
   wire n18789;
   wire n18790;
   wire n18791;
   wire n18792;
   wire n18793;
   wire n18794;
   wire n18795;
   wire n18796;
   wire n18797;
   wire n18798;
   wire n18799;
   wire n18800;
   wire n18801;
   wire n18802;
   wire n18803;
   wire n18804;
   wire n18805;
   wire n18806;
   wire n18807;
   wire n18808;
   wire n18809;
   wire n18810;
   wire n18811;
   wire n18812;
   wire n18813;
   wire n18814;
   wire n18815;
   wire n18816;
   wire n18817;
   wire n18818;
   wire n18819;
   wire n18820;
   wire n18821;
   wire n18822;
   wire n18823;
   wire n18824;
   wire n18825;
   wire n18826;
   wire n18827;
   wire n18828;
   wire n18829;
   wire n18830;
   wire n18831;
   wire n18832;
   wire n18833;
   wire n18834;
   wire n18835;
   wire n18836;
   wire n18837;
   wire n18838;
   wire n18839;
   wire n18840;
   wire n18841;
   wire n18842;
   wire n18843;
   wire n18844;
   wire n18845;
   wire n18846;
   wire n18847;
   wire n18848;
   wire n18849;
   wire n18850;
   wire n18851;
   wire n18852;
   wire n18853;
   wire n18854;
   wire n18855;
   wire n18856;
   wire n18857;
   wire n18858;
   wire n18859;
   wire n18860;
   wire n18861;
   wire n18862;
   wire n18863;
   wire n18864;
   wire n18865;
   wire n18866;
   wire n18867;
   wire n18868;
   wire n18869;
   wire n18870;
   wire n18871;
   wire n18872;
   wire n18873;
   wire n18874;
   wire n18875;
   wire n18876;
   wire n18877;
   wire n18878;
   wire n18879;
   wire n18880;
   wire n18881;
   wire n18882;
   wire n18883;
   wire n18884;
   wire n18885;
   wire n18886;
   wire n18887;
   wire n18888;
   wire n18889;
   wire n18890;
   wire n18891;
   wire n18892;
   wire n18893;
   wire n18894;
   wire n18895;
   wire n18896;
   wire n18897;
   wire n18898;
   wire n18899;
   wire n18900;
   wire n18901;
   wire n18902;
   wire n18903;
   wire n18904;
   wire n18905;
   wire n18906;
   wire n18907;
   wire n18908;
   wire n18909;
   wire n18910;
   wire n18911;
   wire n18912;
   wire n18913;
   wire n18914;
   wire n18915;
   wire n18916;
   wire n18917;
   wire n18918;
   wire n18919;
   wire n18920;
   wire n18921;
   wire n18922;
   wire n18923;
   wire n18924;
   wire n18925;
   wire n18926;
   wire n18927;
   wire n18928;
   wire n18929;
   wire n18930;
   wire n18931;
   wire n18932;
   wire n18933;
   wire n18934;
   wire n18935;
   wire n18936;
   wire n18937;
   wire n18938;
   wire n18939;
   wire n18940;
   wire n18941;
   wire n18942;
   wire n18943;
   wire n18944;
   wire n18945;
   wire n18946;
   wire n18947;
   wire n18948;
   wire n18950;
   wire n18951;
   wire n18952;
   wire n18953;
   wire n18954;
   wire n18955;
   wire n18956;
   wire n18957;
   wire n18958;
   wire n18959;
   wire n18960;
   wire n18961;
   wire n18962;
   wire n18963;
   wire n18964;
   wire n18965;
   wire n18966;
   wire n18967;
   wire n18968;
   wire n18969;
   wire n18970;
   wire n18971;
   wire n18972;
   wire n18973;
   wire n18974;
   wire n18975;
   wire n18976;
   wire n18977;
   wire n18978;
   wire n18979;
   wire n18980;
   wire n18981;
   wire n18982;
   wire n18983;
   wire n18984;
   wire n18985;
   wire n18986;
   wire n18987;
   wire n18988;
   wire n18989;
   wire n18990;
   wire n18991;
   wire n18992;
   wire n18993;
   wire n18994;
   wire n18995;
   wire n18996;
   wire n18997;
   wire n18998;
   wire n18999;
   wire n19000;
   wire n19001;
   wire n19002;
   wire n19003;
   wire n19004;
   wire n19005;
   wire n19006;
   wire n19007;
   wire n19008;
   wire n19009;
   wire n19010;
   wire n19011;
   wire n19012;
   wire n19013;
   wire n19014;
   wire n19015;
   wire n19016;
   wire n19017;
   wire n19018;
   wire n19019;
   wire n19020;
   wire n19021;
   wire n19022;
   wire n19023;
   wire n19024;
   wire n19025;
   wire n19026;
   wire n19027;
   wire n19028;
   wire n19029;
   wire n19030;
   wire n19031;
   wire n19032;
   wire n19033;
   wire n19034;
   wire n19035;
   wire n19036;
   wire n19037;
   wire n19038;
   wire n19039;
   wire n19040;
   wire n19041;
   wire n19042;
   wire n19043;
   wire n19044;
   wire n19045;
   wire n19046;
   wire n19047;
   wire n19048;
   wire n19049;
   wire n19050;
   wire n19051;
   wire n19052;
   wire n19053;
   wire n19054;
   wire n19055;
   wire n19056;
   wire n19057;
   wire n19058;
   wire n19059;
   wire n19060;
   wire n19061;
   wire n19062;
   wire n19063;
   wire n19064;
   wire n19065;
   wire n19066;
   wire n19067;
   wire n19068;
   wire n19069;
   wire n19070;
   wire n19071;
   wire n19072;
   wire n19073;
   wire n19074;
   wire n19075;
   wire n19076;
   wire n19077;
   wire n19078;
   wire n19079;
   wire n19080;
   wire n19081;
   wire n19082;
   wire n19083;
   wire n19084;
   wire n19085;
   wire n19086;
   wire n19087;
   wire n19088;
   wire n19089;
   wire n19090;
   wire n19091;
   wire n19092;
   wire n19093;
   wire n19094;
   wire n19095;
   wire n19096;
   wire n19097;
   wire n19098;
   wire n19099;
   wire n19100;
   wire n19101;
   wire n19102;
   wire n19103;
   wire n19104;
   wire n19105;
   wire n19106;
   wire n19107;
   wire n19108;
   wire n19109;
   wire n19110;
   wire n19111;
   wire n19112;
   wire n19113;
   wire n19114;
   wire n19115;
   wire n19116;
   wire n19117;
   wire n19118;
   wire n19119;
   wire n19120;
   wire n19121;
   wire n19122;
   wire n19123;
   wire n19124;
   wire n19125;
   wire n19126;
   wire n19127;
   wire n19128;
   wire n19129;
   wire n19130;
   wire n19131;
   wire n19132;
   wire n19133;
   wire n19134;
   wire n19135;
   wire n19136;
   wire n19137;
   wire n19138;
   wire n19139;
   wire n19140;
   wire n19141;
   wire n19142;
   wire n19143;
   wire n19144;
   wire n19145;
   wire n19146;
   wire n19147;
   wire n19148;
   wire n19149;
   wire n19150;
   wire n19151;
   wire n19152;
   wire n19153;
   wire n19154;
   wire n19155;
   wire n19156;
   wire n19157;
   wire n19158;
   wire n19159;
   wire n19160;
   wire n19161;
   wire n19162;
   wire n19163;
   wire n19164;
   wire n19165;
   wire n19166;
   wire n19167;
   wire n19168;
   wire n19169;
   wire n19170;
   wire n19171;
   wire n19172;
   wire n19173;
   wire n19174;
   wire n19175;
   wire n19176;
   wire n19177;
   wire n19178;
   wire n19179;
   wire n19180;
   wire n19181;
   wire n19182;
   wire n19183;
   wire n19184;
   wire n19185;
   wire n19186;
   wire n19187;
   wire n19188;
   wire n19189;
   wire n19190;
   wire n19191;
   wire n19192;
   wire n19193;
   wire n19194;
   wire n19195;
   wire n19196;
   wire n19197;
   wire n19198;
   wire n19199;
   wire n19200;
   wire n19201;
   wire n19202;
   wire n19203;
   wire n19204;
   wire n19205;
   wire n19206;
   wire n19207;
   wire n19208;
   wire n19209;
   wire n19210;
   wire n19211;
   wire n19212;
   wire n19213;
   wire n19214;
   wire n19215;
   wire n19216;
   wire n19217;
   wire n19218;
   wire n19219;
   wire n19220;
   wire n19221;
   wire n19222;
   wire n19223;
   wire n19224;
   wire n19225;
   wire n19226;
   wire n19227;
   wire n19228;
   wire n19229;
   wire n19230;
   wire n19231;
   wire n19232;
   wire n19233;
   wire n19234;
   wire n19235;
   wire n19236;
   wire n19237;
   wire n19238;
   wire n19239;
   wire n19240;
   wire n19241;
   wire n19242;
   wire n19243;
   wire n19244;
   wire n19245;
   wire n19246;
   wire n19247;
   wire n19248;
   wire n19249;
   wire n19250;
   wire n19251;
   wire n19252;
   wire n19253;
   wire n19254;
   wire n19255;
   wire n19256;
   wire n19257;
   wire n19258;
   wire n19259;
   wire n19260;
   wire n19261;
   wire n19262;
   wire n19263;
   wire n19264;
   wire n19265;
   wire n19266;
   wire n19267;
   wire n19268;
   wire n19269;
   wire n19270;
   wire n19271;
   wire n19272;
   wire n19273;
   wire n19274;
   wire n19275;
   wire n19276;
   wire n19277;
   wire n19278;
   wire n19279;
   wire n19280;
   wire n19281;
   wire n19282;
   wire n19283;
   wire n19284;
   wire n19285;
   wire n19286;
   wire n19287;
   wire n19288;
   wire n19289;
   wire n19290;
   wire n19291;
   wire n19292;
   wire n19293;
   wire n19294;
   wire n19295;
   wire n19296;
   wire n19297;
   wire n19298;
   wire n19299;
   wire n19300;
   wire n19301;
   wire n19302;
   wire n19303;
   wire n19304;
   wire n19305;
   wire n19306;
   wire n19307;
   wire n19308;
   wire n19309;
   wire n19310;
   wire n19311;
   wire n19312;
   wire n19313;
   wire n19314;
   wire n19315;
   wire n19316;
   wire n19317;
   wire n19318;
   wire n19319;
   wire n19320;
   wire n19321;
   wire n19322;
   wire n19323;
   wire n19324;
   wire n19325;
   wire n19326;
   wire n19327;
   wire n19328;
   wire n19329;
   wire n19330;
   wire n19331;
   wire n19332;
   wire n19333;
   wire n19334;
   wire n19335;
   wire n19336;
   wire n19337;
   wire n19338;
   wire n19339;
   wire n19340;
   wire n19341;
   wire n19342;
   wire n19343;
   wire n19344;
   wire n19345;
   wire n19346;
   wire n19347;
   wire n19348;
   wire n19349;
   wire n19350;
   wire n19351;
   wire n19352;
   wire n19353;
   wire n19354;
   wire n19356;
   wire n19357;
   wire n19358;
   wire n19359;
   wire n19360;
   wire n19361;
   wire n19362;
   wire n19363;
   wire n19364;
   wire n19365;
   wire n19366;
   wire n19367;
   wire n19368;
   wire n19369;
   wire n19370;
   wire n19371;
   wire n19372;
   wire n19373;
   wire n19374;
   wire n19375;
   wire n19376;
   wire n19377;
   wire n19378;
   wire n19379;
   wire n19380;
   wire n19381;
   wire n19382;
   wire n19383;
   wire n19384;
   wire n19385;
   wire n19386;
   wire n19387;
   wire n19388;
   wire n19389;
   wire n19390;
   wire n19391;
   wire n19392;
   wire n19393;
   wire n19394;
   wire n19395;
   wire n19396;
   wire n19397;
   wire n19398;
   wire n19399;
   wire n19400;
   wire n19401;
   wire n19402;
   wire n19403;
   wire n19404;
   wire n19405;
   wire n19406;
   wire n19407;
   wire n19408;
   wire n19409;
   wire n19410;
   wire n19411;
   wire n19412;
   wire n19413;
   wire n19414;
   wire n19415;
   wire n19416;
   wire n19417;
   wire n19418;
   wire n19419;
   wire n19420;
   wire n19421;
   wire n19422;
   wire n19423;
   wire n19424;
   wire n19425;
   wire n19426;
   wire n19427;
   wire n19428;
   wire n19429;
   wire n19430;
   wire n19431;
   wire n19432;
   wire n19433;
   wire n19435;
   wire n19436;
   wire n19437;
   wire n19438;
   wire n19439;
   wire n19440;
   wire n19441;
   wire n19442;
   wire n19443;
   wire n19444;
   wire n19445;
   wire n19446;
   wire n19447;
   wire n19448;
   wire n19449;
   wire n19450;
   wire n19451;
   wire n19452;
   wire n19453;
   wire n19454;
   wire n19455;
   wire n19456;
   wire n19457;
   wire n19458;
   wire n19459;
   wire n19460;
   wire n19461;
   wire n19462;
   wire n19463;
   wire n19464;
   wire n19465;
   wire n19466;
   wire n19467;
   wire n19468;
   wire n19469;
   wire n19470;
   wire n19471;
   wire n19472;
   wire n19473;
   wire n19474;
   wire n19475;
   wire n19476;
   wire n19477;
   wire n19478;
   wire n19479;
   wire n19480;
   wire n19481;
   wire n19482;
   wire n19483;
   wire n19484;
   wire n19485;
   wire n19486;
   wire n19487;
   wire n19488;
   wire n19489;
   wire n19490;
   wire n19491;
   wire n19492;
   wire n19493;
   wire n19494;
   wire n19495;
   wire n19496;
   wire n19497;
   wire n19498;
   wire n19499;
   wire n19500;
   wire n19501;
   wire n19502;
   wire n19503;
   wire n19504;
   wire n19505;
   wire n19506;
   wire n19507;
   wire n19508;
   wire n19509;
   wire n19510;
   wire n19511;
   wire n19512;
   wire n19514;
   wire n19515;
   wire n19516;
   wire n19517;
   wire n19518;
   wire n19519;
   wire n19520;
   wire n19521;
   wire n19522;
   wire n19523;
   wire n19524;
   wire n19525;
   wire n19526;
   wire n19527;
   wire n19528;
   wire n19529;
   wire n19530;
   wire n19531;
   wire n19532;
   wire n19533;
   wire n19534;
   wire n19535;
   wire n19536;
   wire n19537;
   wire n19538;
   wire n19539;
   wire n19540;
   wire n19541;
   wire n19543;
   wire n19544;
   wire n19545;
   wire n19546;
   wire n19547;
   wire n19549;
   wire n19550;
   wire n19551;
   wire n19552;
   wire n19553;
   wire n19554;
   wire n19555;
   wire n19556;
   wire n19557;
   wire n19558;
   wire n19559;
   wire n19560;
   wire n19561;
   wire n19562;
   wire n19563;
   wire n19564;
   wire n19565;
   wire n19566;
   wire n19567;
   wire n19568;
   wire n19569;
   wire n19570;
   wire n19571;
   wire n19572;
   wire n19573;
   wire n19574;
   wire n19575;
   wire n19576;
   wire n19577;
   wire n19578;
   wire n19579;
   wire n19580;
   wire n19581;
   wire n19582;
   wire n19583;
   wire n19584;
   wire n19585;
   wire n19586;
   wire n19587;
   wire n19588;
   wire n19589;
   wire n19590;
   wire n19591;
   wire n19592;
   wire n19593;
   wire n19594;
   wire n19595;
   wire n19596;
   wire n19597;
   wire n19598;
   wire n19599;
   wire n19600;
   wire n19601;
   wire n19602;
   wire n19603;
   wire n19604;
   wire n19605;
   wire n19606;
   wire n19607;
   wire n19608;
   wire n19609;
   wire n19610;
   wire n19611;
   wire n19612;
   wire n19613;
   wire n19614;
   wire n19615;
   wire n19616;
   wire n19617;
   wire n19618;
   wire n19619;
   wire n19620;
   wire n19621;
   wire n19622;
   wire n19623;
   wire n19624;
   wire n19625;
   wire n19626;
   wire n19627;
   wire n19629;
   wire n19630;
   wire n19632;
   wire n19633;
   wire n19634;
   wire n19635;
   wire n19636;
   wire n19637;
   wire n19638;
   wire n19639;
   wire n19640;
   wire n19641;
   wire n19642;
   wire n19643;
   wire n19644;
   wire n19645;
   wire n19646;
   wire n19647;
   wire n19648;
   wire n19649;
   wire n19650;
   wire n19651;
   wire n19652;
   wire n19654;
   wire n19655;
   wire n19656;
   wire n19657;
   wire n19658;
   wire n19659;
   wire n19660;
   wire n19661;
   wire n19662;
   wire n19663;
   wire n19665;
   wire n19666;
   wire n19667;
   wire n19668;
   wire n19669;
   wire n19670;
   wire n19671;
   wire n19672;
   wire n19673;
   wire n19674;
   wire n19675;
   wire n19676;
   wire n19677;
   wire n19678;
   wire n19679;
   wire n19680;
   wire n19681;
   wire n19682;
   wire n19683;
   wire n19684;
   wire n19685;
   wire n19686;
   wire n19687;
   wire n19688;
   wire n19689;
   wire n19690;
   wire n19691;
   wire n19692;
   wire n19693;
   wire n19694;
   wire n19695;
   wire n19696;
   wire n19697;
   wire n19698;
   wire n19699;
   wire n19700;
   wire n19701;
   wire n19702;
   wire n19703;
   wire n19704;
   wire n19705;
   wire n19706;
   wire n19707;
   wire n19708;
   wire n19709;
   wire n19710;
   wire n19711;
   wire n19712;
   wire n19713;
   wire n19714;
   wire n19715;
   wire n19716;
   wire n19717;
   wire n19718;
   wire n19719;
   wire n19720;
   wire n19721;
   wire n19722;
   wire n19723;
   wire n19724;
   wire n19725;
   wire n19726;
   wire n19727;
   wire n19728;
   wire n19729;
   wire n19730;
   wire n19731;
   wire n19732;
   wire n19733;
   wire n19734;
   wire n19735;
   wire n19736;
   wire n19737;
   wire n19738;
   wire n19739;
   wire n19740;
   wire n19741;
   wire n19742;
   wire n19743;
   wire n19744;
   wire n19745;
   wire n19746;
   wire n19747;
   wire n19748;
   wire n19749;
   wire n19750;
   wire n19751;
   wire n19752;
   wire n19753;
   wire n19754;
   wire n19755;
   wire n19756;
   wire n19757;
   wire n19758;
   wire n19759;
   wire n19760;
   wire n19761;
   wire n19762;
   wire n19763;
   wire n19764;
   wire n19765;
   wire n19766;
   wire n19767;
   wire n19769;
   wire n19770;
   wire n19771;
   wire n19772;
   wire n19773;
   wire n19774;
   wire n19775;
   wire n19776;
   wire n19777;
   wire n19778;
   wire n19779;
   wire n19780;
   wire n19781;
   wire n19782;
   wire n19783;
   wire n19784;
   wire n19785;
   wire n19786;
   wire n19787;
   wire n19788;
   wire n19789;
   wire n19790;
   wire n19791;
   wire n19792;
   wire n19793;
   wire n19794;
   wire n19795;
   wire n19796;
   wire n19797;
   wire n19798;
   wire n19799;
   wire n19800;
   wire n19801;
   wire n19802;
   wire n19803;
   wire n19804;
   wire n19805;
   wire n19806;
   wire n19807;
   wire n19808;
   wire n19809;
   wire n19810;
   wire n19811;
   wire n19812;
   wire n19813;
   wire n19814;
   wire n19815;
   wire n19816;
   wire n19817;
   wire n19818;
   wire n19819;
   wire n19820;
   wire n19821;
   wire n19822;
   wire n19823;
   wire n19824;
   wire n19825;
   wire n19826;
   wire n19827;
   wire n19828;
   wire n19829;
   wire n19830;
   wire n19831;
   wire n19832;
   wire n19833;
   wire n19834;
   wire n19835;
   wire n19836;
   wire n19837;
   wire n19838;
   wire n19839;
   wire n19840;
   wire n19841;
   wire n19842;
   wire n19843;
   wire n19844;
   wire n19845;
   wire n19846;
   wire n19847;
   wire n19848;
   wire n19849;
   wire n19850;
   wire n19851;
   wire n19852;
   wire n19853;
   wire n19854;
   wire n19855;
   wire n19856;
   wire n19857;
   wire n19858;
   wire n19859;
   wire n19860;
   wire n19861;
   wire n19862;
   wire n19863;
   wire n19864;
   wire n19865;
   wire n19866;
   wire n19867;
   wire n19868;
   wire n19869;
   wire n19870;
   wire n19871;
   wire n19872;
   wire n19873;
   wire n19874;
   wire n19875;
   wire n19876;
   wire n19877;
   wire n19878;
   wire n19879;
   wire n19880;
   wire n19881;
   wire n19882;
   wire n19883;
   wire n19884;
   wire n19885;
   wire n19886;
   wire n19887;
   wire n19888;
   wire n19889;
   wire n19890;
   wire n19891;
   wire n19892;
   wire n19893;
   wire n19894;
   wire n19895;
   wire n19896;
   wire n19897;
   wire n19898;
   wire n19899;
   wire n19900;
   wire n19901;
   wire n19902;
   wire n19903;
   wire n19904;
   wire n19905;
   wire n19906;
   wire n19907;
   wire n19908;
   wire n19909;
   wire n19910;
   wire n19911;
   wire n19912;
   wire n19913;
   wire n19914;
   wire n19915;
   wire n19916;
   wire n19917;
   wire n19918;
   wire n19919;
   wire n19920;
   wire n19921;
   wire n19922;
   wire n19923;
   wire n19924;
   wire n19925;
   wire n19926;
   wire n19927;
   wire n19928;
   wire n19930;
   wire n19931;
   wire n19932;
   wire n19933;
   wire n19934;
   wire n19935;
   wire n19936;
   wire n19937;
   wire n19938;
   wire n19939;
   wire n19940;
   wire n19941;
   wire n19942;
   wire n19943;
   wire n19944;
   wire n19945;
   wire n19946;
   wire n19947;
   wire n19948;
   wire n19949;
   wire n19950;
   wire n19951;
   wire n19952;
   wire n19953;
   wire n19954;
   wire n19955;
   wire n19956;
   wire n19957;
   wire n19958;
   wire n19959;
   wire n19960;
   wire n19961;
   wire n19962;
   wire n19963;
   wire n19964;
   wire n19965;
   wire n19966;
   wire n19967;
   wire n19968;
   wire n19969;
   wire n19970;
   wire n19971;
   wire n19972;
   wire n19973;
   wire n19974;
   wire n19975;
   wire n19976;
   wire n19977;
   wire n19978;
   wire n19979;
   wire n19980;
   wire n19981;
   wire n19982;
   wire n19983;
   wire n19984;
   wire n19985;
   wire n19986;
   wire n19987;
   wire n19988;
   wire n19989;
   wire n19990;
   wire n19991;
   wire n19992;
   wire n19993;
   wire n19994;
   wire n19995;
   wire n19996;
   wire n19997;
   wire n19998;
   wire n19999;
   wire n20000;
   wire n20001;
   wire n20002;
   wire n20003;
   wire n20004;
   wire n20005;
   wire n20006;
   wire n20007;
   wire n20008;
   wire n20009;
   wire n20010;
   wire n20011;
   wire n20012;
   wire n20013;
   wire n20014;
   wire n20015;
   wire n20016;
   wire n20017;
   wire n20018;
   wire n20019;
   wire n20020;
   wire n20021;
   wire n20022;
   wire n20023;
   wire n20024;
   wire n20025;
   wire n20026;
   wire n20027;
   wire n20028;
   wire n20029;
   wire n20030;
   wire n20031;
   wire n20032;
   wire n20033;
   wire n20034;
   wire n20035;
   wire n20036;
   wire n20037;
   wire n20038;
   wire n20039;
   wire n20040;
   wire n20041;
   wire n20042;
   wire n20043;
   wire n20044;
   wire n20045;
   wire n20046;
   wire n20047;
   wire n20048;
   wire n20050;
   wire n20051;
   wire n20052;
   wire n20053;
   wire n20054;
   wire n20055;
   wire n20056;
   wire n20057;
   wire n20058;
   wire n20059;
   wire n20060;
   wire n20061;
   wire n20062;
   wire n20063;
   wire n20064;
   wire n20065;
   wire n20066;
   wire n20067;
   wire n20068;
   wire n20069;
   wire n20070;
   wire n20071;
   wire n20072;
   wire n20073;
   wire n20074;
   wire n20075;
   wire n20076;
   wire n20077;
   wire n20078;
   wire n20079;
   wire n20080;
   wire n20081;
   wire n20082;
   wire n20083;
   wire n20084;
   wire n20085;
   wire n20086;
   wire n20087;
   wire n20088;
   wire n20089;
   wire n20090;
   wire n20091;
   wire n20092;
   wire n20093;
   wire n20094;
   wire n20095;
   wire n20096;
   wire n20097;
   wire n20098;
   wire n20099;
   wire n20100;
   wire n20101;
   wire n20102;
   wire n20103;
   wire n20104;
   wire n20105;
   wire n20106;
   wire n20107;
   wire n20108;
   wire n20109;
   wire n20110;
   wire n20111;
   wire n20112;
   wire n20113;
   wire n20114;
   wire n20115;
   wire n20116;
   wire n20117;
   wire n20118;
   wire n20119;
   wire n20120;
   wire n20121;
   wire n20122;
   wire n20123;
   wire n20124;
   wire n20125;
   wire n20126;
   wire n20127;
   wire n20128;
   wire n20129;
   wire n20130;
   wire n20131;
   wire n20132;
   wire n20133;
   wire n20134;
   wire n20135;
   wire n20136;
   wire n20137;
   wire n20138;
   wire n20139;
   wire n20140;
   wire n20141;
   wire n20142;
   wire n20143;
   wire n20144;
   wire n20145;
   wire n20146;
   wire n20147;
   wire n20148;
   wire n20149;
   wire n20150;
   wire n20151;
   wire n20152;
   wire n20153;
   wire n20154;
   wire n20155;
   wire n20156;
   wire n20157;
   wire n20158;
   wire n20159;
   wire n20160;
   wire n20161;
   wire n20162;
   wire n20163;
   wire n20164;
   wire n20165;
   wire n20166;
   wire n20167;
   wire n20168;
   wire n20169;
   wire n20170;
   wire n20171;
   wire n20172;
   wire n20173;
   wire n20174;
   wire n20175;
   wire n20176;
   wire n20177;
   wire n20178;
   wire n20179;
   wire n20180;
   wire n20181;
   wire n20182;
   wire n20183;
   wire n20184;
   wire n20185;
   wire n20186;
   wire n20187;
   wire n20188;
   wire n20189;
   wire n20190;
   wire n20191;
   wire n20192;
   wire n20193;
   wire n20194;
   wire n20195;
   wire n20196;
   wire n20197;
   wire n20198;
   wire n20199;
   wire n20200;
   wire n20201;
   wire n20202;
   wire n20203;
   wire n20204;
   wire n20205;
   wire n20206;
   wire n20207;
   wire n20208;
   wire n20209;
   wire n20210;
   wire n20211;
   wire n20212;
   wire n20213;
   wire n20214;
   wire n20215;
   wire n20216;
   wire n20217;
   wire n20218;
   wire n20219;
   wire n20220;
   wire n20221;
   wire n20222;
   wire n20223;
   wire n20224;
   wire n20225;
   wire n20226;
   wire n20227;
   wire n20228;
   wire n20229;
   wire n20230;
   wire n20231;
   wire n20232;
   wire n20233;
   wire n20234;
   wire n20235;
   wire n20236;
   wire n20237;
   wire n20238;
   wire n20239;
   wire n20240;
   wire n20241;
   wire n20242;
   wire n20243;
   wire n20244;
   wire n20245;
   wire n20246;
   wire n20247;
   wire n20248;
   wire n20249;
   wire n20250;
   wire n20251;
   wire n20252;
   wire n20253;
   wire n20254;
   wire n20256;
   wire n20257;
   wire n20258;
   wire n20259;
   wire n20260;
   wire n20261;
   wire n20262;
   wire n20263;
   wire n20264;
   wire n20265;
   wire n20266;
   wire n20267;
   wire n20268;
   wire n20269;
   wire n20270;
   wire n20271;
   wire n20272;
   wire n20273;
   wire n20274;
   wire n20275;
   wire n20276;
   wire n20277;
   wire n20278;
   wire n20279;
   wire n20280;
   wire n20281;
   wire n20282;
   wire n20283;
   wire n20284;
   wire n20285;
   wire n20286;
   wire n20287;
   wire n20288;
   wire n20289;
   wire n20290;
   wire n20291;
   wire n20292;
   wire n20293;
   wire n20294;
   wire n20295;
   wire n20296;
   wire n20297;
   wire n20298;
   wire n20299;
   wire n20300;
   wire n20301;
   wire n20302;
   wire n20303;
   wire n20304;
   wire n20305;
   wire n20306;
   wire n20307;
   wire n20308;
   wire n20309;
   wire n20310;
   wire n20311;
   wire n20312;
   wire n20313;
   wire n20314;
   wire n20315;
   wire n20316;
   wire n20317;
   wire n20318;
   wire n20319;
   wire n20320;
   wire n20321;
   wire n20322;
   wire n20323;
   wire n20324;
   wire n20325;
   wire n20326;
   wire n20327;
   wire n20328;
   wire n20329;
   wire n20330;
   wire n20331;
   wire n20332;
   wire n20333;
   wire n20334;
   wire n20335;
   wire n20336;
   wire n20337;
   wire n20338;
   wire n20339;
   wire n20340;
   wire n20341;
   wire n20342;
   wire n20343;
   wire n20344;
   wire n20345;
   wire n20346;
   wire n20347;
   wire n20348;
   wire n20349;
   wire n20350;
   wire n20351;
   wire n20352;
   wire n20353;
   wire n20354;
   wire n20355;
   wire n20356;
   wire n20357;
   wire n20358;
   wire n20359;
   wire n20360;
   wire n20361;
   wire n20362;
   wire n20363;
   wire n20364;
   wire n20365;
   wire n20366;
   wire n20367;
   wire n20368;
   wire n20369;
   wire n20370;
   wire n20371;
   wire n20372;
   wire n20373;
   wire n20374;
   wire n20375;
   wire n20376;
   wire n20377;
   wire n20378;
   wire n20379;
   wire n20380;
   wire n20381;
   wire n20382;
   wire n20383;
   wire n20384;
   wire n20385;
   wire n20386;
   wire n20387;
   wire n20388;
   wire n20389;
   wire n20390;
   wire n20391;
   wire n20392;
   wire n20393;
   wire n20394;
   wire n20395;
   wire n20396;
   wire n20397;
   wire n20398;
   wire n20399;
   wire n20400;
   wire n20401;
   wire n20402;
   wire n20403;
   wire n20404;
   wire n20405;
   wire n20406;
   wire n20407;
   wire n20408;
   wire n20409;
   wire n20410;
   wire n20411;
   wire n20412;
   wire n20413;
   wire n20414;
   wire n20415;
   wire n20416;
   wire n20417;
   wire n20418;
   wire n20419;
   wire n20420;
   wire n20421;
   wire n20422;
   wire n20423;
   wire n20424;
   wire n20425;
   wire n20426;
   wire n20427;
   wire n20428;
   wire n20429;
   wire n20430;
   wire n20431;
   wire n20432;
   wire n20433;
   wire n20434;
   wire n20435;
   wire n20436;
   wire n20437;
   wire n20438;
   wire n20439;
   wire n20440;
   wire n20441;
   wire n20442;
   wire n20443;
   wire n20444;
   wire n20445;
   wire n20446;
   wire n20447;
   wire n20448;
   wire n20449;
   wire n20450;
   wire n20451;
   wire n20452;
   wire n20453;
   wire n20454;
   wire n20455;
   wire n20456;
   wire n20457;
   wire n20458;
   wire n20459;
   wire n20460;
   wire n20461;
   wire n20462;
   wire n20463;
   wire n20464;
   wire n20465;
   wire n20466;
   wire n20467;
   wire n20468;
   wire n20469;
   wire n20470;
   wire n20471;
   wire n20472;
   wire n20473;
   wire n20474;
   wire n20475;
   wire n20476;
   wire n20477;
   wire n20478;
   wire n20479;
   wire n20480;
   wire n20481;
   wire n20482;
   wire n20483;
   wire n20484;
   wire n20485;
   wire n20486;
   wire n20487;
   wire n20488;
   wire n20489;
   wire n20490;
   wire n20491;
   wire n20492;
   wire n20493;
   wire n20494;
   wire n20495;
   wire n20496;
   wire n20497;
   wire n20498;
   wire n20499;
   wire n20500;
   wire n20501;
   wire n20502;
   wire n20503;
   wire n20504;
   wire n20505;
   wire n20506;
   wire n20507;
   wire n20508;
   wire n20509;
   wire n20510;
   wire n20511;
   wire n20512;
   wire n20513;
   wire n20514;
   wire n20515;
   wire n20516;
   wire n20517;
   wire n20518;
   wire n20519;
   wire n20520;
   wire n20521;
   wire n20522;
   wire n20523;
   wire n20524;
   wire n20525;
   wire n20526;
   wire n20527;
   wire n20528;
   wire n20529;
   wire n20530;
   wire n20531;
   wire n20532;
   wire n20533;
   wire n20534;
   wire n20535;
   wire n20536;
   wire n20537;
   wire n20538;
   wire n20539;
   wire n20540;
   wire n20541;
   wire n20542;
   wire n20543;
   wire n20544;
   wire n20545;
   wire n20546;
   wire n20547;
   wire n20548;
   wire n20549;
   wire n20550;
   wire n20551;
   wire n20552;
   wire n20553;
   wire n20554;
   wire n20555;
   wire n20556;
   wire n20557;
   wire n20558;
   wire n20559;
   wire n20560;
   wire n20561;
   wire n20562;
   wire n20563;
   wire n20564;
   wire n20565;
   wire n20566;
   wire n20567;
   wire n20568;
   wire n20569;
   wire n20570;
   wire n20571;
   wire n20572;
   wire n20573;
   wire n20574;
   wire n20575;
   wire n20576;
   wire n20577;
   wire n20578;
   wire n20579;
   wire n20580;
   wire n20581;
   wire n20582;
   wire n20583;
   wire n20584;
   wire n20585;
   wire n20586;
   wire n20587;
   wire n20588;
   wire n20589;
   wire n20590;
   wire n20591;
   wire n20592;
   wire n20593;
   wire n20594;
   wire n20595;
   wire n20596;
   wire n20597;
   wire n20598;
   wire n20599;
   wire n20600;
   wire n20601;
   wire n20602;
   wire n20603;
   wire n20604;
   wire n20605;
   wire n20606;
   wire n20607;
   wire n20608;
   wire n20609;
   wire n20610;
   wire n20611;
   wire n20612;
   wire n20613;
   wire n20614;
   wire n20615;
   wire n20616;
   wire n20617;
   wire n20618;
   wire n20619;
   wire n20620;
   wire n20621;
   wire n20622;
   wire n20623;
   wire n20624;
   wire n20625;
   wire n20626;
   wire n20627;
   wire n20628;
   wire n20629;
   wire n20630;
   wire n20631;
   wire n20632;
   wire n20633;
   wire n20634;
   wire n20635;
   wire n20636;
   wire n20637;
   wire n20638;
   wire n20639;
   wire n20640;
   wire n20641;
   wire n20642;
   wire n20643;
   wire n20644;
   wire n20645;
   wire n20646;
   wire n20647;
   wire n20648;
   wire n20649;
   wire n20650;
   wire n20651;
   wire n20652;
   wire n20653;
   wire n20654;
   wire n20655;
   wire n20656;
   wire n20657;
   wire n20658;
   wire n20659;
   wire n20660;
   wire n20661;
   wire n20662;
   wire n20663;
   wire n20664;
   wire n20665;
   wire n20666;
   wire n20667;
   wire n20668;
   wire n20669;
   wire n20670;
   wire n20671;
   wire n20672;
   wire n20673;
   wire n20674;
   wire n20675;
   wire n20676;
   wire n20677;
   wire n20678;
   wire n20679;
   wire n20680;
   wire n20681;
   wire n20682;
   wire n20683;
   wire n20684;
   wire n20685;
   wire n20686;
   wire n20687;
   wire n20688;
   wire n20689;
   wire n20690;
   wire n20691;
   wire n20692;
   wire n20693;
   wire n20694;
   wire n20695;
   wire n20696;
   wire n20697;
   wire n20698;
   wire n20699;
   wire n20700;
   wire n20701;
   wire n20702;
   wire n20703;
   wire n20704;
   wire n20705;
   wire n20706;
   wire n20707;
   wire n20708;
   wire n20709;
   wire n20710;
   wire n20711;
   wire n20712;
   wire n20713;
   wire n20714;
   wire n20715;
   wire n20716;
   wire n20717;
   wire n20718;
   wire n20719;
   wire n20720;
   wire n20721;
   wire n20722;
   wire n20723;
   wire n20724;
   wire n20725;
   wire n20726;
   wire n20727;
   wire n20728;
   wire n20729;
   wire n20730;
   wire n20731;
   wire n20732;
   wire n20733;
   wire n20734;
   wire n20735;
   wire n20736;
   wire n20737;
   wire n20738;
   wire n20739;
   wire n20740;
   wire n20741;
   wire n20742;
   wire n20743;
   wire n20744;
   wire n20745;
   wire n20746;
   wire n20747;
   wire n20748;
   wire n20749;
   wire n20750;
   wire n20751;
   wire n20752;
   wire n20753;
   wire n20754;
   wire n20755;
   wire n20756;
   wire n20757;
   wire n20758;
   wire n20759;
   wire n20760;
   wire n20761;
   wire n20762;
   wire n20763;
   wire n20764;
   wire n20765;
   wire n20766;
   wire n20767;
   wire n20768;
   wire n20769;
   wire n20770;
   wire n20771;
   wire n20772;
   wire n20773;
   wire n20774;
   wire n20775;
   wire n20776;
   wire n20777;
   wire n20778;
   wire n20779;
   wire n20780;
   wire n20781;
   wire n20782;
   wire n20783;
   wire n20784;
   wire n20785;
   wire n20786;
   wire n20787;
   wire n20788;
   wire n20789;
   wire n20790;
   wire n20791;
   wire n20792;
   wire n20793;
   wire n20794;
   wire n20795;
   wire n20796;
   wire n20797;
   wire n20798;
   wire n20799;
   wire n20800;
   wire n20801;
   wire n20802;
   wire n20803;
   wire n20804;
   wire n20805;
   wire n20806;
   wire n20807;
   wire n20808;
   wire n20809;
   wire n20810;
   wire n20811;
   wire n20812;
   wire n20813;
   wire n20814;
   wire n20815;
   wire n20816;
   wire n20817;
   wire n20818;
   wire n20819;
   wire n20820;
   wire n20821;
   wire n20822;
   wire n20823;
   wire n20824;
   wire n20825;
   wire n20826;
   wire n20827;
   wire n20828;
   wire n20829;
   wire n20830;
   wire n20831;
   wire n20832;
   wire n20833;
   wire n20834;
   wire n20835;
   wire n20836;
   wire n20837;
   wire n20838;
   wire n20839;
   wire n20840;
   wire n20841;
   wire n20842;
   wire n20843;
   wire n20844;
   wire n20845;
   wire n20846;
   wire n20847;
   wire n20848;
   wire n20849;
   wire n20850;
   wire n20851;
   wire n20852;
   wire n20853;
   wire n20854;
   wire n20855;
   wire n20856;
   wire n20857;
   wire n20858;
   wire n20860;
   wire n20861;
   wire n20862;
   wire n20863;
   wire n20864;
   wire n20865;
   wire n20866;
   wire n20867;
   wire n20868;
   wire n20869;
   wire n20870;
   wire n20871;
   wire n20872;
   wire n20873;
   wire n20874;
   wire n20875;
   wire n20876;
   wire n20877;
   wire n20878;
   wire n20879;
   wire n20880;
   wire n20881;
   wire n20882;
   wire n20883;
   wire n20884;
   wire n20885;
   wire n20886;
   wire n20887;
   wire n20888;
   wire n20889;
   wire n20890;
   wire n20891;
   wire n20892;
   wire n20893;
   wire n20894;
   wire n20895;
   wire n20896;
   wire n20897;
   wire n20898;
   wire n20899;
   wire n20900;
   wire n20901;
   wire n20902;
   wire n20903;
   wire n20904;
   wire n20905;
   wire n20906;
   wire n20907;
   wire n20908;
   wire n20909;
   wire n20910;
   wire n20911;
   wire n20912;
   wire n20913;
   wire n20914;
   wire n20915;
   wire n20916;
   wire n20917;
   wire n20918;
   wire n20919;
   wire n20920;
   wire n20921;
   wire n20922;
   wire n20923;
   wire n20924;
   wire n20925;
   wire n20926;
   wire n20927;
   wire n20928;
   wire n20929;
   wire n20930;
   wire n20931;
   wire n20932;
   wire n20933;
   wire n20934;
   wire n20935;
   wire n20936;
   wire n20937;
   wire n20938;
   wire n20939;
   wire n20940;
   wire n20941;
   wire n20942;
   wire n20943;
   wire n20944;
   wire n20945;
   wire n20946;
   wire n20947;
   wire n20948;
   wire n20949;
   wire n20950;
   wire n20951;
   wire n20952;
   wire n20953;
   wire n20954;
   wire n20955;
   wire n20956;
   wire n20957;
   wire n20958;
   wire n20959;
   wire n20960;
   wire n20961;
   wire n20962;
   wire n20963;
   wire n20964;
   wire n20965;
   wire n20966;
   wire n20967;
   wire n20968;
   wire n20969;
   wire n20970;
   wire n20971;
   wire n20972;
   wire n20973;
   wire n20974;
   wire n20975;
   wire n20976;
   wire n20977;
   wire n20978;
   wire n20979;
   wire n20980;
   wire n20981;
   wire n20982;
   wire n20983;
   wire n20984;
   wire n20985;
   wire n20986;
   wire n20987;
   wire n20988;
   wire n20989;
   wire n20990;
   wire n20991;
   wire n20992;
   wire n20993;
   wire n20994;
   wire n20995;
   wire n20996;
   wire n20997;
   wire n20998;
   wire n20999;
   wire n21000;
   wire n21001;
   wire n21002;
   wire n21003;
   wire n21004;
   wire n21005;
   wire n21006;
   wire n21007;
   wire n21008;
   wire n21009;
   wire n21010;
   wire n21011;
   wire n21012;
   wire n21013;
   wire n21014;
   wire n21015;
   wire n21016;
   wire n21017;
   wire n21018;
   wire n21019;
   wire n21020;
   wire n21021;
   wire n21022;
   wire n21023;
   wire n21024;
   wire n21025;
   wire n21026;
   wire n21027;
   wire n21028;
   wire n21029;
   wire n21030;
   wire n21031;
   wire n21032;
   wire n21033;
   wire n21034;
   wire n21035;
   wire n21036;
   wire n21037;
   wire n21038;
   wire n21039;
   wire n21040;
   wire n21041;
   wire n21042;
   wire n21043;
   wire n21044;
   wire n21045;
   wire n21046;
   wire n21047;
   wire n21048;
   wire n21049;
   wire n21050;
   wire n21051;
   wire n21052;
   wire n21053;
   wire n21054;
   wire n21055;
   wire n21056;
   wire n21057;
   wire n21058;
   wire n21059;
   wire n21060;
   wire n21061;
   wire n21062;
   wire n21063;
   wire n21064;
   wire n21065;
   wire n21066;
   wire n21067;
   wire n21068;
   wire n21069;
   wire n21070;
   wire n21071;
   wire n21072;
   wire n21073;
   wire n21074;
   wire n21075;
   wire n21076;
   wire n21077;
   wire n21078;
   wire n21079;
   wire n21080;
   wire n21081;
   wire n21082;
   wire n21083;
   wire n21084;
   wire n21085;
   wire n21086;
   wire n21087;
   wire n21088;
   wire n21089;
   wire n21090;
   wire n21091;
   wire n21092;
   wire n21093;
   wire n21094;
   wire n21095;
   wire n21096;
   wire n21097;
   wire n21098;
   wire n21099;
   wire n21100;
   wire n21101;
   wire n21102;
   wire n21103;
   wire n21104;
   wire n21105;
   wire n21106;
   wire n21107;
   wire n21108;
   wire n21109;
   wire n21110;
   wire n21111;
   wire n21112;
   wire n21113;
   wire n21114;
   wire n21115;
   wire n21116;
   wire n21117;
   wire n21118;
   wire n21119;
   wire n21120;
   wire n21121;
   wire n21122;
   wire n21123;
   wire n21124;
   wire n21125;
   wire n21126;
   wire n21127;
   wire n21128;
   wire n21129;
   wire n21130;
   wire n21131;
   wire n21132;
   wire n21133;
   wire n21134;
   wire n21135;
   wire n21136;
   wire n21137;
   wire n21138;
   wire n21139;
   wire n21140;
   wire n21141;
   wire n21142;
   wire n21143;
   wire n21144;
   wire n21145;
   wire n21146;
   wire n21147;
   wire n21148;
   wire n21149;
   wire n21150;
   wire n21151;
   wire n21152;
   wire n21153;
   wire n21154;
   wire n21155;
   wire n21156;
   wire n21157;
   wire n21158;
   wire n21159;
   wire n21160;
   wire n21161;
   wire n21162;
   wire n21163;
   wire n21164;
   wire n21165;
   wire n21166;
   wire n21167;
   wire n21168;
   wire n21169;
   wire n21170;
   wire n21171;
   wire n21172;
   wire n21173;
   wire n21174;
   wire n21175;
   wire n21176;
   wire n21177;
   wire n21178;
   wire n21179;
   wire n21180;
   wire n21181;
   wire n21182;
   wire n21183;
   wire n21184;
   wire n21185;
   wire n21186;
   wire n21187;
   wire n21188;
   wire n21189;
   wire n21190;
   wire n21191;
   wire n21192;
   wire n21193;
   wire n21194;
   wire n21195;
   wire n21196;
   wire n21197;
   wire n21198;
   wire n21199;
   wire n21200;
   wire n21201;
   wire n21202;
   wire n21203;
   wire n21204;
   wire n21205;
   wire n21206;
   wire n21207;
   wire n21208;
   wire n21209;
   wire n21210;
   wire n21211;
   wire n21212;
   wire n21213;
   wire n21214;
   wire n21215;
   wire n21216;
   wire n21217;
   wire n21218;
   wire n21219;
   wire n21220;
   wire n21221;
   wire n21222;
   wire n21223;
   wire n21224;
   wire n21225;
   wire n21226;
   wire n21227;
   wire n21228;
   wire n21229;
   wire n21230;
   wire n21231;
   wire n21232;
   wire n21233;
   wire n21234;
   wire n21235;
   wire n21236;
   wire n21237;
   wire n21238;
   wire n21239;
   wire n21240;
   wire n21241;
   wire n21242;
   wire n21243;
   wire n21244;
   wire n21245;
   wire n21246;
   wire n21247;
   wire n21248;
   wire n21249;
   wire n21250;
   wire n21251;
   wire n21252;
   wire n21253;
   wire n21254;
   wire n21255;
   wire n21256;
   wire n21257;
   wire n21258;
   wire n21259;
   wire n21260;
   wire n21261;
   wire n21262;
   wire n21263;
   wire n21264;
   wire n21265;
   wire n21266;
   wire n21267;
   wire n21268;
   wire n21269;
   wire n21270;
   wire n21271;
   wire n21272;
   wire n21273;
   wire n21274;
   wire n21275;
   wire n21276;
   wire n21277;
   wire n21278;
   wire n21279;
   wire n21280;
   wire n21281;
   wire n21282;
   wire n21283;
   wire n21284;
   wire n21285;
   wire n21286;
   wire n21287;
   wire n21288;
   wire n21289;
   wire n21290;
   wire n21291;
   wire n21292;
   wire n21293;
   wire n21294;
   wire n21295;
   wire n21296;
   wire n21297;
   wire n21298;
   wire n21299;
   wire n21300;
   wire n21301;
   wire n21302;
   wire n21303;
   wire n21304;
   wire n21305;
   wire n21306;
   wire n21307;
   wire n21308;
   wire n21309;
   wire n21310;
   wire n21311;
   wire n21312;
   wire n21313;
   wire n21314;
   wire n21315;
   wire n21316;
   wire n21317;
   wire n21318;
   wire n21319;
   wire n21320;
   wire n21321;
   wire n21322;
   wire n21323;
   wire n21324;
   wire n21325;
   wire n21326;
   wire n21327;
   wire n21328;
   wire n21329;
   wire n21330;
   wire n21331;
   wire n21332;
   wire n21333;
   wire n21334;
   wire n21335;
   wire n21336;
   wire n21337;
   wire n21338;
   wire n21339;
   wire n21340;
   wire n21341;
   wire n21342;
   wire n21343;
   wire n21344;
   wire n21345;
   wire n21346;
   wire n21347;
   wire n21348;
   wire n21349;
   wire n21350;
   wire n21351;
   wire n21352;
   wire n21353;
   wire n21354;
   wire n21355;
   wire n21356;
   wire n21357;
   wire n21358;
   wire n21359;
   wire n21360;
   wire n21361;
   wire n21362;
   wire n21363;
   wire n21364;
   wire n21365;
   wire n21366;
   wire n21367;
   wire n21368;
   wire n21369;
   wire n21370;
   wire n21371;
   wire n21372;
   wire n21373;
   wire n21374;
   wire n21375;
   wire n21376;
   wire n21377;
   wire n21378;
   wire n21379;
   wire n21380;
   wire n21381;
   wire n21382;
   wire n21383;
   wire n21384;
   wire n21385;
   wire n21386;
   wire n21387;
   wire n21388;
   wire n21389;
   wire n21390;
   wire n21391;
   wire n21392;
   wire n21393;
   wire n21394;
   wire n21395;
   wire n21396;
   wire n21397;
   wire n21398;
   wire n21399;
   wire n21400;
   wire n21401;
   wire n21402;
   wire n21403;
   wire n21404;
   wire n21405;
   wire n21406;
   wire n21407;
   wire n21408;
   wire n21409;
   wire n21410;
   wire n21411;
   wire n21412;
   wire n21413;
   wire n21414;
   wire n21415;
   wire n21416;
   wire n21417;
   wire n21418;
   wire n21419;
   wire n21420;
   wire n21421;
   wire n21422;
   wire n21423;
   wire n21424;
   wire n21425;
   wire n21426;
   wire n21427;
   wire n21428;
   wire n21429;
   wire n21430;
   wire n21431;
   wire n21432;
   wire n21433;
   wire n21434;
   wire n21435;
   wire n21436;
   wire n21437;
   wire n21438;
   wire n21439;
   wire n21440;
   wire n21441;
   wire n21442;
   wire n21443;
   wire n21444;
   wire n21445;
   wire n21446;
   wire n21447;
   wire n21448;
   wire n21449;
   wire n21450;
   wire n21451;
   wire n21452;
   wire n21453;
   wire n21454;
   wire n21455;
   wire n21456;
   wire n21457;
   wire n21458;
   wire n21459;
   wire n21460;
   wire n21461;
   wire n21462;
   wire n21463;
   wire n21464;
   wire n21465;
   wire n21466;
   wire n21467;
   wire n21468;
   wire n21469;
   wire n21470;
   wire n21471;
   wire n21472;
   wire n21473;
   wire n21474;
   wire n21475;
   wire n21476;
   wire n21477;
   wire n21478;
   wire n21479;
   wire n21480;
   wire n21481;
   wire n21482;
   wire n21483;
   wire n21484;
   wire n21485;
   wire n21486;
   wire n21487;
   wire n21488;
   wire n21489;
   wire n21490;
   wire n21491;
   wire n21492;
   wire n21493;
   wire n21494;
   wire n21495;
   wire n21496;
   wire n21497;
   wire n21498;
   wire n21499;
   wire n21500;
   wire n21501;
   wire n21502;
   wire n21503;
   wire n21504;
   wire n21505;
   wire n21506;
   wire n21507;
   wire n21508;
   wire n21509;
   wire n21510;
   wire n21511;
   wire n21512;
   wire n21513;
   wire n21514;
   wire n21515;
   wire n21516;
   wire n21517;
   wire n21518;
   wire n21519;
   wire n21520;
   wire n21521;
   wire n21522;
   wire n21523;
   wire n21524;
   wire n21525;
   wire n21526;
   wire n21527;
   wire n21528;
   wire n21529;
   wire n21530;
   wire n21531;
   wire n21532;
   wire n21533;
   wire n21534;
   wire n21535;
   wire n21536;
   wire n21537;
   wire n21538;
   wire n21539;
   wire n21540;
   wire n21541;
   wire n21542;
   wire n21543;
   wire n21544;
   wire n21545;
   wire n21546;
   wire n21547;
   wire n21548;
   wire n21549;
   wire n21550;
   wire n21551;
   wire n21552;
   wire n21553;
   wire n21554;
   wire n21555;
   wire n21556;
   wire n21557;
   wire n21558;
   wire n21559;
   wire n21560;
   wire n21561;
   wire n21562;
   wire n21563;
   wire n21564;
   wire n21565;
   wire n21566;
   wire n21567;
   wire n21568;
   wire n21569;
   wire n21570;
   wire n21571;
   wire n21572;
   wire n21573;
   wire n21574;
   wire n21575;
   wire n21576;
   wire n21577;
   wire n21578;
   wire n21579;
   wire n21580;
   wire n21581;
   wire n21582;
   wire n21583;
   wire n21584;
   wire n21585;
   wire n21586;
   wire n21587;
   wire n21588;
   wire n21589;
   wire n21590;
   wire n21591;
   wire n21592;
   wire n21593;
   wire n21594;
   wire n21595;
   wire n21596;
   wire n21597;
   wire n21598;
   wire n21599;
   wire n21600;
   wire n21601;
   wire n21602;
   wire n21603;
   wire n21604;
   wire n21605;
   wire n21606;
   wire n21607;
   wire n21608;
   wire n21609;
   wire n21610;
   wire n21611;
   wire n21612;
   wire n21613;
   wire n21614;
   wire n21615;
   wire n21616;
   wire n21617;
   wire n21618;
   wire n21619;
   wire n21620;
   wire n21621;
   wire n21622;
   wire n21623;
   wire n21624;
   wire n21625;
   wire n21626;
   wire n21627;
   wire n21628;
   wire n21629;
   wire n21630;
   wire n21631;
   wire n21632;
   wire n21633;
   wire n21634;
   wire n21635;
   wire n21636;
   wire n21637;
   wire n21638;
   wire n21639;
   wire n21640;
   wire n21641;
   wire n21643;
   wire n21644;
   wire n21645;
   wire n21647;
   wire n21648;
   wire n21649;
   wire n21650;
   wire n21651;
   wire n21652;
   wire n21653;
   wire n21654;
   wire n21655;
   wire n21656;
   wire n21657;
   wire n21658;
   wire n21659;
   wire n21660;
   wire n21661;
   wire n21662;
   wire n21663;
   wire n21664;
   wire n21665;
   wire n21666;
   wire n21667;
   wire n21668;
   wire n21669;
   wire n21670;
   wire n21671;
   wire n21672;
   wire n21673;
   wire n21674;
   wire n21675;
   wire n21676;
   wire n21677;
   wire n21678;
   wire n21679;
   wire n21680;
   wire n21681;
   wire n21682;
   wire n21683;
   wire n21684;
   wire n21685;
   wire n21686;
   wire n21687;
   wire n21688;
   wire n21689;
   wire n21690;
   wire n21691;
   wire n21692;
   wire n21693;
   wire n21694;
   wire n21695;
   wire n21696;
   wire n21697;
   wire n21698;
   wire n21699;
   wire n21700;
   wire n21701;
   wire n21702;
   wire n21703;
   wire n21704;
   wire n21705;
   wire n21706;
   wire n21707;
   wire n21708;
   wire n21709;
   wire n21710;
   wire n21711;
   wire n21712;
   wire n21713;
   wire n21714;
   wire n21715;
   wire n21716;
   wire n21717;
   wire n21718;
   wire n21719;
   wire n21720;
   wire n21721;
   wire n21722;
   wire n21723;
   wire n21724;
   wire n21725;
   wire n21726;
   wire n21727;
   wire n21728;
   wire n21729;
   wire n21730;
   wire n21731;
   wire n21732;
   wire n21733;
   wire n21734;
   wire n21735;
   wire n21736;
   wire n21737;
   wire n21738;
   wire n21739;
   wire n21740;
   wire n21741;
   wire n21742;
   wire n21743;
   wire n21744;
   wire n21745;
   wire n21746;
   wire n21747;
   wire n21748;
   wire n21749;
   wire n21750;
   wire n21751;
   wire n21752;
   wire n21753;
   wire n21754;
   wire n21755;
   wire n21756;
   wire n21757;
   wire n21758;
   wire n21759;
   wire n21760;
   wire n21761;
   wire n21762;
   wire n21763;
   wire n21764;
   wire n21765;
   wire n21766;
   wire n21767;
   wire n21768;
   wire n21769;
   wire n21770;
   wire n21771;
   wire n21772;
   wire n21773;
   wire n21774;
   wire n21775;
   wire n21776;
   wire n21777;
   wire n21778;
   wire n21779;
   wire n21780;
   wire n21781;
   wire n21782;
   wire n21783;
   wire n21784;
   wire n21785;
   wire n21786;
   wire n21787;
   wire n21788;
   wire n21789;
   wire n21790;
   wire n21791;
   wire n21792;
   wire n21793;
   wire n21794;
   wire n21796;
   wire n21797;
   wire n21798;
   wire n21799;
   wire n21800;
   wire n21801;
   wire n21802;
   wire n21803;
   wire n21804;
   wire n21805;
   wire n21806;
   wire n21807;
   wire n21808;
   wire n21809;
   wire n21810;
   wire n21811;
   wire n21812;
   wire n21813;
   wire n21814;
   wire n21815;
   wire n21816;
   wire n21817;
   wire n21818;
   wire n21819;
   wire n21820;
   wire n21821;
   wire n21822;
   wire n21823;
   wire n21824;
   wire n21825;
   wire n21826;
   wire n21827;
   wire n21828;
   wire n21829;
   wire n21830;
   wire n21831;
   wire n21832;
   wire n21833;
   wire n21834;
   wire n21835;
   wire n21836;
   wire n21837;
   wire n21838;
   wire n21839;
   wire n21840;
   wire n21841;
   wire n21842;
   wire n21843;
   wire n21844;
   wire n21845;
   wire n21847;
   wire n21848;
   wire n21849;
   wire n21850;
   wire n21851;
   wire n21852;
   wire n21853;
   wire n21854;
   wire n21855;
   wire n21856;
   wire n21857;
   wire n21858;
   wire n21859;
   wire n21860;
   wire n21862;
   wire n21863;
   wire n21864;
   wire n21865;
   wire n21866;
   wire n21867;
   wire n21868;
   wire n21869;
   wire n21870;
   wire n21871;
   wire n21872;
   wire n21873;
   wire n21874;
   wire n21875;
   wire n21876;
   wire n21877;
   wire n21878;
   wire n21879;
   wire n21880;
   wire n21881;
   wire n21882;
   wire n21883;
   wire n21884;
   wire n21885;
   wire n21886;
   wire n21887;
   wire n21888;
   wire n21889;
   wire n21890;
   wire n21891;
   wire n21892;
   wire n21893;
   wire n21894;
   wire n21895;
   wire n21896;
   wire n21897;
   wire n21898;
   wire n21899;
   wire n21900;
   wire n21901;
   wire n21902;
   wire n21903;
   wire n21904;
   wire n21905;
   wire n21906;
   wire n21907;
   wire n21908;
   wire n21909;
   wire n21910;
   wire n21911;
   wire n21912;
   wire n21913;
   wire n21914;
   wire n21915;
   wire n21916;
   wire n21917;
   wire n21918;
   wire n21919;
   wire n21920;
   wire n21921;
   wire n21922;
   wire n21923;
   wire n21924;
   wire n21925;
   wire n21926;
   wire n21927;
   wire n21928;
   wire n21929;
   wire n21930;
   wire n21931;
   wire n21932;
   wire n21933;
   wire n21934;
   wire n21935;
   wire n21936;
   wire n21937;
   wire n21938;
   wire n21939;
   wire n21940;
   wire n21941;
   wire n21942;
   wire n21943;
   wire n21944;
   wire n21945;
   wire n21946;
   wire n21947;
   wire n21948;
   wire n21949;
   wire n21950;
   wire n21951;
   wire n21952;
   wire n21953;
   wire n21954;
   wire n21955;
   wire n21956;
   wire n21957;
   wire n21958;
   wire n21959;
   wire n21960;
   wire n21961;
   wire n21962;
   wire n21963;
   wire n21964;
   wire n21965;
   wire n21966;
   wire n21967;
   wire n21968;
   wire n21969;
   wire n21970;
   wire n21971;
   wire n21972;
   wire n21973;
   wire n21974;
   wire n21975;
   wire n21976;
   wire n21977;
   wire n21978;
   wire n21979;
   wire n21980;
   wire n21981;
   wire n21982;
   wire n21983;
   wire n21984;
   wire n21985;
   wire n21986;
   wire n21987;
   wire n21988;
   wire n21989;
   wire n21990;
   wire n21991;
   wire n21992;
   wire n21993;
   wire n21994;
   wire n21995;
   wire n21996;
   wire n21997;
   wire n21998;
   wire n21999;
   wire n22000;
   wire n22001;
   wire n22002;
   wire n22003;
   wire n22004;
   wire n22005;
   wire n22006;
   wire n22007;
   wire n22008;
   wire n22009;
   wire n22010;
   wire n22011;
   wire n22012;
   wire n22013;
   wire n22014;
   wire n22015;
   wire n22016;
   wire n22017;
   wire n22018;
   wire n22019;
   wire n22020;
   wire n22021;
   wire n22022;
   wire n22023;
   wire n22024;
   wire n22025;
   wire n22026;
   wire n22027;
   wire n22028;
   wire n22029;
   wire n22030;
   wire n22031;
   wire n22032;
   wire n22033;
   wire n22034;
   wire n22035;
   wire n22036;
   wire n22037;
   wire n22038;
   wire n22039;
   wire n22040;
   wire n22041;
   wire n22042;
   wire n22043;
   wire n22044;
   wire n22045;
   wire n22046;
   wire n22047;
   wire n22048;
   wire n22049;
   wire n22050;
   wire n22051;
   wire n22052;
   wire n22053;
   wire n22054;
   wire n22055;
   wire n22056;
   wire n22057;
   wire n22058;
   wire n22059;
   wire n22060;
   wire n22061;
   wire n22062;
   wire n22063;
   wire n22064;
   wire n22065;
   wire n22066;
   wire n22067;
   wire n22068;
   wire n22069;
   wire n22070;
   wire n22071;
   wire n22072;
   wire n22073;
   wire n22074;
   wire n22075;
   wire n22076;
   wire n22077;
   wire n22078;
   wire n22079;
   wire n22080;
   wire n22081;
   wire n22082;
   wire n22083;
   wire n22084;
   wire n22085;
   wire n22086;
   wire n22087;
   wire n22088;
   wire n22089;
   wire n22090;
   wire n22091;
   wire n22092;
   wire n22093;
   wire n22094;
   wire n22095;
   wire n22096;
   wire n22097;
   wire n22098;
   wire n22099;
   wire n22100;
   wire n22101;
   wire n22102;
   wire n22103;
   wire n22104;
   wire n22105;
   wire n22106;
   wire n22107;
   wire n22108;
   wire n22109;
   wire n22110;
   wire n22111;
   wire n22112;
   wire n22113;
   wire n22114;
   wire n22115;
   wire n22116;
   wire n22117;
   wire n22118;
   wire n22119;
   wire n22120;
   wire n22121;
   wire n22122;
   wire n22123;
   wire n22124;
   wire n22125;
   wire n22126;
   wire n22127;
   wire n22128;
   wire n22129;
   wire n22130;
   wire n22131;
   wire n22132;
   wire n22133;
   wire n22134;
   wire n22135;
   wire n22136;
   wire n22137;
   wire n22138;
   wire n22139;
   wire n22140;
   wire n22141;
   wire n22142;
   wire n22143;
   wire n22144;
   wire n22145;
   wire n22146;
   wire n22147;
   wire n22148;
   wire n22149;
   wire n22150;
   wire n22151;
   wire n22152;
   wire n22153;
   wire n22154;
   wire n22155;
   wire n22156;
   wire n22157;
   wire n22158;
   wire n22159;
   wire n22160;
   wire n22161;
   wire n22162;
   wire n22163;
   wire n22164;
   wire n22165;
   wire n22166;
   wire n22167;
   wire n22168;
   wire n22169;
   wire n22170;
   wire n22171;
   wire n22172;
   wire n22173;
   wire n22174;
   wire n22175;
   wire n22176;
   wire n22177;
   wire n22178;
   wire n22179;
   wire n22180;
   wire n22181;
   wire n22182;
   wire n22183;
   wire n22184;
   wire n22185;
   wire n22186;
   wire n22187;
   wire n22188;
   wire n22189;
   wire n22190;
   wire n22191;
   wire n22192;
   wire n22193;
   wire n22194;
   wire n22195;
   wire n22196;
   wire n22197;
   wire n22198;
   wire n22199;
   wire n22200;
   wire n22201;
   wire n22202;
   wire n22203;
   wire n22204;
   wire n22205;
   wire n22206;
   wire n22207;
   wire n22208;
   wire n22209;
   wire n22210;
   wire n22211;
   wire n22212;
   wire n22213;
   wire n22214;
   wire n22215;
   wire n22216;
   wire n22217;
   wire n22218;
   wire n22219;
   wire n22220;
   wire n22221;
   wire n22222;
   wire n22223;
   wire n22224;
   wire n22225;
   wire n22226;
   wire n22227;
   wire n22228;
   wire n22229;
   wire n22230;
   wire n22231;
   wire n22232;
   wire n22233;
   wire n22234;
   wire n22235;
   wire n22236;
   wire n22237;
   wire n22238;
   wire n22239;
   wire n22240;
   wire n22241;
   wire n22242;
   wire n22243;
   wire n22244;
   wire n22245;
   wire n22246;
   wire n22247;
   wire n22248;
   wire n22249;
   wire n22250;
   wire n22251;
   wire n22252;
   wire n22253;
   wire n22254;
   wire n22255;
   wire n22256;
   wire n22257;
   wire n22258;
   wire n22259;
   wire n22260;
   wire n22261;
   wire n22262;
   wire n22263;
   wire n22264;
   wire n22265;
   wire n22266;
   wire n22267;
   wire n22268;
   wire n22269;
   wire n22270;
   wire n22271;
   wire n22272;
   wire n22273;
   wire n22274;
   wire n22275;
   wire n22276;
   wire n22277;
   wire n22278;
   wire n22279;
   wire n22280;
   wire n22281;
   wire n22282;
   wire n22283;
   wire n22284;
   wire n22285;
   wire n22286;
   wire n22287;
   wire n22288;
   wire n22289;
   wire n22290;
   wire n22291;
   wire n22292;
   wire n22293;
   wire n22294;
   wire n22295;
   wire n22296;
   wire n22297;
   wire n22298;
   wire n22299;
   wire n22300;
   wire n22301;
   wire n22302;
   wire n22303;
   wire n22304;
   wire n22305;
   wire n22306;
   wire n22307;
   wire n22308;
   wire n22309;
   wire n22310;
   wire n22311;
   wire n22312;
   wire n22313;
   wire n22314;
   wire n22315;
   wire n22316;
   wire n22317;
   wire n22318;
   wire n22319;
   wire n22320;
   wire n22321;
   wire n22322;
   wire n22323;
   wire n22324;
   wire n22325;
   wire n22326;
   wire n22327;
   wire n22328;
   wire n22329;
   wire n22330;
   wire n22331;
   wire n22332;
   wire n22333;
   wire n22334;
   wire n22335;
   wire n22336;
   wire n22337;
   wire n22338;
   wire n22339;
   wire n22340;
   wire n22341;
   wire n22342;
   wire n22343;
   wire n22344;
   wire n22345;
   wire n22346;
   wire n22347;
   wire n22348;
   wire n22349;
   wire n22350;
   wire n22351;
   wire n22352;
   wire n22353;
   wire n22354;
   wire n22355;
   wire n22356;
   wire n22357;
   wire n22358;
   wire n22359;
   wire n22360;
   wire n22361;
   wire n22362;
   wire n22363;
   wire n22364;
   wire n22365;
   wire n22366;
   wire n22367;
   wire n22368;
   wire n22369;
   wire n22370;
   wire n22371;
   wire n22372;
   wire n22373;
   wire n22374;
   wire n22375;
   wire n22376;
   wire n22377;
   wire n22378;
   wire n22379;
   wire n22380;
   wire n22381;
   wire n22382;
   wire n22383;
   wire n22384;
   wire n22385;
   wire n22386;
   wire n22387;
   wire n22388;
   wire n22389;
   wire n22390;
   wire n22391;
   wire n22392;
   wire n22393;
   wire n22394;
   wire n22395;
   wire n22396;
   wire n22397;
   wire n22398;
   wire n22399;
   wire n22400;
   wire n22401;
   wire n22402;
   wire n22403;
   wire n22404;
   wire n22405;
   wire n22406;
   wire n22407;
   wire n22408;
   wire n22409;
   wire n22410;
   wire n22411;
   wire n22412;
   wire n22413;
   wire n22414;
   wire n22415;
   wire n22416;
   wire n22417;
   wire n22418;
   wire n22419;
   wire n22420;
   wire n22421;
   wire n22422;
   wire n22423;
   wire n22424;
   wire n22425;
   wire n22426;
   wire n22427;
   wire n22428;
   wire n22429;
   wire n22430;
   wire n22431;
   wire n22432;
   wire n22433;
   wire n22434;
   wire n22435;
   wire n22436;
   wire n22437;
   wire n22438;
   wire n22439;
   wire n22440;
   wire n22441;
   wire n22442;
   wire n22443;
   wire n22444;
   wire n22445;
   wire n22446;
   wire n22447;
   wire n22448;
   wire n22449;
   wire n22450;
   wire n22451;
   wire n22452;
   wire n22453;
   wire n22454;
   wire n22455;
   wire n22456;
   wire n22457;
   wire n22458;
   wire n22459;
   wire n22460;
   wire n22461;
   wire n22462;
   wire n22463;
   wire n22464;
   wire n22465;
   wire n22466;
   wire n22467;
   wire n22468;
   wire n22469;
   wire n22470;
   wire n22471;
   wire n22472;
   wire n22473;
   wire n22474;
   wire n22475;
   wire n22476;
   wire n22477;
   wire n22478;
   wire n22479;
   wire n22480;
   wire n22481;
   wire n22482;
   wire n22483;
   wire n22484;
   wire n22485;
   wire n22486;
   wire n22487;
   wire n22488;
   wire n22489;
   wire n22490;
   wire n22491;
   wire n22492;
   wire n22493;
   wire n22494;
   wire n22495;
   wire n22496;
   wire n22497;
   wire n22498;
   wire n22499;
   wire n22500;
   wire n22501;
   wire n22502;
   wire n22503;
   wire n22504;
   wire n22505;
   wire n22506;
   wire n22507;
   wire n22508;
   wire n22509;
   wire n22510;
   wire n22511;
   wire n22512;
   wire n22513;
   wire n22514;
   wire n22515;
   wire n22516;
   wire n22517;
   wire n22518;
   wire n22519;
   wire n22520;
   wire n22521;
   wire n22522;
   wire n22523;
   wire n22524;
   wire n22525;
   wire n22526;
   wire n22527;
   wire n22528;
   wire n22529;
   wire n22530;
   wire n22531;
   wire n22532;
   wire n22533;
   wire n22534;
   wire n22535;
   wire n22536;
   wire n22537;
   wire n22538;
   wire n22539;
   wire n22540;
   wire n22541;
   wire n22542;
   wire n22543;
   wire n22544;
   wire n22545;
   wire n22546;
   wire n22547;
   wire n22548;
   wire n22549;
   wire n22550;
   wire n22551;
   wire n22552;
   wire n22553;
   wire n22554;
   wire n22555;
   wire n22556;
   wire n22557;
   wire n22558;
   wire n22559;
   wire n22560;
   wire n22561;
   wire n22562;
   wire n22563;
   wire n22564;
   wire n22565;
   wire n22566;
   wire n22567;
   wire n22568;
   wire n22569;
   wire n22570;
   wire n22571;
   wire n22572;
   wire n22573;
   wire n22574;
   wire n22575;
   wire n22576;
   wire n22577;
   wire n22578;
   wire n22579;
   wire n22580;
   wire n22581;
   wire n22582;
   wire n22583;
   wire n22584;
   wire n22585;
   wire n22586;
   wire n22587;
   wire n22588;
   wire n22589;
   wire n22590;
   wire n22591;
   wire n22592;
   wire n22593;
   wire n22594;
   wire n22595;
   wire n22596;
   wire n22597;
   wire n22598;
   wire n22599;
   wire n22600;
   wire n22601;
   wire n22602;
   wire n22603;
   wire n22604;
   wire n22605;
   wire n22606;
   wire n22607;
   wire n22608;
   wire n22609;
   wire n22610;
   wire n22611;
   wire n22612;
   wire n22613;
   wire n22614;
   wire n22615;
   wire n22616;
   wire n22617;
   wire n22618;
   wire n22619;
   wire n22620;
   wire n22621;
   wire n22622;
   wire n22623;
   wire n22624;
   wire n22625;
   wire n22626;
   wire n22627;
   wire n22628;
   wire n22629;
   wire n22630;
   wire n22631;
   wire n22632;
   wire n22633;
   wire n22634;
   wire n22635;
   wire n22636;
   wire n22637;
   wire n22638;
   wire n22639;
   wire n22640;
   wire n22641;
   wire n22642;
   wire n22643;
   wire n22644;
   wire n22645;
   wire n22646;
   wire n22647;
   wire n22648;
   wire n22649;
   wire n22650;
   wire n22651;
   wire n22652;
   wire n22653;
   wire n22654;
   wire n22655;
   wire n22656;
   wire n22657;
   wire n22658;
   wire n22659;
   wire n22660;
   wire n22661;
   wire n22662;
   wire n22663;
   wire n22664;
   wire n22665;
   wire n22666;
   wire n22667;
   wire n22668;
   wire n22669;
   wire n22670;
   wire n22671;
   wire n22672;
   wire n22673;
   wire n22674;
   wire n22675;
   wire n22676;
   wire n22677;
   wire n22678;
   wire n22679;
   wire n22680;
   wire n22681;
   wire n22682;
   wire n22683;
   wire n22684;
   wire n22685;
   wire n22686;
   wire n22687;
   wire n22688;
   wire n22689;
   wire n22690;
   wire n22691;
   wire n22692;
   wire n22693;
   wire n22694;
   wire n22695;
   wire n22696;
   wire n22697;
   wire n22698;
   wire n22699;
   wire n22700;
   wire n22701;
   wire n22702;
   wire n22703;
   wire n22704;
   wire n22705;
   wire n22706;
   wire n22707;
   wire n22708;
   wire n22709;
   wire n22710;
   wire n22711;
   wire n22712;
   wire n22713;
   wire n22714;
   wire n22715;
   wire n22716;
   wire n22717;
   wire n22718;
   wire n22719;
   wire n22720;
   wire n22721;
   wire n22722;
   wire n22723;
   wire n22724;
   wire n22725;
   wire n22726;
   wire n22727;
   wire n22728;
   wire n22729;
   wire n22730;
   wire n22731;
   wire n22732;
   wire n22733;
   wire n22734;
   wire n22735;
   wire n22736;
   wire n22737;
   wire n22738;
   wire n22739;
   wire n22740;
   wire n22741;
   wire n22742;
   wire n22743;
   wire n22744;
   wire n22745;
   wire n22746;
   wire n22747;
   wire n22748;
   wire n22749;
   wire n22750;
   wire n22751;
   wire n22752;
   wire n22753;
   wire n22754;
   wire n22755;
   wire n22756;
   wire n22757;
   wire n22758;
   wire n22759;
   wire n22760;
   wire n22761;
   wire n22762;
   wire n22763;
   wire n22764;
   wire n22765;
   wire n22766;
   wire n22767;
   wire n22768;
   wire n22769;
   wire n22770;
   wire n22771;
   wire n22772;
   wire n22773;
   wire n22774;
   wire n22775;
   wire n22776;
   wire n22777;
   wire n22778;
   wire n22779;
   wire n22780;
   wire n22781;
   wire n22782;
   wire n22783;
   wire n22784;
   wire n22785;
   wire n22786;
   wire n22787;
   wire n22788;
   wire n22789;
   wire n22790;
   wire n22791;
   wire n22792;
   wire n22793;
   wire n22794;
   wire n22795;
   wire n22796;
   wire n22797;
   wire n22798;
   wire n22799;
   wire n22800;
   wire n22801;
   wire n22802;
   wire n22803;
   wire n22804;
   wire n22805;
   wire n22806;
   wire n22807;
   wire n22808;
   wire n22809;
   wire n22810;
   wire n22811;
   wire n22812;
   wire n22813;
   wire n22814;
   wire n22815;
   wire n22816;
   wire n22817;
   wire n22818;
   wire n22819;
   wire n22820;
   wire n22821;
   wire n22822;
   wire n22823;
   wire n22824;
   wire n22825;
   wire n22826;
   wire n22827;
   wire n22828;
   wire n22829;
   wire n22830;
   wire n22831;
   wire n22832;
   wire n22833;
   wire n22834;
   wire n22835;
   wire n22836;
   wire n22837;
   wire n22838;
   wire n22839;
   wire n22840;
   wire n22841;
   wire n22842;
   wire n22843;
   wire n22844;
   wire n22845;
   wire n22846;
   wire n22847;
   wire n22848;
   wire n22849;
   wire n22850;
   wire n22851;
   wire n22852;
   wire n22853;
   wire n22854;
   wire n22855;
   wire n22856;
   wire n22857;
   wire n22858;
   wire n22859;
   wire n22860;
   wire n22861;
   wire n22862;
   wire n22863;
   wire n22864;
   wire n22865;
   wire n22866;
   wire n22867;
   wire n22868;
   wire n22869;
   wire n22870;
   wire n22871;
   wire n22872;
   wire n22873;
   wire n22874;
   wire n22875;
   wire n22876;
   wire n22877;
   wire n22878;
   wire n22879;
   wire n22880;
   wire n22881;
   wire n22882;
   wire n22883;
   wire n22884;
   wire n22885;
   wire n22886;
   wire n22887;
   wire n22888;
   wire n22889;
   wire n22890;
   wire n22891;
   wire n22892;
   wire n22893;
   wire n22894;
   wire n22895;
   wire n22896;
   wire n22897;
   wire n22898;
   wire n22899;
   wire n22900;
   wire n22901;
   wire n22902;
   wire n22903;
   wire n22904;
   wire n22905;
   wire n22906;
   wire n22907;
   wire n22908;
   wire n22909;
   wire n22910;
   wire n22911;
   wire n22912;
   wire n22913;
   wire n22914;
   wire n22915;
   wire n22916;
   wire n22917;
   wire n22918;
   wire n22919;
   wire n22920;
   wire n22921;
   wire n22922;
   wire n22923;
   wire n22924;
   wire n22925;
   wire n22926;
   wire n22927;
   wire n22928;
   wire n22929;
   wire n22930;
   wire n22931;
   wire n22932;
   wire n22933;
   wire n22934;
   wire n22935;
   wire n22936;
   wire n22937;
   wire n22938;
   wire n22939;
   wire n22940;
   wire n22941;
   wire n22942;
   wire n22943;
   wire n22944;
   wire n22945;
   wire n22946;
   wire n22947;
   wire n22948;
   wire n22949;
   wire n22950;
   wire n22951;
   wire n22952;
   wire n22953;
   wire n22954;
   wire n22955;
   wire n22956;
   wire n22957;
   wire n22958;
   wire n22959;
   wire n22960;
   wire n22961;
   wire n22962;
   wire n22963;
   wire n22964;
   wire n22965;
   wire n22966;
   wire n22967;
   wire n22968;
   wire n22969;
   wire n22970;
   wire n22971;
   wire n22972;
   wire n22973;
   wire n22974;
   wire n22975;
   wire n22976;
   wire n22977;
   wire n22978;
   wire n22979;
   wire n22980;
   wire n22981;
   wire n22982;
   wire n22983;
   wire n22984;
   wire n22985;
   wire n22986;
   wire n22987;
   wire n22988;
   wire n22989;
   wire n22990;
   wire n22991;
   wire n22992;
   wire n22993;
   wire n22994;
   wire n22995;
   wire n22996;
   wire n22997;
   wire n22998;
   wire n22999;
   wire n23000;
   wire n23001;
   wire n23002;
   wire n23003;
   wire n23004;
   wire n23005;
   wire n23006;
   wire n23007;
   wire n23008;
   wire n23009;
   wire n23010;
   wire n23011;
   wire n23012;
   wire n23013;
   wire n23014;
   wire n23015;
   wire n23016;
   wire n23017;
   wire n23018;
   wire n23019;
   wire n23020;
   wire n23021;
   wire n23022;
   wire n23023;
   wire n23024;
   wire n23025;
   wire n23026;
   wire n23027;
   wire n23028;
   wire n23029;
   wire n23030;
   wire n23031;
   wire n23032;
   wire n23033;
   wire n23034;
   wire n23035;
   wire n23036;
   wire n23037;
   wire n23038;
   wire n23039;
   wire n23040;
   wire n23041;
   wire n23042;
   wire n23043;
   wire n23044;
   wire n23045;
   wire n23046;
   wire n23047;
   wire n23048;
   wire n23049;
   wire n23050;
   wire n23051;
   wire n23052;
   wire n23053;
   wire n23054;
   wire n23055;
   wire n23056;
   wire n23057;
   wire n23058;
   wire n23059;
   wire n23060;
   wire n23061;
   wire n23062;
   wire n23063;
   wire n23064;
   wire n23065;
   wire n23066;
   wire n23067;
   wire n23068;
   wire n23069;
   wire n23070;
   wire n23071;
   wire n23072;
   wire n23073;
   wire n23074;
   wire n23075;
   wire n23076;
   wire n23077;
   wire n23078;
   wire n23079;
   wire n23080;
   wire n23081;
   wire n23082;
   wire n23083;
   wire n23084;
   wire n23085;
   wire n23086;
   wire n23087;
   wire n23088;
   wire n23089;
   wire n23090;
   wire n23091;
   wire n23092;
   wire n23093;
   wire n23094;
   wire n23095;
   wire n23096;
   wire n23097;
   wire n23098;
   wire n23099;
   wire n23100;
   wire n23101;
   wire n23102;
   wire n23103;
   wire n23104;
   wire n23105;
   wire n23106;
   wire n23107;
   wire n23108;
   wire n23109;
   wire n23110;
   wire n23111;
   wire n23112;
   wire n23113;
   wire n23114;
   wire n23115;
   wire n23116;
   wire n23117;
   wire n23118;
   wire n23119;
   wire n23120;
   wire n23121;
   wire n23122;
   wire n23123;
   wire n23124;
   wire n23125;
   wire n23126;
   wire n23127;
   wire n23128;
   wire n23129;
   wire n23130;
   wire n23131;
   wire n23132;
   wire n23133;
   wire n23134;
   wire n23135;
   wire n23136;
   wire n23137;
   wire n23138;
   wire n23139;
   wire n23140;
   wire n23141;
   wire n23142;
   wire n23143;
   wire n23144;
   wire n23145;
   wire n23146;
   wire n23147;
   wire n23148;
   wire n23149;
   wire n23150;
   wire n23151;
   wire n23152;
   wire n23153;
   wire n23154;
   wire n23155;
   wire n23156;
   wire n23157;
   wire n23158;
   wire n23159;
   wire n23160;
   wire n23161;
   wire n23162;
   wire n23163;
   wire n23164;
   wire n23165;
   wire n23166;
   wire n23167;
   wire n23168;
   wire n23169;
   wire n23170;
   wire n23171;
   wire n23172;
   wire n23173;
   wire n23174;
   wire n23175;
   wire n23176;
   wire n23177;
   wire n23178;
   wire n23179;
   wire n23180;
   wire n23181;
   wire n23182;
   wire n23183;
   wire n23184;
   wire n23185;
   wire n23186;
   wire n23187;
   wire n23188;
   wire n23189;
   wire n23190;
   wire n23191;
   wire n23192;
   wire n23193;
   wire n23194;
   wire n23195;
   wire n23196;
   wire n23197;
   wire n23198;
   wire n23199;
   wire n23200;
   wire n23201;
   wire n23202;
   wire n23203;
   wire n23204;
   wire n23205;
   wire n23206;
   wire n23207;
   wire n23208;
   wire n23209;
   wire n23210;
   wire n23211;
   wire n23212;
   wire n23213;
   wire n23214;
   wire n23215;
   wire n23216;
   wire n23217;
   wire n23218;
   wire n23219;
   wire n23220;
   wire n23221;
   wire n23222;
   wire n23223;
   wire n23224;
   wire n23225;
   wire n23226;
   wire n23227;
   wire n23228;
   wire n23229;
   wire n23230;
   wire n23231;
   wire n23232;
   wire n23233;
   wire n23234;
   wire n23235;
   wire n23236;
   wire n23237;
   wire n23238;
   wire n23239;
   wire n23240;
   wire n23241;
   wire n23242;
   wire n23243;
   wire n23244;
   wire n23245;
   wire n23246;
   wire n23247;
   wire n23248;
   wire n23249;
   wire n23250;
   wire n23251;
   wire n23252;
   wire n23253;
   wire n23254;
   wire n23255;
   wire n23256;
   wire n23257;
   wire n23258;
   wire n23259;
   wire n23260;
   wire n23261;
   wire n23262;
   wire n23263;
   wire n23264;
   wire n23265;
   wire n23266;
   wire n23267;
   wire n23268;
   wire n23269;
   wire n23270;
   wire n23271;
   wire n23272;
   wire n23273;
   wire n23274;
   wire n23275;
   wire n23276;
   wire n23277;
   wire n23278;
   wire n23279;
   wire n23280;
   wire n23281;
   wire n23282;
   wire n23283;
   wire n23284;
   wire n23285;
   wire n23286;
   wire n23287;
   wire n23288;
   wire n23289;
   wire n23290;
   wire n23291;
   wire n23292;
   wire n23293;
   wire n23294;
   wire n23295;
   wire n23296;
   wire n23297;
   wire n23298;
   wire n23299;
   wire n23300;
   wire n23301;
   wire n23302;
   wire n23303;
   wire n23304;
   wire n23305;
   wire n23306;
   wire n23307;
   wire n23308;
   wire n23309;
   wire n23310;
   wire n23311;
   wire n23312;
   wire n23313;
   wire n23314;
   wire n23315;
   wire n23316;
   wire n23317;
   wire n23318;
   wire n23319;
   wire n23320;
   wire n23321;
   wire n23322;
   wire n23323;
   wire n23324;
   wire n23325;
   wire n23326;
   wire n23327;
   wire n23328;
   wire n23329;
   wire n23330;
   wire n23331;
   wire n23332;
   wire n23333;
   wire n23334;
   wire n23335;
   wire n23336;
   wire n23337;
   wire n23338;
   wire n23339;
   wire n23340;
   wire n23341;
   wire n23342;
   wire n23343;
   wire n23344;
   wire n23345;
   wire n23346;
   wire n23347;
   wire n23348;
   wire n23349;
   wire n23350;
   wire n23351;
   wire n23352;
   wire n23353;
   wire n23354;
   wire n23355;
   wire n23356;
   wire n23357;
   wire n23358;
   wire n23359;
   wire n23360;
   wire n23361;
   wire n23362;
   wire n23363;
   wire n23364;
   wire n23365;
   wire n23366;
   wire n23367;
   wire n23368;
   wire n23369;
   wire n23370;
   wire n23371;
   wire n23372;
   wire n23373;
   wire n23374;
   wire n23375;
   wire n23376;
   wire n23377;
   wire n23378;
   wire n23379;
   wire n23380;
   wire n23381;
   wire n23382;
   wire n23383;
   wire n23384;
   wire n23385;
   wire n23386;
   wire n23387;
   wire n23388;
   wire n23389;
   wire n23390;
   wire n23391;
   wire n23392;
   wire n23393;
   wire n23394;
   wire n23395;
   wire n23396;
   wire n23397;
   wire n23398;
   wire n23399;
   wire n23400;
   wire n23401;
   wire n23402;
   wire n23403;
   wire n23404;
   wire n23405;
   wire n23406;
   wire n23407;
   wire n23408;
   wire n23409;
   wire n23410;
   wire n23411;
   wire n23412;
   wire n23413;
   wire n23414;
   wire n23415;
   wire n23416;
   wire n23417;
   wire n23418;
   wire n23419;
   wire n23420;
   wire n23421;
   wire n23422;
   wire n23423;
   wire n23424;
   wire n23425;
   wire n23426;
   wire n23427;
   wire n23428;
   wire n23429;
   wire n23430;
   wire n23431;
   wire n23432;
   wire n23433;
   wire n23434;
   wire n23435;
   wire n23436;
   wire n23437;
   wire n23438;
   wire n23439;
   wire n23440;
   wire n23441;
   wire n23442;
   wire n23443;
   wire n23444;
   wire n23445;
   wire n23446;
   wire n23447;
   wire n23448;
   wire n23449;
   wire n23450;
   wire n23451;
   wire n23452;
   wire n23453;
   wire n23454;
   wire n23455;
   wire n23456;
   wire n23457;
   wire n23458;
   wire n23459;
   wire n23460;
   wire n23461;
   wire n23462;
   wire n23463;
   wire n23464;
   wire n23465;
   wire n23466;
   wire n23467;
   wire n23468;
   wire n23469;
   wire n23470;
   wire n23471;
   wire n23472;
   wire n23473;
   wire n23474;
   wire n23475;
   wire n23477;
   wire n23478;
   wire n23479;
   wire n23480;
   wire n23481;
   wire n23482;
   wire n23483;
   wire n23484;
   wire n23485;
   wire n23486;
   wire n23487;
   wire n23488;
   wire n23489;
   wire n23490;
   wire n23491;
   wire n23492;
   wire n23493;
   wire n23494;
   wire n23495;
   wire n23496;
   wire n23497;
   wire n23498;
   wire n23499;
   wire n23500;
   wire n23501;
   wire n23502;
   wire n23503;
   wire n23504;
   wire n23505;
   wire n23506;
   wire n23507;
   wire n23508;
   wire n23509;
   wire n23510;
   wire n23511;
   wire n23512;
   wire n23513;
   wire n23514;
   wire n23515;
   wire n23516;
   wire n23517;
   wire n23518;
   wire n23519;
   wire n23520;
   wire n23521;
   wire n23522;
   wire n23523;
   wire n23524;
   wire n23525;
   wire n23526;
   wire n23527;
   wire n23528;
   wire n23529;
   wire n23530;
   wire n23531;
   wire n23532;
   wire n23533;
   wire n23534;
   wire n23535;
   wire n23536;
   wire n23537;
   wire n23538;
   wire n23539;
   wire n23540;
   wire n23541;
   wire n23542;
   wire n23543;
   wire n23544;
   wire n23545;
   wire n23546;
   wire n23547;
   wire n23548;
   wire n23549;
   wire n23550;
   wire n23551;
   wire n23552;
   wire n23553;
   wire n23554;
   wire n23555;
   wire n23556;
   wire n23557;
   wire n23558;
   wire n23559;
   wire n23560;
   wire n23561;
   wire n23562;
   wire n23563;
   wire n23564;
   wire n23565;
   wire n23566;
   wire n23567;
   wire n23568;
   wire n23569;
   wire n23570;
   wire n23571;
   wire n23572;
   wire n23573;
   wire n23574;
   wire n23575;
   wire n23576;
   wire n23577;
   wire n23578;
   wire n23579;
   wire n23580;
   wire n23581;
   wire n23582;
   wire n23583;
   wire n23584;
   wire n23585;
   wire n23586;
   wire n23587;
   wire n23588;
   wire n23589;
   wire n23590;
   wire n23591;
   wire n23592;
   wire n23593;
   wire n23594;
   wire n23595;
   wire n23596;
   wire n23597;
   wire n23598;
   wire n23599;
   wire n23600;
   wire n23601;
   wire n23602;
   wire n23603;
   wire n23604;
   wire n23605;
   wire n23606;
   wire n23607;
   wire n23608;
   wire n23609;
   wire n23610;
   wire n23611;
   wire n23612;
   wire n23613;
   wire n23614;
   wire n23615;
   wire n23616;
   wire n23617;
   wire n23618;
   wire n23619;
   wire n23620;
   wire n23621;
   wire n23622;
   wire n23623;
   wire n23624;
   wire n23625;
   wire n23626;
   wire n23627;
   wire n23628;
   wire n23629;
   wire n23630;
   wire n23631;
   wire n23632;
   wire n23633;
   wire n23634;
   wire n23635;
   wire n23636;
   wire n23637;
   wire n23638;
   wire n23639;
   wire n23640;
   wire n23641;
   wire n23642;
   wire n23643;
   wire n23644;
   wire n23645;
   wire n23646;
   wire n23647;
   wire n23648;
   wire n23649;
   wire n23650;
   wire n23651;
   wire n23652;
   wire n23653;
   wire n23654;
   wire n23655;
   wire n23656;
   wire n23657;
   wire n23658;
   wire n23659;
   wire n23660;
   wire n23661;
   wire n23662;
   wire n23663;
   wire n23664;
   wire n23665;
   wire n23666;
   wire n23667;
   wire n23668;
   wire n23669;
   wire n23670;
   wire n23671;
   wire n23672;
   wire n23673;
   wire n23674;
   wire n23675;
   wire n23676;
   wire n23677;
   wire n23678;
   wire n23679;
   wire n23680;
   wire n23681;
   wire n23682;
   wire n23683;
   wire n23684;
   wire n23685;
   wire n23686;
   wire n23687;
   wire n23688;
   wire n23689;
   wire n23690;
   wire n23691;
   wire n23692;
   wire n23693;
   wire n23694;
   wire n23695;
   wire n23696;
   wire n23697;
   wire n23698;
   wire n23699;
   wire n23700;
   wire n23701;
   wire n23702;
   wire n23703;
   wire n23704;
   wire n23705;
   wire n23706;
   wire n23707;
   wire n23708;
   wire n23709;
   wire n23710;
   wire n23711;
   wire n23712;
   wire n23713;
   wire n23714;
   wire n23715;
   wire n23716;
   wire n23717;
   wire n23718;
   wire n23719;
   wire n23720;
   wire n23721;
   wire n23722;
   wire n23723;
   wire n23724;
   wire n23725;
   wire n23726;
   wire n23727;
   wire n23728;
   wire n23729;
   wire n23730;
   wire n23731;
   wire n23732;
   wire n23733;
   wire n23734;
   wire n23735;
   wire n23736;
   wire n23737;
   wire n23738;
   wire n23739;
   wire n23740;
   wire n23741;
   wire n23742;
   wire n23743;
   wire n23744;
   wire n23745;
   wire n23746;
   wire n23747;
   wire n23748;
   wire n23749;
   wire n23750;
   wire n23751;
   wire n23752;
   wire n23753;
   wire n23754;
   wire n23755;
   wire n23756;
   wire n23757;
   wire n23758;
   wire n23759;
   wire n23760;
   wire n23761;
   wire n23762;
   wire n23763;
   wire n23764;
   wire n23765;
   wire n23766;
   wire n23767;
   wire n23768;
   wire n23769;
   wire n23770;
   wire n23771;
   wire n23772;
   wire n23773;
   wire n23774;
   wire n23775;
   wire n23776;
   wire n23777;
   wire n23778;
   wire n23779;
   wire n23780;
   wire n23781;
   wire n23782;
   wire n23783;
   wire n23784;
   wire n23785;
   wire n23786;
   wire n23787;
   wire n23788;
   wire n23789;
   wire n23790;
   wire n23791;
   wire n23792;
   wire n23793;
   wire n23794;
   wire n23795;
   wire n23796;
   wire n23797;
   wire n23798;
   wire n23799;
   wire n23800;
   wire n23801;
   wire n23802;
   wire n23803;
   wire n23804;
   wire n23805;
   wire n23806;
   wire n23807;
   wire n23808;
   wire n23809;
   wire n23810;
   wire n23811;
   wire n23812;
   wire n23813;
   wire n23814;
   wire n23815;
   wire n23816;
   wire n23817;
   wire n23818;
   wire n23819;
   wire n23820;
   wire n23821;
   wire n23822;
   wire n23823;
   wire n23824;
   wire n23825;
   wire n23826;
   wire n23827;
   wire n23828;
   wire n23829;
   wire n23830;
   wire n23831;
   wire n23832;
   wire n23833;
   wire n23834;
   wire n23835;
   wire n23836;
   wire n23837;
   wire n23838;
   wire n23839;
   wire n23840;
   wire n23841;
   wire n23842;
   wire n23843;
   wire n23844;
   wire n23845;
   wire n23846;
   wire n23847;
   wire n23848;
   wire n23849;
   wire n23850;
   wire n23851;
   wire n23852;
   wire n23853;
   wire n23854;
   wire n23855;
   wire n23856;
   wire n23857;
   wire n23858;
   wire n23859;
   wire n23860;
   wire n23861;
   wire n23862;
   wire n23863;
   wire n23864;
   wire n23865;
   wire n23866;
   wire n23867;
   wire n23868;
   wire n23869;
   wire n23870;
   wire n23871;
   wire n23872;
   wire n23873;
   wire n23874;
   wire n23875;
   wire n23876;
   wire n23877;
   wire n23878;
   wire n23879;
   wire n23880;
   wire n23881;
   wire n23882;
   wire n23883;
   wire n23884;
   wire n23885;
   wire n23886;
   wire n23887;
   wire n23888;
   wire n23889;
   wire n23890;
   wire n23891;
   wire n23892;
   wire n23893;
   wire n23894;
   wire n23895;
   wire n23896;
   wire n23897;
   wire n23898;
   wire n23899;
   wire n23900;
   wire n23901;
   wire n23902;
   wire n23903;
   wire n23904;
   wire n23905;
   wire n23906;
   wire n23907;
   wire n23908;
   wire n23909;
   wire n23910;
   wire n23911;
   wire n23912;
   wire n23913;
   wire n23914;
   wire n23915;
   wire n23916;
   wire n23917;
   wire n23918;
   wire n23919;
   wire n23920;
   wire n23921;
   wire n23922;
   wire n23923;
   wire n23924;
   wire n23925;
   wire n23926;
   wire n23927;
   wire n23928;
   wire n23929;
   wire n23930;
   wire n23931;
   wire n23932;
   wire n23933;
   wire n23934;
   wire n23935;
   wire n23936;
   wire n23937;
   wire n23938;
   wire n23939;
   wire n23940;
   wire n23941;
   wire n23942;
   wire n23943;
   wire n23944;
   wire n23945;
   wire n23946;
   wire n23947;
   wire n23948;
   wire n23949;
   wire n23950;
   wire n23951;
   wire n23952;
   wire n23953;
   wire n23954;
   wire n23955;
   wire n23956;
   wire n23957;
   wire n23958;
   wire n23959;
   wire n23960;
   wire n23961;
   wire n23962;
   wire n23963;
   wire n23964;
   wire n23965;
   wire n23966;
   wire n23967;
   wire n23968;
   wire n23969;
   wire n23970;
   wire n23971;
   wire n23972;
   wire n23973;
   wire n23974;
   wire n23975;
   wire n23976;
   wire n23977;
   wire n23978;
   wire n23979;
   wire n23980;
   wire n23981;
   wire n23982;
   wire n23983;
   wire n23984;
   wire n23985;
   wire n23986;
   wire n23987;
   wire n23988;
   wire n23989;
   wire n23990;
   wire n23991;
   wire n23992;
   wire n23993;
   wire n23994;
   wire n23995;
   wire n23996;
   wire n23997;
   wire n23998;
   wire n23999;
   wire n24000;
   wire n24001;
   wire n24002;
   wire n24003;
   wire n24004;
   wire n24005;
   wire n24006;
   wire n24007;
   wire n24008;
   wire n24009;
   wire n24010;
   wire n24011;
   wire n24012;
   wire n24013;
   wire n24014;
   wire n24015;
   wire n24016;
   wire n24017;
   wire n24018;
   wire n24019;
   wire n24020;
   wire n24021;
   wire n24022;
   wire n24023;
   wire n24024;
   wire n24025;
   wire n24026;
   wire n24027;
   wire n24028;
   wire n24029;
   wire n24030;
   wire n24031;
   wire n24032;
   wire n24033;
   wire n24034;
   wire n24035;
   wire n24036;
   wire n24038;
   wire n24039;
   wire n24040;
   wire n24041;
   wire n24042;
   wire n24043;
   wire n24044;
   wire n24045;
   wire n24046;
   wire n24047;
   wire n24048;
   wire n24049;
   wire n24050;
   wire n24051;
   wire n24052;
   wire n24053;
   wire n24054;
   wire n24055;
   wire n24056;
   wire n24057;
   wire n24058;
   wire n24059;
   wire n24060;
   wire n24061;
   wire n24062;
   wire n24063;
   wire n24064;
   wire n24065;
   wire n24066;
   wire n24067;
   wire n24068;
   wire n24069;
   wire n24070;
   wire n24071;
   wire n24072;
   wire n24073;
   wire n24074;
   wire n24075;
   wire n24076;
   wire n24077;
   wire n24078;
   wire n24079;
   wire n24080;
   wire n24081;
   wire n24082;
   wire n24083;
   wire n24084;
   wire n24085;
   wire n24086;
   wire n24087;
   wire n24089;
   wire n24090;
   wire n24091;
   wire n24092;
   wire n24093;
   wire n24094;
   wire n24095;
   wire n24096;
   wire n24097;
   wire n24098;
   wire n24099;
   wire n24100;
   wire n24101;
   wire n24102;
   wire n24103;
   wire n24104;
   wire n24105;
   wire n24106;
   wire n24107;
   wire n24108;
   wire n24109;
   wire n24110;
   wire n24111;
   wire n24112;
   wire n24113;
   wire n24114;
   wire n24115;
   wire n24116;
   wire n24117;
   wire n24118;
   wire n24119;
   wire n24120;
   wire n24121;
   wire n24122;
   wire n24123;
   wire n24124;
   wire n24125;
   wire n24126;
   wire n24127;
   wire n24128;
   wire n24130;
   wire n24131;
   wire n24132;
   wire n24133;
   wire n24134;
   wire n24135;
   wire n24136;
   wire n24137;
   wire n24138;
   wire n24139;
   wire n24140;
   wire n24141;
   wire n24142;
   wire n24143;
   wire n24144;
   wire n24145;
   wire n24146;
   wire n24147;
   wire n24148;
   wire n24149;
   wire n24150;
   wire n24151;
   wire n24152;
   wire n24153;
   wire n24154;
   wire n24155;
   wire n24156;
   wire n24157;
   wire n24158;
   wire n24159;
   wire n24160;
   wire n24161;
   wire n24162;
   wire n24163;
   wire n24164;
   wire n24165;
   wire n24166;
   wire n24167;
   wire n24168;
   wire n24169;
   wire n24170;
   wire n24171;
   wire n24172;
   wire n24173;
   wire n24174;
   wire n24175;
   wire n24176;
   wire n24177;
   wire n24178;
   wire n24179;
   wire n24180;
   wire n24181;
   wire n24182;
   wire n24183;
   wire n24184;
   wire n24185;
   wire n24186;
   wire n24187;
   wire n24188;
   wire n24189;
   wire n24190;
   wire n24191;
   wire n24192;
   wire n24193;
   wire n24194;
   wire n24195;
   wire n24196;
   wire n24197;
   wire n24198;
   wire n24199;
   wire n24200;
   wire n24201;
   wire n24202;
   wire n24203;
   wire n24204;
   wire n24205;
   wire n24206;
   wire n24207;
   wire n24208;
   wire n24209;
   wire n24210;
   wire n24211;
   wire n24212;
   wire n24213;
   wire n24214;
   wire n24215;
   wire n24216;
   wire n24217;
   wire n24218;
   wire n24219;
   wire n24220;
   wire n24222;
   wire n24223;
   wire n24224;
   wire n24225;
   wire n24226;
   wire n24227;
   wire n24228;
   wire n24229;
   wire n24230;
   wire n24231;
   wire n24232;
   wire n24233;
   wire n24234;
   wire n24235;
   wire n24236;
   wire n24237;
   wire n24238;
   wire n24239;
   wire n24240;
   wire n24241;
   wire n24242;
   wire n24243;
   wire n24244;
   wire n24245;
   wire n24246;
   wire n24247;
   wire n24248;
   wire n24249;
   wire n24250;
   wire n24251;
   wire n24252;
   wire n24253;
   wire n24254;
   wire n24255;
   wire n24256;
   wire n24257;
   wire n24258;
   wire n24259;
   wire n24260;
   wire n24261;
   wire n24262;
   wire n24263;
   wire n24264;
   wire n24265;
   wire n24266;
   wire n24267;
   wire n24268;
   wire n24269;
   wire n24270;
   wire n24271;
   wire n24272;
   wire n24273;
   wire n24274;
   wire n24275;
   wire n24276;
   wire n24277;
   wire n24278;
   wire n24279;
   wire n24280;
   wire n24281;
   wire n24282;
   wire n24283;
   wire n24284;
   wire n24285;
   wire n24286;
   wire n24287;
   wire n24288;
   wire n24289;
   wire n24290;
   wire n24291;
   wire n24292;
   wire n24293;
   wire n24294;
   wire n24295;
   wire n24296;
   wire n24297;
   wire n24298;
   wire n24299;
   wire n24300;
   wire n24301;
   wire n24302;
   wire n24303;
   wire n24304;
   wire n24305;
   wire n24306;
   wire n24307;
   wire n24308;
   wire n24309;
   wire n24310;
   wire n24311;
   wire n24312;
   wire n24313;
   wire n24314;
   wire n24315;
   wire n24316;
   wire n24317;
   wire n24318;
   wire n24319;
   wire n24320;
   wire n24321;
   wire n24322;
   wire n24323;
   wire n24324;
   wire n24325;
   wire n24326;
   wire n24327;
   wire n24328;
   wire n24329;
   wire n24330;
   wire n24331;
   wire n24332;
   wire n24333;
   wire n24334;
   wire n24335;
   wire n24336;
   wire n24337;
   wire n24338;
   wire n24339;
   wire n24340;
   wire n24341;
   wire n24342;
   wire n24343;
   wire n24345;
   wire n24346;
   wire n24347;
   wire n24348;
   wire n24351;
   wire n24352;
   wire n24353;
   wire n24354;
   wire n24355;
   wire n24356;
   wire n24357;
   wire n24358;
   wire n24359;
   wire n24360;
   wire n24361;
   wire n24362;
   wire n24363;
   wire n24364;
   wire n24365;
   wire n24366;
   wire n24367;
   wire n24368;
   wire n24369;
   wire n24370;
   wire n24371;
   wire n24372;
   wire n24373;
   wire n24374;
   wire n24375;
   wire n24376;
   wire n24377;
   wire n24378;
   wire n24379;
   wire n24380;
   wire n24381;
   wire n24382;
   wire n24383;
   wire n24384;
   wire n24385;
   wire n24386;
   wire n24387;
   wire n24388;
   wire n24389;
   wire n24390;
   wire n24391;
   wire n24392;
   wire n24393;
   wire n24394;
   wire n24395;
   wire n24396;
   wire n24398;
   wire n24399;
   wire n24400;
   wire n24401;
   wire n24402;
   wire n24403;
   wire n24404;
   wire n24405;
   wire n24406;
   wire n24407;
   wire n24408;
   wire n24409;
   wire n24410;
   wire n24411;
   wire n24412;
   wire n24413;
   wire n24414;
   wire n24415;
   wire n24416;
   wire n24417;
   wire n24418;
   wire n24419;
   wire n24420;
   wire n24421;
   wire n24422;
   wire n24423;
   wire n24424;
   wire n24425;
   wire n24426;
   wire n24427;
   wire n24428;
   wire n24429;
   wire n24430;
   wire n24431;
   wire n24432;
   wire n24433;
   wire n24434;
   wire n24435;
   wire n24436;
   wire n24437;
   wire n24438;
   wire n24439;
   wire n24440;
   wire n24441;
   wire n24442;
   wire n24443;
   wire n24444;
   wire n24445;
   wire n24446;
   wire n24447;
   wire n24449;
   wire n24450;
   wire n24451;
   wire n24452;
   wire n24453;
   wire n24454;
   wire n24455;
   wire n24456;
   wire n24457;
   wire n24458;
   wire n24459;
   wire n24460;
   wire n24461;
   wire n24463;
   wire n24464;
   wire n24465;
   wire n24466;
   wire n24467;
   wire n24468;
   wire n24470;
   wire n24471;
   wire n24472;
   wire n24473;
   wire n24474;
   wire n24475;
   wire n24476;
   wire n24477;
   wire n24478;
   wire n24479;
   wire n24480;
   wire n24481;
   wire n24482;
   wire n24483;
   wire n24484;
   wire n24485;
   wire n24486;
   wire n24487;
   wire n24488;
   wire n24489;
   wire n24490;
   wire n24491;
   wire n24492;
   wire n24493;
   wire n24494;
   wire n24495;
   wire n24496;
   wire n24497;
   wire n24498;
   wire n24499;
   wire n24500;
   wire n24501;
   wire n24502;
   wire n24503;
   wire n24504;
   wire n24505;
   wire n24506;
   wire n24507;
   wire n24508;
   wire n24509;
   wire n24510;
   wire n24511;
   wire n24512;
   wire n24513;
   wire n24514;
   wire n24515;
   wire n24516;
   wire n24517;
   wire n24518;
   wire n24519;
   wire n24520;
   wire n24521;
   wire n24522;
   wire n24523;
   wire n24524;
   wire n24525;
   wire n24526;
   wire n24527;
   wire n24528;
   wire n24529;
   wire n24530;
   wire n24531;
   wire n24532;
   wire n24533;
   wire n24534;
   wire n24535;
   wire n24536;
   wire n24537;
   wire n24538;
   wire n24539;
   wire n24540;
   wire n24541;
   wire n24542;
   wire n24543;
   wire n24544;
   wire n24545;
   wire n24546;
   wire n24547;
   wire n24548;
   wire n24549;
   wire n24550;
   wire n24551;
   wire n24552;
   wire n24553;
   wire n24554;
   wire n24555;
   wire n24556;
   wire n24557;
   wire n24558;
   wire n24559;
   wire n24560;
   wire n24561;
   wire n24562;
   wire n24563;
   wire n24564;
   wire n24565;
   wire n24566;
   wire n24567;
   wire n24568;
   wire n24569;
   wire n24570;
   wire n24571;
   wire n24572;
   wire n24573;
   wire n24574;
   wire n24575;
   wire n24576;
   wire n24577;
   wire n24578;
   wire n24579;
   wire n24580;
   wire n24581;
   wire n24582;
   wire n24583;
   wire n24584;
   wire n24585;
   wire n24586;
   wire n24587;
   wire n24588;
   wire n24589;
   wire n24590;
   wire n24591;
   wire n24592;
   wire n24593;
   wire n24594;
   wire n24595;
   wire n24596;
   wire n24597;
   wire n24598;
   wire n24599;
   wire n24600;
   wire n24601;
   wire n24602;
   wire n24603;
   wire n24604;
   wire n24605;
   wire n24606;
   wire n24607;
   wire n24608;
   wire n24609;
   wire n24610;
   wire n24611;
   wire n24612;
   wire n24613;
   wire n24614;
   wire n24615;
   wire n24616;
   wire n24617;
   wire n24618;
   wire n24619;
   wire n24620;
   wire n24621;
   wire n24622;
   wire n24623;
   wire n24624;
   wire n24625;
   wire n24626;
   wire n24627;
   wire n24628;
   wire n24629;
   wire n24630;
   wire n24631;
   wire n24632;
   wire n24633;
   wire n24634;
   wire n24635;
   wire n24636;
   wire n24637;
   wire n24638;
   wire n24639;
   wire n24640;
   wire n24641;
   wire n24642;
   wire n24643;
   wire n24644;
   wire n24645;
   wire n24646;
   wire n24647;
   wire n24648;
   wire n24649;
   wire n24650;
   wire n24651;
   wire n24652;
   wire n24653;
   wire n24654;
   wire n24655;
   wire n24656;
   wire n24657;
   wire n24658;
   wire n24659;
   wire n24660;
   wire n24661;
   wire n24662;
   wire n24663;
   wire n24664;
   wire n24665;
   wire n24666;
   wire n24667;
   wire n24668;
   wire n24669;
   wire n24670;
   wire n24671;
   wire n24672;
   wire n24673;
   wire n24674;
   wire n24675;
   wire n24676;
   wire n24677;
   wire n24678;
   wire n24679;
   wire n24680;
   wire n24681;
   wire n24682;
   wire n24683;
   wire n24684;
   wire n24685;
   wire n24686;
   wire n24687;
   wire n24688;
   wire n24689;
   wire n24690;
   wire n24691;
   wire n24692;
   wire n24693;
   wire n24694;
   wire n24695;
   wire n24696;
   wire n24697;
   wire n24698;
   wire n24699;
   wire n24700;
   wire n24701;
   wire n24702;
   wire n24703;
   wire n24704;
   wire n24705;
   wire n24706;
   wire n24707;
   wire n24708;
   wire n24709;
   wire n24710;
   wire n24711;
   wire n24712;
   wire n24713;
   wire n24714;
   wire n24715;
   wire n24716;
   wire n24717;
   wire n24718;
   wire n24719;
   wire n24720;
   wire n24721;
   wire n24722;
   wire n24723;
   wire n24724;
   wire n24725;
   wire n24726;
   wire n24727;
   wire n24728;
   wire n24729;
   wire n24730;
   wire n24731;
   wire n24732;
   wire n24733;
   wire n24734;
   wire n24735;
   wire n24736;
   wire n24737;
   wire n24738;
   wire n24739;
   wire n24740;
   wire n24741;
   wire n24742;
   wire n24743;
   wire n24744;
   wire n24745;
   wire n24746;
   wire n24747;
   wire n24748;
   wire n24749;
   wire n24750;
   wire n24751;
   wire n24752;
   wire n24754;
   wire n24755;
   wire n24756;
   wire n24757;
   wire n24758;
   wire n24759;
   wire n24760;
   wire n24761;
   wire n24762;
   wire n24763;
   wire n24764;
   wire n24765;
   wire n24766;
   wire n24767;
   wire n24768;
   wire n24769;
   wire n24770;
   wire n24771;
   wire n24772;
   wire n24773;
   wire n24774;
   wire n24775;
   wire n24776;
   wire n24777;
   wire n24778;
   wire n24779;
   wire n24780;
   wire n24781;
   wire n24782;
   wire n24783;
   wire n24784;
   wire n24785;
   wire n24786;
   wire n24787;
   wire n24788;
   wire n24789;
   wire n24790;
   wire n24791;
   wire n24792;
   wire n24793;
   wire n24794;
   wire n24795;
   wire n24796;
   wire n24797;
   wire n24798;
   wire n24799;
   wire n24800;
   wire n24801;
   wire n24802;
   wire n24803;
   wire n24804;
   wire n24805;
   wire n24806;
   wire n24807;
   wire n24808;
   wire n24809;
   wire n24810;
   wire n24811;
   wire n24812;
   wire n24813;
   wire n24814;
   wire n24815;
   wire n24816;
   wire n24817;
   wire n24818;
   wire n24819;
   wire n24820;
   wire n24821;
   wire n24822;
   wire n24823;
   wire n24824;
   wire n24825;
   wire n24826;
   wire n24827;
   wire n24828;
   wire n24829;
   wire n24830;
   wire n24831;
   wire n24832;
   wire n24833;
   wire n24834;
   wire n24835;
   wire n24836;
   wire n24837;
   wire n24838;
   wire n24839;
   wire n24840;
   wire n24841;
   wire n24842;
   wire n24843;
   wire n24844;
   wire n24845;
   wire n24846;
   wire n24847;
   wire n24848;
   wire n24849;
   wire n24850;
   wire n24851;
   wire n24852;
   wire n24853;
   wire n24854;
   wire n24855;
   wire n24856;
   wire n24857;
   wire n24858;
   wire n24859;
   wire n24860;
   wire n24861;
   wire n24862;
   wire n24863;
   wire n24864;
   wire n24865;
   wire n24866;
   wire n24867;
   wire n24868;
   wire n24869;
   wire n24870;
   wire n24871;
   wire n24872;
   wire n24873;
   wire n24874;
   wire n24875;
   wire n24876;
   wire n24877;
   wire n24878;
   wire n24879;
   wire n24880;
   wire n24881;
   wire n24882;
   wire n24883;
   wire n24884;
   wire n24885;
   wire n24886;
   wire n24887;
   wire n24888;
   wire n24889;
   wire n24890;
   wire n24891;
   wire n24892;
   wire n24893;
   wire n24894;
   wire n24895;
   wire n24896;
   wire n24897;
   wire n24898;
   wire n24899;
   wire n24900;
   wire n24901;
   wire n24902;
   wire n24903;
   wire n24904;
   wire n24905;
   wire n24906;
   wire n24907;
   wire n24908;
   wire n24909;
   wire n24910;
   wire n24911;
   wire n24912;
   wire n24913;
   wire n24914;
   wire n24915;
   wire n24916;
   wire n24917;
   wire n24918;
   wire n24919;
   wire n24920;
   wire n24921;
   wire n24922;
   wire n24923;
   wire n24924;
   wire n24925;
   wire n24926;
   wire n24927;
   wire n24928;
   wire n24929;
   wire n24930;
   wire n24931;
   wire n24932;
   wire n24933;
   wire n24934;
   wire n24935;
   wire n24936;
   wire n24937;
   wire n24938;
   wire n24939;
   wire n24940;
   wire n24941;
   wire n24942;
   wire n24943;
   wire n24944;
   wire n24945;
   wire n24946;
   wire n24947;
   wire n24948;
   wire n24949;
   wire n24950;
   wire n24951;
   wire n24952;
   wire n24953;
   wire n24954;
   wire n24955;
   wire n24956;
   wire n24957;
   wire n24958;
   wire n24959;
   wire n24960;
   wire n24961;
   wire n24962;
   wire n24963;
   wire n24964;
   wire n24965;
   wire n24966;
   wire n24967;
   wire n24968;
   wire n24970;
   wire n24971;
   wire n24972;
   wire n24973;
   wire n24974;
   wire n24975;
   wire n24976;
   wire n24977;
   wire n24978;
   wire n24979;
   wire n24980;
   wire n24981;
   wire n24982;
   wire n24983;
   wire n24984;
   wire n24985;
   wire n24986;
   wire n24987;
   wire n24988;
   wire n24989;
   wire n24990;
   wire n24991;
   wire n24992;
   wire n24993;
   wire n24994;
   wire n24995;
   wire n24996;
   wire n24997;
   wire n24998;
   wire n24999;
   wire n25000;
   wire n25001;
   wire n25002;
   wire n25003;
   wire n25004;
   wire n25005;
   wire n25006;
   wire n25007;
   wire n25008;
   wire n25009;
   wire n25010;
   wire n25011;
   wire n25012;
   wire n25013;
   wire n25014;
   wire n25015;
   wire n25016;
   wire n25017;
   wire n25018;
   wire n25019;
   wire n25020;
   wire n25021;
   wire n25022;
   wire n25023;
   wire n25024;
   wire n25025;
   wire n25026;
   wire n25027;
   wire n25028;
   wire n25029;
   wire n25030;
   wire n25031;
   wire n25032;
   wire n25033;
   wire n25034;
   wire n25035;
   wire n25036;
   wire n25037;
   wire n25038;
   wire n25039;
   wire n25040;
   wire n25041;
   wire n25042;
   wire n25043;
   wire n25044;
   wire n25045;
   wire n25046;
   wire n25047;
   wire n25048;
   wire n25049;
   wire n25050;
   wire n25051;
   wire n25052;
   wire n25053;
   wire n25054;
   wire n25055;
   wire n25056;
   wire n25057;
   wire n25058;
   wire n25059;
   wire n25060;
   wire n25061;
   wire n25062;
   wire n25063;
   wire n25064;
   wire n25065;
   wire n25066;
   wire n25067;
   wire n25068;
   wire n25069;
   wire n25070;
   wire n25071;
   wire n25072;
   wire n25073;
   wire n25074;
   wire n25076;
   wire n25077;
   wire n25078;
   wire n25079;
   wire n25080;
   wire n25081;
   wire n25082;
   wire n25083;
   wire n25084;
   wire n25085;
   wire n25086;
   wire n25087;
   wire n25088;
   wire n25089;
   wire n25090;
   wire n25091;
   wire n25092;
   wire n25093;
   wire n25094;
   wire n25095;
   wire n25096;
   wire n25097;
   wire n25098;
   wire n25099;
   wire n25100;
   wire n25101;
   wire n25102;
   wire n25103;
   wire n25104;
   wire n25105;
   wire n25106;
   wire n25107;
   wire n25108;
   wire n25109;
   wire n25110;
   wire n25111;
   wire n25112;
   wire n25113;
   wire n25114;
   wire n25115;
   wire n25116;
   wire n25117;
   wire n25118;
   wire n25119;
   wire n25121;
   wire n25122;
   wire n25123;
   wire n25124;
   wire n25125;
   wire n25126;
   wire n25127;
   wire n25128;
   wire n25129;
   wire n25130;
   wire n25131;
   wire n25132;
   wire n25133;
   wire n25134;
   wire n25135;
   wire n25136;
   wire n25137;
   wire n25138;
   wire n25139;
   wire n25140;
   wire n25141;
   wire n25142;
   wire n25143;
   wire n25144;
   wire n25145;
   wire n25146;
   wire n25147;
   wire n25148;
   wire n25149;
   wire n25150;
   wire n25151;
   wire n25152;
   wire n25153;
   wire n25154;
   wire n25155;
   wire n25156;
   wire n25157;
   wire n25158;
   wire n25159;
   wire n25160;
   wire n25161;
   wire n25162;
   wire n25163;
   wire n25164;
   wire n25165;
   wire n25166;
   wire n25167;
   wire n25168;
   wire n25169;
   wire n25170;
   wire n25171;
   wire n25172;
   wire n25173;
   wire n25174;
   wire n25175;
   wire n25176;
   wire n25177;
   wire n25178;
   wire n25179;
   wire n25180;
   wire n25181;
   wire n25182;
   wire n25183;
   wire n25184;
   wire n25185;
   wire n25186;
   wire n25187;
   wire n25188;
   wire n25189;
   wire n25190;
   wire n25191;
   wire n25192;
   wire n25193;
   wire n25194;
   wire n25195;
   wire n25196;
   wire n25197;
   wire n25198;
   wire n25199;
   wire n25200;
   wire n25201;
   wire n25202;
   wire n25203;
   wire n25204;
   wire n25205;
   wire n25206;
   wire n25207;
   wire n25208;
   wire n25209;
   wire n25210;
   wire n25211;
   wire n25212;
   wire n25213;
   wire n25214;
   wire n25215;
   wire n25216;
   wire n25217;
   wire n25218;
   wire n25219;
   wire n25220;
   wire n25221;
   wire n25222;
   wire n25223;
   wire n25224;
   wire n25225;
   wire n25226;
   wire n25227;
   wire n25228;
   wire n25229;
   wire n25230;
   wire n25231;
   wire n25232;
   wire n25233;
   wire n25234;
   wire n25235;
   wire n25236;
   wire n25237;
   wire n25238;
   wire n25239;
   wire n25240;
   wire n25241;
   wire n25242;
   wire n25243;
   wire n25244;
   wire n25245;
   wire n25246;
   wire n25247;
   wire n25248;
   wire n25249;
   wire n25250;
   wire n25251;
   wire n25252;
   wire n25253;
   wire n25254;
   wire n25255;
   wire n25256;
   wire n25257;
   wire n25258;
   wire n25259;
   wire n25260;
   wire n25261;
   wire n25262;
   wire n25263;
   wire n25264;
   wire n25265;
   wire n25266;
   wire n25267;
   wire n25268;
   wire n25269;
   wire n25270;
   wire n25271;
   wire n25272;
   wire n25273;
   wire n25274;
   wire n25275;
   wire n25276;
   wire n25277;
   wire n25278;
   wire n25279;
   wire n25280;
   wire n25281;
   wire n25282;
   wire n25283;
   wire n25284;
   wire n25285;
   wire n25286;
   wire n25287;
   wire n25288;
   wire n25289;
   wire n25290;
   wire n25291;
   wire n25292;
   wire n25293;
   wire n25294;
   wire n25295;
   wire n25296;
   wire n25297;
   wire n25298;
   wire n25299;
   wire n25300;
   wire n25301;
   wire n25302;
   wire n25303;
   wire n25304;
   wire n25305;
   wire n25306;
   wire n25307;
   wire n25308;
   wire n25309;
   wire n25310;
   wire n25311;
   wire n25312;
   wire n25313;
   wire n25314;
   wire n25315;
   wire n25316;
   wire n25317;
   wire n25318;
   wire n25319;
   wire n25320;
   wire n25321;
   wire n25322;
   wire n25323;
   wire n25324;
   wire n25325;
   wire n25326;
   wire n25327;
   wire n25328;
   wire n25329;
   wire n25330;
   wire n25331;
   wire n25332;
   wire n25333;
   wire n25334;
   wire n25335;
   wire n25336;
   wire n25337;
   wire n25338;
   wire n25339;
   wire n25340;
   wire n25341;
   wire n25342;
   wire n25343;
   wire n25344;
   wire n25345;
   wire n25346;
   wire n25347;
   wire n25348;
   wire n25349;
   wire n25350;
   wire n25351;
   wire n25352;
   wire n25353;
   wire n25354;
   wire n25355;
   wire n25356;
   wire n25357;
   wire n25358;
   wire n25359;
   wire n25360;
   wire n25361;
   wire n25362;
   wire n25363;
   wire n25364;
   wire n25365;
   wire n25366;
   wire n25367;
   wire n25368;
   wire n25369;
   wire n25370;
   wire n25371;
   wire n25372;
   wire n25373;
   wire n25374;
   wire n25375;
   wire n25376;
   wire n25377;
   wire n25378;
   wire n25379;
   wire n25380;
   wire n25381;
   wire n25382;
   wire n25383;
   wire n25384;
   wire n25386;
   wire n25387;
   wire n25388;
   wire n25389;
   wire n25390;
   wire n25391;
   wire n25392;
   wire n25393;
   wire n25394;
   wire n25395;
   wire n25396;
   wire n25397;
   wire n25398;
   wire n25399;
   wire n25400;
   wire n25401;
   wire n25402;
   wire n25403;
   wire n25404;
   wire n25405;
   wire n25406;
   wire n25407;
   wire n25408;
   wire n25409;
   wire n25410;
   wire n25411;
   wire n25412;
   wire n25413;
   wire n25414;
   wire n25415;
   wire n25416;
   wire n25417;
   wire n25418;
   wire n25419;
   wire n25420;
   wire n25421;
   wire n25422;
   wire n25423;
   wire n25425;
   wire n25426;
   wire n25427;
   wire n25428;
   wire n25429;
   wire n25430;
   wire n25431;
   wire n25432;
   wire n25433;
   wire n25434;
   wire n25435;
   wire n25436;
   wire n25437;
   wire n25438;
   wire n25439;
   wire n25440;
   wire n25441;
   wire n25442;
   wire n25443;
   wire n25444;
   wire n25445;
   wire n25446;
   wire n25447;
   wire n25448;
   wire n25449;
   wire n25450;
   wire n25451;
   wire n25452;
   wire n25453;
   wire n25454;
   wire n25455;
   wire n25456;
   wire n25457;
   wire n25458;
   wire n25459;
   wire n25460;
   wire n25461;
   wire n25462;
   wire n25463;
   wire n25464;
   wire n25465;
   wire n25466;
   wire n25467;
   wire n25468;
   wire n25469;
   wire n25470;
   wire n25471;
   wire n25472;
   wire n25473;
   wire n25474;
   wire n25475;
   wire n25476;
   wire n25477;
   wire n25478;
   wire n25479;
   wire n25480;
   wire n25481;
   wire n25482;
   wire n25483;
   wire n25484;
   wire n25485;
   wire n25486;
   wire n25487;
   wire n25488;
   wire n25489;
   wire n25490;
   wire n25491;
   wire n25492;
   wire n25493;
   wire n25494;
   wire n25495;
   wire n25496;
   wire n25497;
   wire n25498;
   wire n25499;
   wire n25500;
   wire n25501;
   wire n25502;
   wire n25503;
   wire n25504;
   wire n25505;
   wire n25506;
   wire n25507;
   wire n25508;
   wire n25509;
   wire n25510;
   wire n25511;
   wire n25512;
   wire n25513;
   wire n25514;
   wire n25515;
   wire n25516;
   wire n25517;
   wire n25518;
   wire n25519;
   wire n25520;
   wire n25521;
   wire n25522;
   wire n25523;
   wire n25524;
   wire n25525;
   wire n25526;
   wire n25527;
   wire n25528;
   wire n25529;
   wire n25530;
   wire n25531;
   wire n25532;
   wire n25533;
   wire n25534;
   wire n25535;
   wire n25536;
   wire n25537;
   wire n25538;
   wire n25539;
   wire n25540;
   wire n25541;
   wire n25542;
   wire n25543;
   wire n25544;
   wire n25545;
   wire n25546;
   wire n25547;
   wire n25548;
   wire n25549;
   wire n25550;
   wire n25551;
   wire n25552;
   wire n25553;
   wire n25554;
   wire n25555;
   wire n25556;
   wire n25557;
   wire n25558;
   wire n25559;
   wire n25560;
   wire n25561;
   wire n25562;
   wire n25563;
   wire n25564;
   wire n25565;
   wire n25566;
   wire n25567;
   wire n25568;
   wire n25569;
   wire n25570;
   wire n25571;
   wire n25572;
   wire n25573;
   wire n25574;
   wire n25575;
   wire n25576;
   wire n25577;
   wire n25578;
   wire n25579;
   wire n25580;
   wire n25581;
   wire n25582;
   wire n25583;
   wire n25584;
   wire n25585;
   wire n25586;
   wire n25587;
   wire n25588;
   wire n25589;
   wire n25590;
   wire n25591;
   wire n25592;
   wire n25593;
   wire n25594;
   wire n25595;
   wire n25596;
   wire n25597;
   wire n25598;
   wire n25599;
   wire n25600;
   wire n25601;
   wire n25602;
   wire n25603;
   wire n25604;
   wire n25605;
   wire n25606;
   wire n25607;
   wire n25608;
   wire n25609;
   wire n25610;
   wire n25611;
   wire n25612;
   wire n25613;
   wire n25614;
   wire n25615;
   wire n25616;
   wire n25617;
   wire n25618;
   wire n25619;
   wire n25620;
   wire n25621;
   wire n25622;
   wire n25623;
   wire n25624;
   wire n25625;
   wire n25626;
   wire n25627;
   wire n25628;
   wire n25629;
   wire n25630;
   wire n25631;
   wire n25632;
   wire n25633;
   wire n25634;
   wire n25635;
   wire n25636;
   wire n25637;
   wire n25638;
   wire n25639;
   wire n25640;
   wire n25641;
   wire n25642;
   wire n25643;
   wire n25644;
   wire n25645;
   wire n25646;
   wire n25647;
   wire n25648;
   wire n25649;
   wire n25650;
   wire n25651;
   wire n25652;
   wire n25653;
   wire n25654;
   wire n25655;
   wire n25656;
   wire n25657;
   wire n25658;
   wire n25659;
   wire n25660;
   wire n25661;
   wire n25662;
   wire n25663;
   wire n25664;
   wire n25665;
   wire n25666;
   wire n25667;
   wire n25668;
   wire n25669;
   wire n25670;
   wire n25671;
   wire n25672;
   wire n25673;
   wire n25674;
   wire n25675;
   wire n25676;
   wire n25677;
   wire n25678;
   wire n25679;
   wire n25680;
   wire n25681;
   wire n25682;
   wire n25683;
   wire n25684;
   wire n25685;
   wire n25686;
   wire n25687;
   wire n25688;
   wire n25689;
   wire n25690;
   wire n25691;
   wire n25692;
   wire n25693;
   wire n25694;
   wire n25695;
   wire n25696;
   wire n25697;
   wire n25698;
   wire n25699;
   wire n25700;
   wire n25701;
   wire n25702;
   wire n25703;
   wire n25704;
   wire n25705;
   wire n25706;
   wire n25707;
   wire n25708;
   wire n25709;
   wire n25710;
   wire n25711;
   wire n25712;
   wire n25713;
   wire n25714;
   wire n25715;
   wire n25716;
   wire n25717;
   wire n25718;
   wire n25719;
   wire n25720;
   wire n25721;
   wire n25722;
   wire n25723;
   wire n25724;
   wire n25725;
   wire n25726;
   wire n25727;
   wire n25728;
   wire n25729;
   wire n25730;
   wire n25731;
   wire n25732;
   wire n25733;
   wire n25734;
   wire n25735;
   wire n25736;
   wire n25737;
   wire n25738;
   wire n25739;
   wire n25740;
   wire n25741;
   wire n25742;
   wire n25743;
   wire n25744;
   wire n25745;
   wire n25746;
   wire n25747;
   wire n25748;
   wire n25749;
   wire n25750;
   wire n25751;
   wire n25752;
   wire n25753;
   wire n25754;
   wire n25755;
   wire n25756;
   wire n25757;
   wire n25758;
   wire n25759;
   wire n25760;
   wire n25761;
   wire n25762;
   wire n25763;
   wire n25764;
   wire n25765;
   wire n25766;
   wire n25767;
   wire n25768;
   wire n25769;
   wire n25770;
   wire n25771;
   wire n25772;
   wire n25773;
   wire n25774;
   wire n25775;
   wire n25776;
   wire n25777;
   wire n25778;
   wire n25779;
   wire n25780;
   wire n25781;
   wire n25782;
   wire n25783;
   wire n25784;
   wire n25785;
   wire n25786;
   wire n25787;
   wire n25788;
   wire n25789;
   wire n25790;
   wire n25791;
   wire n25792;
   wire n25793;
   wire n25794;
   wire n25795;
   wire n25796;
   wire n25797;
   wire n25798;
   wire n25799;
   wire n25800;
   wire n25801;
   wire n25802;
   wire n25803;
   wire n25804;
   wire n25805;
   wire n25806;
   wire n25807;
   wire n25808;
   wire n25809;
   wire n25810;
   wire n25811;
   wire n25812;
   wire n25813;
   wire n25814;
   wire n25815;
   wire n25816;
   wire n25817;
   wire n25818;
   wire n25819;
   wire n25820;
   wire n25821;
   wire n25822;
   wire n25823;
   wire n25824;
   wire n25825;
   wire n25826;
   wire n25827;
   wire n25828;
   wire n25829;
   wire n25830;
   wire n25831;
   wire n25832;
   wire n25833;
   wire n25834;
   wire n25835;
   wire n25836;
   wire n25837;
   wire n25838;
   wire n25839;
   wire n25840;
   wire n25841;
   wire n25842;
   wire n25843;
   wire n25844;
   wire n25845;
   wire n25846;
   wire n25847;
   wire n25848;
   wire n25849;
   wire n25850;
   wire n25851;
   wire n25852;
   wire n25853;
   wire n25854;
   wire n25855;
   wire n25856;
   wire n25857;
   wire n25858;
   wire n25859;
   wire n25860;
   wire n25861;
   wire n25862;
   wire n25863;
   wire n25864;
   wire n25865;
   wire n25866;
   wire n25867;
   wire n25868;
   wire n25869;
   wire n25870;
   wire n25871;
   wire n25872;
   wire n25873;
   wire n25874;
   wire n25875;
   wire n25876;
   wire n25877;
   wire n25878;
   wire n25879;
   wire n25880;
   wire n25881;
   wire n25882;
   wire n25883;
   wire n25884;
   wire n25885;
   wire n25886;
   wire n25887;
   wire n25888;
   wire n25889;
   wire n25890;
   wire n25891;
   wire n25892;
   wire n25893;
   wire n25894;
   wire n25895;
   wire n25896;
   wire n25897;
   wire n25898;
   wire n25899;
   wire n25900;
   wire n25901;
   wire n25902;
   wire n25903;
   wire n25904;
   wire n25905;
   wire n25906;
   wire n25907;
   wire n25908;
   wire n25909;
   wire n25910;
   wire n25911;
   wire n25912;
   wire n25913;
   wire n25914;
   wire n25915;
   wire n25916;
   wire n25917;
   wire n25918;
   wire n25919;
   wire n25920;
   wire n25921;
   wire n25922;
   wire n25923;
   wire n25924;
   wire n25925;
   wire n25926;
   wire n25927;
   wire n25928;
   wire n25929;
   wire n25930;
   wire n25931;
   wire n25932;
   wire n25933;
   wire n25934;
   wire n25935;
   wire n25936;
   wire n25937;
   wire n25938;
   wire n25939;
   wire n25940;
   wire n25941;
   wire n25942;
   wire n25943;
   wire n25944;
   wire n25945;
   wire n25946;
   wire n25947;
   wire n25948;
   wire n25949;
   wire n25950;
   wire n25951;
   wire n25952;
   wire n25953;
   wire n25954;
   wire n25955;
   wire n25956;
   wire n25957;
   wire n25958;
   wire n25959;
   wire n25960;
   wire n25961;
   wire n25962;
   wire n25963;
   wire n25964;
   wire n25965;
   wire n25966;
   wire n25967;
   wire n25968;
   wire n25969;
   wire n25970;
   wire n25971;
   wire n25972;
   wire n25973;
   wire n25974;
   wire n25975;
   wire n25976;
   wire n25977;
   wire n25978;
   wire n25979;
   wire n25980;
   wire n25981;
   wire n25982;
   wire n25983;
   wire n25984;
   wire n25985;
   wire n25986;
   wire n25987;
   wire n25988;
   wire n25989;
   wire n25990;
   wire n25991;
   wire n25992;
   wire n25993;
   wire n25994;
   wire n25995;
   wire n25997;
   wire n25998;
   wire n25999;
   wire n26000;
   wire n26003;
   wire n26006;
   wire n26008;
   wire n26009;
   wire n26010;
   wire n26011;
   wire n26012;
   wire n26013;
   wire n26014;
   wire n26015;
   wire n26016;
   wire n26017;
   wire n26018;
   wire n26019;
   wire n26020;
   wire n26021;
   wire n26022;
   wire n26023;
   wire n26024;
   wire n26025;
   wire n26026;
   wire n26027;
   wire n26028;

   assign store_meter_ack_non_partner = 1'b0 ;
   assign store_meter_ack_partner = 1'b0 ;
   assign external_interrupt = 1'b0 ;

   in01f01 FE_OFC2735_n21666 (.o(FE_OFN25981_n21666),
	.a(FE_OFN25974_n21666));
   in01f01 FE_OFC2734_n21666 (.o(FE_OFN25980_n21666),
	.a(FE_OFN25974_n21666));
   in01f01 FE_OFC2733_n21666 (.o(FE_OFN25979_n21666),
	.a(FE_OFN25974_n21666));
   in01f01 FE_OFC2732_n21666 (.o(FE_OFN25978_n21666),
	.a(FE_OFN25974_n21666));
   in01f01 FE_OFC2731_n21666 (.o(FE_OFN25977_n21666),
	.a(FE_OFN25974_n21666));
   in01f01 FE_OFC2730_n21666 (.o(FE_OFN25976_n21666),
	.a(FE_OFN25973_n21666));
   in01f01 FE_OFC2729_n21666 (.o(FE_OFN25975_n21666),
	.a(FE_OFN25973_n21666));
   in01f01 FE_OFC2728_n21666 (.o(FE_OFN25974_n21666),
	.a(n21666));
   in01f01 FE_OFC2727_n21666 (.o(FE_OFN25973_n21666),
	.a(n21666));
   in01f06 FE_OFC2726_n20135 (.o(FE_OFN25972_n20135),
	.a(FE_OFN25971_n20135));
   in01f03 FE_OFC2725_n20135 (.o(FE_OFN25971_n20135),
	.a(n20135));
   in01f40 FE_OCPC2610_n19306_dup (.o(FE_RN_69),
	.a(FE_OFN24736_n19306));
   na04f03 FE_RC_130_0 (.o(n24093),
	.a(n24090),
	.b(n24091),
	.c(n24089),
	.d(n24092));
   oa12m02 FE_RC_129_0 (.o(FE_OFN643_dataOut_E_17),
	.a(n24411),
	.b(FE_OFN219_n24645),
	.c(FE_OFN25892_n25395));
   oa12m02 FE_RC_128_0 (.o(FE_OFN787_dataOut_W_21),
	.a(n24571),
	.b(FE_OFN233_n24719),
	.c(FE_OFN394_n19446));
   ao22f01 FE_RC_127_0 (.o(n21135),
	.a(n23949),
	.b(n19056),
	.c(FE_OFN138_n23948),
	.d(n19054));
   in01f02 FE_OCPC2724_FE_OFN141_n23964 (.o(FE_OFN142_n23964),
	.a(FE_OFN141_n23964));
   in01f06 FE_OCPC2723_n24342 (.o(FE_OCPN25970_n24342),
	.a(n24342));
   in01f08 FE_OCPC2722_n24342 (.o(FE_OCPN25841_n24342),
	.a(n24342));
   in01f04 FE_OCPC2721_n24342 (.o(FE_OCPN25835_n24342),
	.a(n24342));
   in01f06 FE_OCPC2720_n24342 (.o(n19654),
	.a(n24342));
   in01f03 FE_OCPC2719_n24342 (.o(FE_OCPN25838_n24342),
	.a(n24342));
   in01f08 FE_OCPC2718_n24342 (.o(FE_OCPN25839_n24342),
	.a(n24342));
   in01f08 FE_OCPC2717_n24342 (.o(FE_OCPN25830_n),
	.a(n24342));
   in01f10 FE_OCPC2716_n24342 (.o(FE_OCPN25836_n24342),
	.a(n24342));
   na04m04 FE_RC_126_0 (.o(n24230),
	.a(n24229),
	.b(n24226),
	.c(n24228),
	.d(n24227));
   oa12m02 FE_RC_125_0 (.o(FE_OFN883_dataOut_P_0),
	.a(n24661),
	.b(FE_OFN239_n24739),
	.c(FE_OFN524_n24728));
   ao22f01 FE_RC_124_0 (.o(n24417),
	.a(FE_OFN237_n24730),
	.b(FE_OFN44_n19054),
	.c(FE_OFN528_n24732),
	.d(n19057));
   oa12m02 FE_RC_123_0 (.o(FE_OFN986_dataOut_E_18),
	.a(n24403),
	.b(n24759),
	.c(FE_OFN25895_n25395));
   oa12m02 FE_RC_122_0 (.o(FE_OFN1032_dataOut_W_18),
	.a(n24547),
	.b(n24759),
	.c(FE_OFN25878_n19446));
   in01f01 FE_RC_121_0 (.o(FE_RN_54_0),
	.a(n25515));
   in01f01 FE_RC_120_0 (.o(FE_RN_55_0),
	.a(n25513));
   in01f01 FE_RC_119_0 (.o(FE_RN_56_0),
	.a(n25514));
   in01f01 FE_RC_118_0 (.o(dataOut_N_51_),
	.a(FE_RN_57_0));
   no03f02 FE_RC_117_0 (.o(FE_RN_57_0),
	.a(FE_RN_56_0),
	.b(FE_RN_55_0),
	.c(FE_RN_54_0));
   oa12m02 FE_RC_116_0 (.o(FE_OFN1058_dataOut_P_12),
	.a(n24592),
	.b(n24593),
	.c(n24728));
   oa12m02 FE_RC_115_0 (.o(FE_OFN799_dataOut_W_13),
	.a(n24539),
	.b(n24606),
	.c(FE_OFN25878_n19446));
   ao22f01 FE_RC_114_0 (.o(n24117),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__11_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__11_));
   oa12m02 FE_RC_113_0 (.o(FE_OFN1008_dataOut_S_18),
	.a(n24674),
	.b(n24759),
	.c(FE_OFN25652_n25499));
   ao22m02 FE_RC_112_0 (.o(n21757),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__8_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__8_));
   in01f04 FE_OCPC2715_FE_OFN143_n23991 (.o(FE_OFN144_n23991),
	.a(FE_OFN143_n23991));
   in01f01 FE_RC_111_0 (.o(FE_RN_51_0),
	.a(n21794));
   in01f01 FE_RC_110_0 (.o(FE_RN_52_0),
	.a(n21793));
   no02f02 FE_RC_109_0 (.o(FE_RN_53_0),
	.a(FE_RN_52_0),
	.b(FE_RN_51_0));
   na03f02 FE_RC_108_0 (.o(n21801),
	.a(n21791),
	.b(n21792),
	.c(FE_RN_53_0));
   oa12m02 FE_RC_107_0 (.o(FE_OFN659_dataOut_E_0),
	.a(n24371),
	.b(FE_OFN239_n24739),
	.c(FE_OFN25895_n25395));
   oa12m02 FE_RC_106_0 (.o(FE_OFN998_dataOut_E_5),
	.a(n21325),
	.b(n23982),
	.c(FE_OFN25892_n25395));
   ao22m02 FE_RC_105_0 (.o(n24251),
	.a(FE_OCPN25840_n24342),
	.b(proc_input_NIB_storage_data_f_0__14_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__14_));
   na02f20 U23427_dup (.o(FE_RN_68),
	.a(n18676),
	.b(n18675));
   ao22f02 FE_RC_104_0 (.o(n20008),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__22_),
	.c(FE_OCPN25953_n18039),
	.d(proc_input_NIB_storage_data_f_10__22_));
   no02f20 U21678_dup (.o(FE_RN_67),
	.a(n19053),
	.b(n19052));
   ao22f01 FE_RC_103_0 (.o(n20010),
	.a(FE_RN_35),
	.b(proc_input_NIB_storage_data_f_12__22_),
	.c(FE_OFN191_n24454),
	.d(proc_input_NIB_storage_data_f_13__22_));
   in01f20 FE_OFC1798_n18815_dup (.o(FE_RN_66),
	.a(n18974));
   na02f10 U21213_dup (.o(FE_RN_65),
	.a(n18916),
	.b(n18915));
   no02f40 U23965_dup2 (.o(FE_RN_64),
	.a(n18827),
	.b(FE_OCPN25899_west_input_NIB_head_ptr_f_0));
   in01f01 FE_RC_102_0 (.o(FE_RN_48_0),
	.a(n25483));
   no02f02 FE_RC_100_0 (.o(FE_RN_50_0),
	.a(n25972),
	.b(FE_RN_48_0));
   na02f06 FE_RC_99_0 (.o(n25484),
	.a(thanksIn_P),
	.b(FE_RN_50_0));
   ao22f10 FE_RC_98_0 (.o(n18901),
	.a(n23993),
	.b(myChipID_f_4_),
	.c(n23587),
	.d(n19575));
   in01f03 FE_RC_97_0 (.o(FE_RN_45_0),
	.a(n19805));
   in01f04 FE_RC_96_0 (.o(FE_RN_46_0),
	.a(n19806));
   no02f06 FE_RC_95_0 (.o(FE_RN_47_0),
	.a(FE_RN_46_0),
	.b(FE_RN_45_0));
   no02f06 FE_RC_94_0 (.o(n19807),
	.a(n19804),
	.b(FE_RN_47_0));
   in01f10 FE_OFC1207_n18683_dup (.o(FE_RN_63),
	.a(FE_RN_40));
   in01f40 FE_OCPC2584_n18648_dup (.o(FE_RN_62),
	.a(n24964));
   na03f06 FE_RC_93_0 (.o(n18458),
	.a(n20523),
	.b(n20521),
	.c(n25339));
   no03f02 FE_RC_92_0 (.o(n18187),
	.a(n18458),
	.b(n18197),
	.c(n18199));
   ao22f08 FE_RC_91_0 (.o(n19988),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__25_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__25_));
   ao22f08 FE_RC_90_0 (.o(n19999),
	.a(FE_OFN28_n18974),
	.b(west_input_NIB_storage_data_f_0__23_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__23_));
   in01f01 FE_RC_89_0 (.o(FE_RN_42_0),
	.a(FE_OFN25596_reset));
   in01f04 FE_RC_88_0 (.o(FE_RN_43_0),
	.a(n25339));
   no02f06 FE_RC_87_0 (.o(FE_RN_44_0),
	.a(FE_RN_43_0),
	.b(FE_RN_42_0));
   na03f06 FE_RC_86_0 (.o(n25322),
	.a(n25324),
	.b(n25321),
	.c(FE_RN_44_0));
   na04f06 FE_RC_85_0 (.o(n20458),
	.a(n25172),
	.b(n20530),
	.c(n25170),
	.d(n20514));
   na02f10 U20207_dup (.o(FE_RN_61),
	.a(n19264),
	.b(n19263));
   na03f20 U23581_dup (.o(FE_RN_60),
	.a(n18582),
	.b(n18581),
	.c(n18580));
   na02f20 U23923_dup (.o(FE_RN_44),
	.a(n18678),
	.b(n18677));
   ao22f10 FE_RC_84_0 (.o(n19153),
	.a(FE_OFN48_n19193),
	.b(north_input_NIB_storage_data_f_3__52_),
	.c(FE_OFN24773_n19075),
	.d(north_input_NIB_storage_data_f_0__52_));
   ao22f08 FE_RC_83_0 (.o(n17919),
	.a(FE_OFN156_n24129),
	.b(proc_input_NIB_storage_data_f_1__37_),
	.c(FE_OFN25637_n19595),
	.d(proc_input_NIB_storage_data_f_15__37_));
   na02f04 FE_RC_82_0 (.o(FE_RN_39_0),
	.a(n20064),
	.b(n20063));
   na02f04 FE_RC_81_0 (.o(FE_RN_40_0),
	.a(n20066),
	.b(n20065));
   in01f06 FE_RC_80_0 (.o(n20072),
	.a(FE_RN_41_0));
   no02f06 FE_RC_79_0 (.o(FE_RN_41_0),
	.a(FE_RN_40_0),
	.b(FE_RN_39_0));
   ao22f08 FE_RC_78_0 (.o(n19581),
	.a(FE_OCPN25838_n24342),
	.b(proc_input_NIB_storage_data_f_0__61_),
	.c(FE_RN_59),
	.d(proc_input_NIB_storage_data_f_4__61_));
   in01f02 FE_OCPC2714_n19500 (.o(FE_OCPN25969_n19500),
	.a(FE_OFN25675_n17777));
   in01f20 FE_OCPC2713_n19500 (.o(FE_OCPN25968_n19500),
	.a(FE_OFN25675_n17777));
   in01f02 FE_OCPC2712_n19500 (.o(FE_OCPN25967_n19500),
	.a(FE_OFN25675_n17777));
   in01f08 FE_OCPC2711_n19500 (.o(FE_OFN25688_n19500),
	.a(FE_OFN25675_n17777));
   in01f06 FE_OCPC2710_n19500 (.o(n21739),
	.a(FE_OFN25675_n17777));
   in01f02 FE_OCPC2709_n19500 (.o(FE_OFN25686_n19500),
	.a(FE_OFN25675_n17777));
   in01f02 FE_OCPC2708_n19500 (.o(FE_RN_35),
	.a(FE_OFN25675_n17777));
   in01f01 FE_OCPC2707_n19500 (.o(FE_OCPN25832_n19500),
	.a(FE_OFN25675_n17777));
   in01f02 FE_OCPC2706_n19500 (.o(FE_RN_54),
	.a(FE_OFN25675_n17777));
   in01f08 FE_OCPC2705_n19500 (.o(n17747),
	.a(FE_OFN25675_n17777));
   in01f20 FE_OCPC2704_n19500 (.o(FE_OFN25675_n17777),
	.a(n19500));
   in01f10 FE_OFC2264_n19508_dup (.o(FE_RN_59),
	.a(FE_OFN25606_n19508));
   ao22f08 FE_RC_77_0 (.o(n19676),
	.a(n24060),
	.b(proc_input_NIB_storage_data_f_9__49_),
	.c(FE_OCPN25949_n18039),
	.d(proc_input_NIB_storage_data_f_10__49_));
   in01f08 FE_OCPC2703_proc_input_NIB_head_ptr_f_2 (.o(FE_OCPN25966_proc_input_NIB_head_ptr_f_2),
	.a(proc_input_NIB_head_ptr_f_2_));
   in01f01 FE_OCPC2702_proc_input_NIB_head_ptr_f_2 (.o(FE_OCPN25965_proc_input_NIB_head_ptr_f_2),
	.a(proc_input_NIB_head_ptr_f_2_));
   in01f20 FE_OCPC2701_proc_input_NIB_head_ptr_f_2 (.o(n19502),
	.a(proc_input_NIB_head_ptr_f_2_));
   oa22f10 FE_RC_76_0 (.o(n19650),
	.a(n19634),
	.b(n19635),
	.c(n23318),
	.d(n19633));
   ao12f06 FE_RC_75_0 (.o(n18711),
	.a(n18351),
	.b(FE_OFN24741_n18683),
	.c(south_input_NIB_storage_data_f_1__34_));
   ao22f06 U21927_dup (.o(FE_RN_58),
	.a(FE_OCPN25810_n18959),
	.b(west_input_NIB_storage_data_f_3__44_),
	.c(FE_OFN27_n18974),
	.d(west_input_NIB_storage_data_f_0__44_));
   in01f20 FE_OCPC2604_n19306_dup (.o(FE_RN_57),
	.a(n19306));
   na02f10 U23911_dup (.o(FE_RN_56),
	.a(n18662),
	.b(n18661));
   na04f06 FE_RC_74_0 (.o(n19117),
	.a(n19246),
	.b(n20168),
	.c(n20167),
	.d(n19245));
   in01f10 FE_OFC1208_n18683_dup (.o(FE_RN_55),
	.a(FE_RN_40));
   na02f06 FE_RC_73_0 (.o(FE_RN_36_0),
	.a(FE_OCPN25901_west_input_NIB_head_ptr_f_0),
	.b(n18824));
   na02f03 FE_RC_72_0 (.o(FE_RN_37_0),
	.a(n18825),
	.b(west_input_NIB_head_ptr_f_0_));
   in01f08 FE_RC_71_0 (.o(n21342),
	.a(FE_RN_38_0));
   na02f06 FE_RC_70_0 (.o(FE_RN_38_0),
	.a(FE_RN_37_0),
	.b(FE_RN_36_0));
   ao22f10 FE_RC_69_0 (.o(n18649),
	.a(n18061),
	.b(south_input_NIB_storage_data_f_1__63_),
	.c(n19973),
	.d(south_input_NIB_storage_data_f_2__63_));
   in01f20 FE_OFC1875_n19225_dup (.o(FE_RN_10),
	.a(n19225));
   in01f40 FE_OCPC2700_n19530 (.o(n24454),
	.a(n19530));
   in01f40 FE_OCPC2699_n21739 (.o(FE_OFN24803_n19500),
	.a(FE_OFN25675_n17777));
   in01f02 FE_OCPC2698_n18039 (.o(FE_OCPN25964_n18039),
	.a(n18036));
   in01f02 FE_OCPC2697_n18039 (.o(FE_OCPN25963_n18039),
	.a(n18036));
   in01f10 FE_OCPC2696_n18039 (.o(FE_OCPN25962_n18039),
	.a(n18036));
   in01f02 FE_OCPC2695_n18039 (.o(FE_OCPN25961_n18039),
	.a(n18036));
   in01f04 FE_OCPC2694_n18039 (.o(FE_OCPN25960_n18039),
	.a(n18036));
   in01f06 FE_OCPC2693_n18039 (.o(FE_OCPN25959_n18039),
	.a(n18036));
   in01f02 FE_OCPC2692_n18039 (.o(FE_OCPN25958_n18039),
	.a(n18036));
   in01f06 FE_OCPC2691_n18039 (.o(FE_OCPN25957_n18039),
	.a(n18036));
   in01f02 FE_OCPC2690_n18039 (.o(FE_OCPN25956_n18039),
	.a(n18036));
   in01f02 FE_OCPC2689_n18039 (.o(FE_OCPN25955_n18039),
	.a(n18036));
   in01f10 FE_OCPC2688_n18039 (.o(FE_OCPN25954_n18039),
	.a(n18036));
   in01f01 FE_OCPC2687_n18039 (.o(FE_OCPN25953_n18039),
	.a(n18036));
   in01f04 FE_OCPC2686_n18039 (.o(FE_OCPN25952_n18039),
	.a(n18036));
   in01f01 FE_OCPC2685_n18039 (.o(FE_OCPN25951_n18039),
	.a(n18036));
   in01f03 FE_OCPC2684_n18039 (.o(FE_OCPN25950_n18039),
	.a(n18036));
   in01f04 FE_OCPC2683_n18039 (.o(FE_OCPN25949_n18039),
	.a(n18036));
   in01f02 FE_OCPC2682_n18039 (.o(n18035),
	.a(n18036));
   in01f01 FE_OCPC2681_n18039 (.o(n18034),
	.a(n18036));
   in01f02 FE_OCPC2680_n18039 (.o(n18051),
	.a(n18036));
   in01f01 FE_OCPC2679_n18039 (.o(FE_OFN25668_n18038),
	.a(n18036));
   in01f02 FE_OCPC2678_n18039 (.o(n18037),
	.a(n18036));
   in01f04 FE_OCPC2677_n18039 (.o(n18038),
	.a(n18036));
   in01f20 FE_OCPC2676_n18039 (.o(n18036),
	.a(n18039));
   in01f20 FE_OFC2260_n19508_dup (.o(FE_RN_53),
	.a(n19508));
   in01f02 FE_RC_68_0 (.o(FE_RN_33_0),
	.a(n20094));
   in01f02 FE_RC_67_0 (.o(FE_RN_34_0),
	.a(n20093));
   no02f06 FE_RC_66_0 (.o(FE_RN_35_0),
	.a(FE_RN_34_0),
	.b(FE_RN_33_0));
   na02f06 FE_RC_65_0 (.o(n20103),
	.a(FE_RN_17_0),
	.b(FE_RN_35_0));
   no03f04 FE_RC_64_0 (.o(n20461),
	.a(n20456),
	.b(n20453),
	.c(FE_RN_2_0));
   in01f01 FE_OCPC2675_n19595 (.o(FE_OCPN25948_n19595),
	.a(FE_RN_34));
   in01f40 FE_OCPC2674_n19595 (.o(FE_OCPN25947_n19595),
	.a(FE_RN_34));
   in01f02 FE_OCPC2673_n19595 (.o(n19544),
	.a(FE_RN_34));
   in01f06 FE_OCPC2672_n19595 (.o(FE_OFN25635_n19595),
	.a(FE_RN_34));
   in01f02 FE_OCPC2671_n19595 (.o(FE_OFN25634_n19595),
	.a(FE_RN_34));
   in01f01 FE_OCPC2670_n19595 (.o(n20097),
	.a(FE_RN_34));
   in01f02 FE_OCPC2669_n19595 (.o(FE_OFN25633_n19595),
	.a(FE_RN_34));
   in01f01 FE_OCPC2668_n19595 (.o(FE_OFN25632_n19595),
	.a(FE_RN_34));
   in01f03 FE_OCPC2667_n19595 (.o(n17780),
	.a(FE_RN_34));
   in01f08 FE_OCPC2666_n19595 (.o(FE_OFN25637_n19595),
	.a(FE_RN_34));
   in01f02 FE_OCPC2665_n19595 (.o(FE_RN_50),
	.a(FE_RN_34));
   in01f03 FE_OCPC2664_n19595 (.o(FE_OFN25636_n19595),
	.a(FE_RN_34));
   in01f01 FE_OCPC2663_n19595 (.o(n24065),
	.a(FE_RN_34));
   in01f20 FE_OCPC2662_n19595 (.o(FE_RN_34),
	.a(n19595));
   in01f10 FE_OFC1802_n19505_dup (.o(FE_RN_52),
	.a(n19505));
   in01f03 FE_OFC2036_n21747_dup (.o(FE_RN_51),
	.a(FE_RN_48));
   no03m04 FE_RC_63_0 (.o(n20766),
	.a(n19919),
	.b(n19921),
	.c(n19920));
   in01f40 FE_OCPC2627_n19550_dup (.o(FE_RN_49),
	.a(n19550));
   in01f40 FE_OCPC2661_n21747 (.o(FE_OFN161_n24129),
	.a(n21747));
   ao22f10 FE_RC_62_0 (.o(n19612),
	.a(FE_OCPN25947_n19595),
	.b(proc_input_NIB_storage_data_f_15__60_),
	.c(n17754),
	.d(proc_input_NIB_storage_data_f_3__60_));
   ao22f20 FE_RC_61_0 (.o(n19172),
	.a(FE_OFN96_n21865),
	.b(north_input_NIB_storage_data_f_2__54_),
	.c(FE_OFN25610_n19071),
	.d(north_input_NIB_storage_data_f_1__54_));
   na02f40 U23443_dup (.o(FE_RN_48),
	.a(FE_OFN24793_n17934),
	.b(FE_OCPN25946_n19501));
   in01f01 FE_RC_60_0 (.o(FE_RN_30_0),
	.a(n25167));
   in01f02 FE_RC_59_0 (.o(FE_RN_31_0),
	.a(n25184));
   no02f04 FE_RC_58_0 (.o(FE_RN_32_0),
	.a(FE_RN_31_0),
	.b(FE_RN_30_0));
   no02f02 FE_RC_57_0 (.o(west_output_control_N469),
	.a(n25166),
	.b(FE_RN_32_0));
   in01f10 FE_OCPC2407_n18959_dup (.o(FE_RN_47),
	.a(n18959));
   in01f10 U23903_dup (.o(FE_RN_46),
	.a(n18651));
   in01f40 FE_OFC1761_north_input_NIB_head_ptr_f_1_dup (.o(FE_RN_45),
	.a(north_input_NIB_head_ptr_f_1_));
   ao22f10 FE_RC_56_0 (.o(n18650),
	.a(n24473),
	.b(south_input_NIB_storage_data_f_3__63_),
	.c(FE_OFN24744_n18648),
	.d(south_input_NIB_storage_data_f_0__63_));
   ao22f20 FE_RC_55_0 (.o(n18916),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__62_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__62_));
   oa22f10 FE_RC_54_0 (.o(n18579),
	.a(n23995),
	.b(FE_OFN53_n19355),
	.c(n21407),
	.d(n19347));
   no03f20 U23907_dup (.o(FE_RN_43),
	.a(n18659),
	.b(n18658),
	.c(n18657));
   in01f10 FE_OFC1805_south_input_NIB_head_ptr_f_1_dup1 (.o(FE_RN_42),
	.a(south_input_NIB_head_ptr_f_1_));
   no02f80 U23588_dup (.o(FE_RN_41),
	.a(south_input_NIB_head_ptr_f_0_),
	.b(FE_RN_30));
   na02f40 U23604_dup (.o(FE_RN_40),
	.a(FE_OFN15_south_input_NIB_head_ptr_f_1),
	.b(south_input_NIB_head_ptr_f_0_));
   no04f06 FE_RC_53_0 (.o(n20223),
	.a(n20218),
	.b(n20219),
	.c(n20220),
	.d(n18099));
   na02f10 U21470_dup (.o(FE_RN_39),
	.a(n18002),
	.b(n17995));
   in01f08 FE_OCPC2447_n21745_dup (.o(FE_RN_38),
	.a(FE_RN_15));
   na02f40 U23454_dup (.o(FE_RN_37),
	.a(n19502),
	.b(proc_input_NIB_head_ptr_f_3_));
   na03f20 U23506_dup (.o(FE_RN_36),
	.a(n18311),
	.b(n18309),
	.c(n18306));
   na03f04 FE_RC_52_0 (.o(n25046),
	.a(n25469),
	.b(n25470),
	.c(proc_input_NIB_elements_in_array_f_2_));
   ao22f10 FE_RC_51_0 (.o(n19614),
	.a(FE_OCPN25962_n18039),
	.b(proc_input_NIB_storage_data_f_10__60_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__60_));
   in01f20 FE_OCPC2660_n19501 (.o(FE_OCPN25946_n19501),
	.a(FE_OCPN25931_n19501));
   in01f20 FE_OCPC2659_n19501 (.o(FE_OCPN25932_n19501),
	.a(FE_OCPN25931_n19501));
   in01f20 FE_OCPC2658_n19501 (.o(FE_OCPN25931_n19501),
	.a(n19501));
   in01f10 FE_OCPC2657_n19501 (.o(n18533),
	.a(n19501));
   in01f08 FE_OFC2117_n19655_dup (.o(FE_RN_33),
	.a(FE_OFN25671_n19655));
   in01f01 FE_RC_50_0 (.o(FE_RN_27_0),
	.a(n25064));
   in01f02 FE_RC_49_0 (.o(FE_RN_28_0),
	.a(FE_OFN570_n25395));
   no02f02 FE_RC_48_0 (.o(FE_RN_29_0),
	.a(FE_RN_28_0),
	.b(FE_RN_27_0));
   na02f02 FE_RC_47_0 (.o(n25066),
	.a(n25396),
	.b(FE_RN_29_0));
   na04f20 FE_RC_46_0 (.o(n18120),
	.a(n17949),
	.b(n17948),
	.c(n17947),
	.d(n17941));
   in01f04 FE_RC_45_0 (.o(FE_RN_24_0),
	.a(proc_input_NIB_storage_data_f_11__53_));
   in01f04 FE_RC_44_0 (.o(FE_RN_25_0),
	.a(FE_OCPN25920_n19547));
   no02f06 FE_RC_43_0 (.o(FE_RN_26_0),
	.a(FE_RN_25_0),
	.b(FE_RN_24_0));
   no02f08 FE_RC_42_0 (.o(n19665),
	.a(FE_RN_26_0),
	.b(n17932));
   no04f06 FE_RC_41_0 (.o(n25107),
	.a(n25104),
	.b(n25103),
	.c(n25105),
	.d(n25106));
   in01f20 FE_OFC1800_n18815_dup (.o(FE_RN_32),
	.a(n18837));
   in01f10 FE_OCPC2656_n23612 (.o(n17797),
	.a(n23612));
   in01f10 FE_OCPC2655_n19071 (.o(n24364),
	.a(FE_OFN177_n24364));
   in01f40 FE_OCPC2654_n19071 (.o(FE_OFN25610_n19071),
	.a(FE_OFN177_n24364));
   in01f20 FE_OCPC2653_n19071 (.o(FE_OFN178_n24364),
	.a(FE_OFN177_n24364));
   in01f20 FE_OCPC2652_n19071 (.o(FE_OFN177_n24364),
	.a(n19071));
   in01f03 FE_OCPC2651_n19071 (.o(n19223),
	.a(n19071));
   in01f04 FE_OCPC2650_n19071 (.o(FE_OFN176_n24364),
	.a(n19071));
   in01f02 FE_OCPC2649_n24965 (.o(FE_OCPN25945_n24965),
	.a(n24965));
   in01f06 FE_OCPC2648_n24965 (.o(FE_OCPN25944_n24965),
	.a(n24965));
   in01f06 FE_OCPC2647_n24965 (.o(FE_OCPN25943_n24965),
	.a(n24965));
   in01f01 FE_OCPC2646_n24965 (.o(FE_OCPN25942_n24965),
	.a(n24965));
   in01f08 FE_OCPC2645_n24965 (.o(FE_OCPN25941_n24965),
	.a(n24965));
   in01f01 FE_OCPC2644_n24965 (.o(FE_OCPN25940_n24965),
	.a(n24965));
   in01f06 FE_OCPC2643_n24965 (.o(FE_OCPN25939_n24965),
	.a(n24965));
   in01f01 FE_OCPC2642_n24965 (.o(FE_OCPN25938_n24965),
	.a(n24965));
   in01f01 FE_OCPC2641_n24965 (.o(FE_OCPN25937_n24965),
	.a(n24965));
   in01f01 FE_OCPC2640_n24965 (.o(FE_OCPN25936_n24965),
	.a(n24965));
   in01f01 FE_OCPC2639_n24965 (.o(FE_OCPN25935_n24965),
	.a(n24965));
   in01f02 FE_OCPC2638_n24965 (.o(FE_RN_13),
	.a(n24965));
   in01f01 FE_OCPC2637_n24965 (.o(FE_OFN24791_n24965),
	.a(n24965));
   in01f01 FE_OCPC2636_n24965 (.o(FE_OFN24788_n24965),
	.a(n24965));
   in01f40 FE_OCPC2635_n24965 (.o(n24473),
	.a(n24965));
   na02f20 U24007_dup (.o(FE_RN_25),
	.a(n18887),
	.b(n18886));
   no03f08 FE_RC_40_0 (.o(n21426),
	.a(n18958),
	.b(n18956),
	.c(n18957));
   no02f80 U23979_dup (.o(FE_RN_31),
	.a(west_input_NIB_head_ptr_f_1_),
	.b(FE_OCPN25900_west_input_NIB_head_ptr_f_0));
   in01f40 FE_OFC1805_south_input_NIB_head_ptr_f_1_dup (.o(FE_RN_30),
	.a(south_input_NIB_head_ptr_f_1_));
   in01f10 FE_OCPC2634_n19914 (.o(FE_OFN25661_n19914),
	.a(FE_OFN25664_n19914));
   in01f40 FE_OCPC2633_n19914 (.o(FE_OFN25659_n19914),
	.a(FE_OFN25663_n19914));
   in01f20 FE_OCPC2632_n19914 (.o(FE_OFN25662_n19914),
	.a(FE_OFN25663_n19914));
   in01f10 FE_OCPC2631_n19914 (.o(n24359),
	.a(FE_OFN25663_n19914));
   in01f08 FE_OCPC2630_n19914 (.o(FE_OFN25664_n19914),
	.a(n19914));
   in01f40 FE_OCPC2628_n19914 (.o(FE_OFN25663_n19914),
	.a(n19914));
   in01f20 FE_OCPC2627_n19550 (.o(n18077),
	.a(n19550));
   in01f40 FE_OCPC2626_n19980 (.o(FE_OFN28_n18974),
	.a(n19980));
   in01f40 FE_OCPC2625_n19498 (.o(FE_OFN20_n17779),
	.a(FE_OFN25640_n19498));
   in01f10 FE_OCPC2624_n19498 (.o(n17779),
	.a(FE_OFN25640_n19498));
   in01f20 FE_OCPC2623_n19498 (.o(FE_OFN25640_n19498),
	.a(n19498));
   in01f10 FE_OCPC2622_n24342 (.o(FE_OCPN25934_n24342),
	.a(FE_OCPN25933_n24342));
   in01f40 FE_OCPC2621_n24342 (.o(FE_OCPN25933_n24342),
	.a(n24342));
   in01f40 FE_OCPC2613_n19504 (.o(n19769),
	.a(FE_OFN25643_n19504));
   in01f40 FE_OCPC2612_n19504 (.o(FE_OFN25644_n19504),
	.a(FE_OFN25643_n19504));
   in01f20 FE_OCPC2611_n19504 (.o(FE_OFN25643_n19504),
	.a(n19504));
   in01f40 FE_OCPC2610_n19306 (.o(FE_OCPN25813_FE_OFN24735_n19306),
	.a(FE_OFN24736_n19306));
   in01f02 FE_OCPC2609_n19306 (.o(FE_OFN24737_n19306),
	.a(FE_RN_57));
   in01f02 FE_OCPC2608_n19306 (.o(FE_OFN24732_n19306),
	.a(FE_RN_57));
   in01f04 FE_OCPC2607_n19306 (.o(FE_OCPN25906_n19306),
	.a(FE_RN_57));
   in01f06 FE_OCPC2606_n19306 (.o(FE_OCPN25907_n19306),
	.a(FE_RN_57));
   in01f06 FE_OCPC2605_n19306 (.o(FE_OFN24735_n19306),
	.a(FE_RN_57));
   in01f40 FE_OCPC2604_n19306 (.o(FE_OFN24736_n19306),
	.a(n19306));
   in01f01 FE_OCPC2600_n19503 (.o(FE_OFN25690_n19503),
	.a(n19503));
   in01f01 FE_OCPC2599_n19503 (.o(FE_OFN24798_n19503),
	.a(n19503));
   in01f01 FE_OCPC2598_n19503 (.o(n21746),
	.a(n19503));
   in01f01 FE_OCPC2597_n19503 (.o(n19656),
	.a(n19503));
   in01f04 FE_OCPC2595_n18828 (.o(FE_OCPN25929_n18828),
	.a(FE_RN_31));
   in01f01 FE_OCPC2593_n18828 (.o(FE_OCPN25927_n18828),
	.a(n18828));
   in01f04 FE_OCPC2592_n18828 (.o(FE_OCPN25926_n18828),
	.a(n18828));
   in01f08 FE_OCPC2591_n18828 (.o(FE_OCPN25925_n18828),
	.a(n18828));
   in01f02 FE_OCPC2590_n18828 (.o(FE_OFN183_n24390),
	.a(n18828));
   in01f06 FE_OCPC2589_n18828 (.o(n18997),
	.a(n18828));
   in01f10 FE_OCPC2588_n18828 (.o(FE_RN_7),
	.a(n18828));
   in01f01 FE_OCPC2587_n18828 (.o(FE_OFN24748_n18828),
	.a(n18828));
   in01f06 FE_OCPC2586_n18828 (.o(n24390),
	.a(n18828));
   in01f20 FE_OCPC2413_n19499_dup (.o(FE_RN_29),
	.a(n19499));
   in01f08 FE_OFC1716_n25140_dup (.o(FE_RN_28),
	.a(n25140));
   in01f06 FE_OCPC2548_n18828_dup1 (.o(FE_RN_27),
	.a(FE_OCPN25929_n18828));
   no02f06 U21478_dup (.o(FE_RN_26),
	.a(n18014),
	.b(n24954));
   in01f08 FE_OFC1741_n17934_dup (.o(FE_RN_24),
	.a(n17934));
   no02f06 U18697_dup (.o(FE_RN_23),
	.a(n20413),
	.b(n20412));
   ao12f08 U20103_dup (.o(FE_RN_16),
	.a(n20006),
	.b(n20007),
	.c(n21539));
   in01f20 FE_OCPC2585_n18648 (.o(n24472),
	.a(n24964));
   in01f40 FE_OCPC2584_n18648 (.o(FE_OFN24744_n18648),
	.a(n24964));
   in01f40 FE_OCPC2583_n18648 (.o(n24964),
	.a(n18648));
   in01f20 FE_OCPC2582_n18648 (.o(FE_OFN24745_n18648),
	.a(n18648));
   in01f06 FE_OCPC2581_n19547 (.o(FE_OCPN25924_n19547),
	.a(n19547));
   in01f01 FE_OCPC2580_n19547 (.o(FE_OCPN25923_n19547),
	.a(n19547));
   in01f04 FE_OCPC2579_n19547 (.o(FE_OCPN25922_n19547),
	.a(n19547));
   in01f02 FE_OCPC2578_n19547 (.o(FE_OCPN25921_n19547),
	.a(n19547));
   in01f02 FE_OCPC2577_n19547 (.o(FE_OCPN25920_n19547),
	.a(n19547));
   in01f04 FE_OCPC2576_n19547 (.o(FE_OCPN25919_n19547),
	.a(n19547));
   in01f03 FE_OCPC2575_n19547 (.o(FE_OCPN25918_n19547),
	.a(n19547));
   in01f02 FE_OCPC2574_n19547 (.o(FE_OCPN25917_n19547),
	.a(n19547));
   in01f01 FE_OCPC2573_n19547 (.o(FE_OCPN25916_n19547),
	.a(n19547));
   in01f01 FE_OCPC2572_n19547 (.o(FE_OCPN25915_n19547),
	.a(n19547));
   in01f02 FE_OCPC2571_n19547 (.o(FE_OCPN25914_n19547),
	.a(n19547));
   in01f02 FE_OCPC2570_n19547 (.o(FE_OCPN25913_n19547),
	.a(n19547));
   in01f02 FE_OCPC2569_n19547 (.o(FE_OCPN25912_n19547),
	.a(n19547));
   in01f01 FE_OCPC2568_n19547 (.o(FE_OCPN25911_n19547),
	.a(n19547));
   in01f02 FE_OCPC2567_n19547 (.o(FE_OCPN25910_n19547),
	.a(n19547));
   in01f10 FE_OCPC2566_n19547 (.o(FE_OCPN25909_n19547),
	.a(n19547));
   in01f01 FE_OCPC2565_n19547 (.o(FE_OCPN25908_n19547),
	.a(n19547));
   in01f02 FE_OCPC2564_n19547 (.o(n24455),
	.a(n19547));
   in01f02 FE_OCPC2563_n19547 (.o(n18033),
	.a(n19547));
   in01f02 FE_OCPC2562_n19547 (.o(FE_OFN25674_n18033),
	.a(n19547));
   in01f10 FE_OCPC2561_FE_RN_6 (.o(FE_OCPN25816_n20147),
	.a(FE_RN_6));
   no02f10 U23952_dup (.o(FE_RN_22),
	.a(n19044),
	.b(n18734));
   no02f08 U21544_dup (.o(FE_RN_21),
	.a(n19540),
	.b(n19539));
   na04f20 U23393_dup (.o(FE_RN_20),
	.a(n19407),
	.b(n19406),
	.c(n19405),
	.d(n19404));
   in01f08 FE_OFC1896_n21748_dup (.o(FE_RN_19),
	.a(n21748));
   na02f40 U23383_dup (.o(FE_RN_18),
	.a(FE_OFN24792_n17934),
	.b(FE_RN_52));
   in01f40 U23417_dup (.o(FE_RN_17),
	.a(n18754));
   na02f40 U23447_dup (.o(FE_RN_15),
	.a(n17785),
	.b(FE_OCPN25932_n19501));
   na02f20 U24213_dup (.o(FE_RN_14),
	.a(n19345),
	.b(n19344));
   oa12f02 U21828_dup (.o(FE_RN_12),
	.a(n18205),
	.b(n18206),
	.c(n18202));
   no02f20 U24067_dup (.o(FE_RN_11),
	.a(north_input_NIB_head_ptr_f_0_),
	.b(FE_OFN25617_north_input_NIB_head_ptr_f_1));
   no02f20 U24156_dup (.o(FE_RN_9),
	.a(n19244),
	.b(n20297));
   in01f08 U21373_dup (.o(FE_RN_2),
	.a(n17867));
   in01f06 FE_OCPC2558_n19306 (.o(FE_OCPN25905_n19306),
	.a(FE_RN_57));
   oa22f10 FE_RC_39_0 (.o(n19669),
	.a(FE_RN_36),
	.b(n19666),
	.c(n18146),
	.d(myChipID_f_0_));
   no02f40 U23965_dup1 (.o(FE_RN_8),
	.a(n18827),
	.b(FE_OCPN25899_west_input_NIB_head_ptr_f_0));
   no03f40 U23394_dup (.o(FE_RN_6),
	.a(n19410),
	.b(n19409),
	.c(n19408));
   ao22f20 FE_RC_38_0 (.o(n19402),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__58_),
	.c(FE_OCPN25813_FE_OFN24735_n19306),
	.d(east_input_NIB_storage_data_f_1__58_));
   no02f40 U23965_dup (.o(FE_RN_5),
	.a(n18827),
	.b(FE_OCPN25899_west_input_NIB_head_ptr_f_0));
   in01f01 FE_RC_36_0 (.o(FE_RN_22_0),
	.a(n25463));
   no02f01 FE_RC_35_0 (.o(FE_RN_23_0),
	.a(FE_RN_22_0),
	.b(n19496));
   na02f02 FE_RC_34_0 (.o(n25150),
	.a(n25149),
	.b(FE_RN_23_0));
   no04f40 U21564_dup (.o(FE_RN_4),
	.a(FE_RN_46),
	.b(n18699),
	.c(n18700),
	.d(n18698));
   in01f08 FE_OCPC2551_n18927 (.o(FE_OCPN25904_n18927),
	.a(n18927));
   in01f01 FE_OCPC2550_n18927 (.o(n22890),
	.a(FE_RN_65));
   in01f08 U23593_dup (.o(FE_RN_3),
	.a(n18614));
   no02f08 U18583_dup (.o(FE_RN_1),
	.a(FE_OFN25600_reset),
	.b(n18575));
   in01f10 FE_OCPC2549_n23508 (.o(n18913),
	.a(n23508));
   ao22f20 FE_RC_33_0 (.o(n20746),
	.a(FE_RN_64),
	.b(west_input_NIB_storage_data_f_3__60_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__60_));
   in01f02 FE_RC_32_0 (.o(FE_RN_18_0),
	.a(FE_OFN25651_n25499));
   in01f04 FE_RC_31_0 (.o(FE_RN_19_0),
	.a(n24968));
   na02f08 FE_RC_30_0 (.o(FE_RN_20_0),
	.a(FE_RN_19_0),
	.b(FE_RN_18_0));
   no03f08 FE_RC_29_0 (.o(n24972),
	.a(FE_RN_20_0),
	.b(n24971),
	.c(n24970));
   in01f01 FE_OCPC2544_west_input_NIB_head_ptr_f_0 (.o(FE_OCPN25903_west_input_NIB_head_ptr_f_0),
	.a(FE_OFN24761_west_input_NIB_head_ptr_f_0));
   in01f40 FE_OCPC2543_west_input_NIB_head_ptr_f_0 (.o(FE_OCPN25902_west_input_NIB_head_ptr_f_0),
	.a(FE_OFN24761_west_input_NIB_head_ptr_f_0));
   in01f01 FE_OCPC2542_west_input_NIB_head_ptr_f_0 (.o(FE_OCPN25901_west_input_NIB_head_ptr_f_0),
	.a(west_input_NIB_head_ptr_f_0_));
   in01f20 FE_OCPC2541_west_input_NIB_head_ptr_f_0 (.o(FE_OCPN25900_west_input_NIB_head_ptr_f_0),
	.a(west_input_NIB_head_ptr_f_0_));
   in01f20 FE_OCPC2540_west_input_NIB_head_ptr_f_0 (.o(FE_OCPN25899_west_input_NIB_head_ptr_f_0),
	.a(west_input_NIB_head_ptr_f_0_));
   in01f20 FE_OCPC2539_west_input_NIB_head_ptr_f_0 (.o(FE_OFN24761_west_input_NIB_head_ptr_f_0),
	.a(west_input_NIB_head_ptr_f_0_));
   in01f04 FE_OFC2535_n25395 (.o(FE_OFN25895_n25395),
	.a(FE_OFN25889_n25395));
   in01f02 FE_OFC2532_n25395 (.o(FE_OFN25892_n25395),
	.a(FE_OFN25889_n25395));
   in01f10 FE_OFC2531_n25395 (.o(FE_OFN25891_n25395),
	.a(FE_OFN25888_n25395));
   in01f01 FE_OFC2529_n25395 (.o(FE_OFN25889_n25395),
	.a(n25395));
   in01f04 FE_OFC2528_n25395 (.o(FE_OFN25888_n25395),
	.a(n25395));
   in01f01 FE_OFC2527_dataOut_S_48 (.o(dataOut_S_48_),
	.a(FE_OFN25887_dataOut_S_48));
   in01f01 FE_OFC2526_dataOut_S_48 (.o(FE_OFN25887_dataOut_S_48),
	.a(FE_OFN25886_dataOut_S_48));
   in01f01 FE_OFC2525_dataOut_N_48 (.o(dataOut_N_48_),
	.a(FE_OFN25885_dataOut_N_48));
   in01f01 FE_OFC2524_dataOut_N_48 (.o(FE_OFN25885_dataOut_N_48),
	.a(FE_OFN25884_dataOut_N_48));
   in01f01 FE_OFC2523_n19446 (.o(FE_OFN25883_n19446),
	.a(FE_OFN25882_n19446));
   in01f01 FE_OFC2522_n19446 (.o(FE_OFN25882_n19446),
	.a(FE_OFN25878_n19446));
   in01f01 FE_OFC2521_n19446 (.o(FE_OFN25881_n19446),
	.a(FE_OFN25877_n19446));
   in01f10 FE_OFC2520_n19446 (.o(FE_OFN25880_n19446),
	.a(FE_OFN25877_n19446));
   in01f01 FE_OFC2519_n19446 (.o(FE_OFN25879_n19446),
	.a(FE_OFN25877_n19446));
   in01f03 FE_OFC2518_n19446 (.o(FE_OFN25878_n19446),
	.a(FE_OFN25877_n19446));
   in01f08 FE_OFC2517_n19446 (.o(FE_OFN25877_n19446),
	.a(n19446));
   in01f10 FE_OFC2516_n25842 (.o(FE_OFN25876_n25842),
	.a(FE_OFN25874_n25842));
   in01f01 FE_OFC2515_n25842 (.o(FE_OFN25875_n25842),
	.a(FE_OFN25874_n25842));
   in01f03 FE_OFC2514_n25842 (.o(FE_OFN25874_n25842),
	.a(n25842));
   in01f01 FE_OFC2512_FE_OFN42_n19022 (.o(FE_OFN25872_FE_OFN42_n19022),
	.a(FE_OFN25871_FE_OFN42_n19022));
   in01f01 FE_OFC2511_FE_OFN42_n19022 (.o(FE_OFN25871_FE_OFN42_n19022),
	.a(FE_OFN42_n19022));
   in01f01 FE_OFC2509_n21666 (.o(FE_OFN25869_n21666),
	.a(FE_OFN25868_n21666));
   in01f01 FE_OFC2508_n21666 (.o(FE_OFN25868_n21666),
	.a(FE_OFN25976_n21666));
   in01f08 FE_OFC2506_FE_OFN24766_n21069 (.o(FE_OFN25866_FE_OFN24766_n21069),
	.a(FE_OFN25861_FE_OFN24766_n21069));
   in01f01 FE_OFC2505_FE_OFN24766_n21069 (.o(FE_OFN25865_FE_OFN24766_n21069),
	.a(FE_OFN25861_FE_OFN24766_n21069));
   in01f01 FE_OFC2502_FE_OFN24766_n21069 (.o(FE_OFN25862_FE_OFN24766_n21069),
	.a(FE_OFN25860_FE_OFN24766_n21069));
   in01f02 FE_OFC2501_FE_OFN24766_n21069 (.o(FE_OFN25861_FE_OFN24766_n21069),
	.a(FE_OFN24766_n21069));
   in01f01 FE_OFC2500_FE_OFN24766_n21069 (.o(FE_OFN25860_FE_OFN24766_n21069),
	.a(FE_OFN24766_n21069));
   in01f02 FE_OFC2497_FE_OFN899_n17770 (.o(FE_OFN25857_FE_OFN899_n17770),
	.a(FE_OFN25847_FE_OFN899_n17770));
   in01f01 FE_OFC2495_FE_OFN899_n17770 (.o(FE_OFN25855_FE_OFN899_n17770),
	.a(FE_OFN25846_FE_OFN899_n17770));
   in01f01 FE_OFC2494_FE_OFN899_n17770 (.o(FE_OFN25854_FE_OFN899_n17770),
	.a(FE_OFN25846_FE_OFN899_n17770));
   in01f01 FE_OFC2493_FE_OFN899_n17770 (.o(FE_OFN25853_FE_OFN899_n17770),
	.a(FE_OFN25846_FE_OFN899_n17770));
   in01f01 FE_OFC2490_FE_OFN899_n17770 (.o(FE_OFN25850_FE_OFN899_n17770),
	.a(FE_OFN25846_FE_OFN899_n17770));
   in01f01 FE_OFC2489_FE_OFN899_n17770 (.o(FE_OFN25849_FE_OFN899_n17770),
	.a(FE_OFN25846_FE_OFN899_n17770));
   in01f01 FE_OFC2487_FE_OFN899_n17770 (.o(FE_OFN25847_FE_OFN899_n17770),
	.a(FE_OFN899_n17770));
   in01f04 FE_OFC2486_FE_OFN899_n17770 (.o(FE_OFN25846_FE_OFN899_n17770),
	.a(FE_OFN899_n17770));
   in01f01 FE_OFC2485_n20699 (.o(FE_OFN25845_n20699),
	.a(n20700));
   in01f01 FE_OFC2483_n25972 (.o(FE_OFN25843_n25972),
	.a(FE_OFN958_n25972));
   in01f20 FE_OCPC2481_FE_OFN97_n21865 (.o(n19220),
	.a(FE_OFN97_n21865));
   in01f02 FE_RC_28_0 (.o(FE_RN_15_0),
	.a(n20096));
   in01f02 FE_RC_27_0 (.o(FE_RN_16_0),
	.a(n20095));
   no02f06 FE_RC_26_0 (.o(FE_RN_17_0),
	.a(FE_RN_16_0),
	.b(FE_RN_15_0));
   in01f02 FE_RC_24_0 (.o(FE_RN_12_0),
	.a(n20084));
   in01f02 FE_RC_23_0 (.o(FE_RN_13_0),
	.a(n20083));
   no02f04 FE_RC_22_0 (.o(FE_RN_14_0),
	.a(FE_RN_13_0),
	.b(FE_RN_12_0));
   na03f06 FE_RC_21_0 (.o(n20092),
	.a(n20085),
	.b(FE_RN_14_0),
	.c(n20086));
   in01f01 FE_RC_20_0 (.o(FE_RN_9_0),
	.a(n25250));
   in01f01 FE_RC_19_0 (.o(FE_RN_10_0),
	.a(n25249));
   na02f01 FE_RC_18_0 (.o(FE_RN_11_0),
	.a(FE_RN_10_0),
	.b(FE_RN_9_0));
   na02f02 FE_RC_17_0 (.o(n25462),
	.a(n25248),
	.b(FE_RN_11_0));
   in01f01 FE_OCPC2479_n24342 (.o(FE_OCPN25840_n24342),
	.a(FE_OCPN25934_n24342));
   in01f03 FE_OCPC2476_n24342 (.o(FE_OCPN25837_n24342),
	.a(FE_OCPN25934_n24342));
   in01f01 FE_OCPC2473_n24342 (.o(FE_OFN24731_n18131),
	.a(FE_OCPN25934_n24342));
   in01f01 FE_OCPC2472_n24342 (.o(n21740),
	.a(FE_OCPN25934_n24342));
   in01f02 FE_OCPC2469_n25298 (.o(n25307),
	.a(n25298));
   in01f02 FE_OCPC2468_n18593 (.o(n18592),
	.a(n18593));
   in01f10 FE_OCPC2467_n24342 (.o(FE_OCPN25834_n),
	.a(FE_OCPN25934_n24342));
   in01f02 FE_OCPC2465_n20535 (.o(FE_OCPN25831_n20535),
	.a(n20535));
   in01f02 FE_OCPC2464_n20535 (.o(n25172),
	.a(n20535));
   ao22f08 FE_RC_16_0 (.o(n19659),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__53_),
	.c(FE_OFN20_n17779),
	.d(proc_input_NIB_storage_data_f_7__53_));
   in01f01 FE_RC_15_0 (.o(FE_RN_6_0),
	.a(proc_input_NIB_elements_in_array_f_4_));
   no02f01 FE_RC_13_0 (.o(FE_RN_8_0),
	.a(FE_RN_22_0),
	.b(FE_RN_6_0));
   na02f04 FE_RC_12_0 (.o(n25489),
	.a(n25484),
	.b(FE_RN_8_0));
   in01f01 FE_RC_11_0 (.o(FE_RN_3_0),
	.a(n20259));
   in01f01 FE_RC_10_0 (.o(FE_RN_4_0),
	.a(n20545));
   na02f04 FE_RC_9_0 (.o(FE_RN_5_0),
	.a(FE_RN_4_0),
	.b(FE_RN_3_0));
   no03f06 FE_RC_8_0 (.o(n20317),
	.a(n20313),
	.b(n25389),
	.c(FE_RN_5_0));
   in01f01 FE_OCPC2448_n24342 (.o(FE_OCPN25819_n24342),
	.a(FE_OCPN25934_n24342));
   in01f10 FE_OCPC2447_n21745 (.o(FE_OCPN25829_n21745),
	.a(FE_RN_15));
   in01f01 FE_OCPC2446_n21745 (.o(FE_OCPN25828_n21745),
	.a(FE_RN_15));
   in01f01 FE_OCPC2445_n21745 (.o(FE_OCPN25827_n21745),
	.a(FE_RN_15));
   in01f01 FE_OCPC2444_n21745 (.o(FE_OCPN25826_n21745),
	.a(FE_RN_15));
   in01f01 FE_OCPC2443_n21745 (.o(FE_OCPN25825_n21745),
	.a(FE_RN_15));
   in01f02 FE_OCPC2442_n21745 (.o(FE_OCPN25824_n21745),
	.a(n21745));
   in01f02 FE_OCPC2441_n21745 (.o(FE_OCPN25823_n21745),
	.a(n21745));
   in01f03 FE_OCPC2440_n21745 (.o(FE_OCPN25822_n21745),
	.a(n21745));
   in01f02 FE_OCPC2439_n21745 (.o(FE_OFN186_n24453),
	.a(n21745));
   in01f02 FE_OCPC2438_n21745 (.o(n24453),
	.a(n21745));
   no03f06 FE_RC_7_0 (.o(n20125),
	.a(n19859),
	.b(n19889),
	.c(n24954));
   no03f04 FE_RC_6_0 (.o(n25401),
	.a(n25391),
	.b(n25390),
	.c(n25403));
   in01f06 FE_OCPC2437_n25147 (.o(n18575),
	.a(n25147));
   in01f02 FE_OCPC2436_n19632 (.o(FE_OCPN25821_n19632),
	.a(n19632));
   in01f10 FE_OCPC2435_n19632 (.o(n22873),
	.a(n19632));
   in01f40 FE_OCPC2434_west_input_NIB_head_ptr_f_1 (.o(FE_OCPN25820_west_input_NIB_head_ptr_f_1),
	.a(west_input_NIB_head_ptr_f_1_));
   in01f40 FE_OCPC2433_west_input_NIB_head_ptr_f_1 (.o(n18827),
	.a(west_input_NIB_head_ptr_f_1_));
   in01f20 FE_OCPC2423_FE_OFN186_n24453 (.o(FE_OCPN25814_FE_OFN186_n24453),
	.a(FE_RN_15));
   in01f40 FE_OCPC2418_proc_input_NIB_head_ptr_f_1 (.o(n19495),
	.a(proc_input_NIB_head_ptr_f_1_));
   in01f20 FE_OCPC2414_n19499 (.o(FE_OFN24743_n19499),
	.a(FE_RN_29));
   in01f10 FE_OCPC2413_n19499 (.o(n19506),
	.a(n19499));
   in01f10 FE_OCPC2411_n18959 (.o(FE_OCPN25811_n18959),
	.a(FE_OFN25667_n18959));
   in01f06 FE_OCPC2410_n18959 (.o(FE_OCPN25810_n18959),
	.a(n24465));
   in01f02 FE_OCPC2409_n18959 (.o(FE_OCPN25809_n18959),
	.a(FE_RN_5));
   in01f10 FE_OCPC2407_n18959 (.o(FE_OCPN25807_n18959),
	.a(n18959));
   in01f04 FE_OCPC2406_n18959 (.o(FE_OFN25667_n18959),
	.a(n18959));
   in01f20 FE_OCPC2404_n18959 (.o(n24465),
	.a(FE_RN_5));
   ao12f08 FE_RC_5_0 (.o(n20141),
	.a(n18010),
	.b(n25078),
	.c(n20140));
   in01f02 FE_RC_4_0 (.o(FE_RN_0_0),
	.a(n20455));
   in01f02 FE_RC_3_0 (.o(FE_RN_1_0),
	.a(n20454));
   na02f04 FE_RC_2_0 (.o(FE_RN_2_0),
	.a(FE_RN_1_0),
	.b(FE_RN_0_0));
   in01f02 FE_OFC2403_n23051 (.o(FE_OFN25806_n23051),
	.a(FE_OFN25797_n23051));
   in01f02 FE_OFC2399_n23051 (.o(FE_OFN25802_n23051),
	.a(FE_OFN25797_n23051));
   in01f04 FE_OFC2398_n23051 (.o(FE_OFN25801_n23051),
	.a(FE_OFN25796_n23051));
   in01f06 FE_OFC2395_n23051 (.o(FE_OFN25798_n23051),
	.a(FE_OFN25795_n23051));
   in01f02 FE_OFC2394_n23051 (.o(FE_OFN25797_n23051),
	.a(n23051));
   in01f02 FE_OFC2393_n23051 (.o(FE_OFN25796_n23051),
	.a(n23051));
   in01f02 FE_OFC2392_n23051 (.o(FE_OFN25795_n23051),
	.a(n23051));
   in01f01 FE_OFC2391_n21053 (.o(FE_OFN25794_n21053),
	.a(FE_OFN25790_n21053));
   in01f06 FE_OFC2389_n21053 (.o(FE_OFN25792_n21053),
	.a(FE_OFN25789_n21053));
   in01f06 FE_OFC2388_n21053 (.o(FE_OFN25791_n21053),
	.a(FE_OFN25788_n21053));
   in01f01 FE_OFC2387_n21053 (.o(FE_OFN25790_n21053),
	.a(n21053));
   in01f06 FE_OFC2386_n21053 (.o(FE_OFN25789_n21053),
	.a(n21053));
   in01f02 FE_OFC2385_n21053 (.o(FE_OFN25788_n21053),
	.a(n21053));
   in01f02 FE_OFC2384_n17770 (.o(FE_OFN25787_n17770),
	.a(FE_OFN25783_n17770));
   in01f10 FE_OFC2382_n17770 (.o(FE_OFN25785_n17770),
	.a(FE_OFN25783_n17770));
   in01f04 FE_OFC2380_n17770 (.o(FE_OFN25783_n17770),
	.a(n17770));
   in01f10 FE_OFC2379_FE_OFN448_n23236 (.o(FE_OFN25782_FE_OFN448_n23236),
	.a(FE_OFN25780_FE_OFN448_n23236));
   in01f06 FE_OFC2378_FE_OFN448_n23236 (.o(FE_OFN25781_FE_OFN448_n23236),
	.a(FE_OFN25779_FE_OFN448_n23236));
   in01f10 FE_OFC2377_FE_OFN448_n23236 (.o(FE_OFN25780_FE_OFN448_n23236),
	.a(FE_OFN448_n23236));
   in01f01 FE_OFC2376_FE_OFN448_n23236 (.o(FE_OFN25779_FE_OFN448_n23236),
	.a(FE_OFN448_n23236));
   in01f03 FE_OFC2375_FE_OFN582_n25619 (.o(FE_OFN25778_FE_OFN582_n25619),
	.a(FE_OFN25772_FE_OFN582_n25619));
   in01f10 FE_OFC2374_FE_OFN582_n25619 (.o(FE_OFN25777_FE_OFN582_n25619),
	.a(FE_OFN25772_FE_OFN582_n25619));
   in01f01 FE_OFC2373_FE_OFN582_n25619 (.o(FE_OFN25776_FE_OFN582_n25619),
	.a(FE_OFN25771_FE_OFN582_n25619));
   in01f04 FE_OFC2372_FE_OFN582_n25619 (.o(FE_OFN25775_FE_OFN582_n25619),
	.a(FE_OFN25770_FE_OFN582_n25619));
   in01f01 FE_OFC2371_FE_OFN582_n25619 (.o(FE_OFN25774_FE_OFN582_n25619),
	.a(FE_OFN25770_FE_OFN582_n25619));
   in01f01 FE_OFC2370_FE_OFN582_n25619 (.o(FE_OFN25773_FE_OFN582_n25619),
	.a(FE_OFN25769_FE_OFN582_n25619));
   in01f06 FE_OFC2369_FE_OFN582_n25619 (.o(FE_OFN25772_FE_OFN582_n25619),
	.a(FE_OFN582_n25619));
   in01f01 FE_OFC2368_FE_OFN582_n25619 (.o(FE_OFN25771_FE_OFN582_n25619),
	.a(FE_OFN582_n25619));
   in01f01 FE_OFC2367_FE_OFN582_n25619 (.o(FE_OFN25770_FE_OFN582_n25619),
	.a(FE_OFN582_n25619));
   in01f01 FE_OFC2366_FE_OFN582_n25619 (.o(FE_OFN25769_FE_OFN582_n25619),
	.a(FE_OFN582_n25619));
   in01f08 FE_OFC2365_FE_OFN1077_n17766 (.o(FE_OFN25768_FE_OFN1077_n17766),
	.a(FE_OFN25759_FE_OFN1077_n17766));
   in01f01 FE_OFC2364_FE_OFN1077_n17766 (.o(FE_OFN25767_FE_OFN1077_n17766),
	.a(FE_OFN25759_FE_OFN1077_n17766));
   in01f01 FE_OFC2363_FE_OFN1077_n17766 (.o(FE_OFN25766_FE_OFN1077_n17766),
	.a(FE_OFN25758_FE_OFN1077_n17766));
   in01f01 FE_OFC2362_FE_OFN1077_n17766 (.o(FE_OFN25765_FE_OFN1077_n17766),
	.a(FE_OFN25757_FE_OFN1077_n17766));
   in01f06 FE_OFC2360_FE_OFN1077_n17766 (.o(FE_OFN25763_FE_OFN1077_n17766),
	.a(FE_OFN25756_FE_OFN1077_n17766));
   in01f01 FE_OFC2359_FE_OFN1077_n17766 (.o(FE_OFN25762_FE_OFN1077_n17766),
	.a(FE_OFN25755_FE_OFN1077_n17766));
   in01f01 FE_OFC2358_FE_OFN1077_n17766 (.o(FE_OFN25761_FE_OFN1077_n17766),
	.a(FE_OFN25754_FE_OFN1077_n17766));
   in01f01 FE_OFC2357_FE_OFN1077_n17766 (.o(FE_OFN25760_FE_OFN1077_n17766),
	.a(FE_OFN25754_FE_OFN1077_n17766));
   in01f08 FE_OFC2356_FE_OFN1077_n17766 (.o(FE_OFN25759_FE_OFN1077_n17766),
	.a(FE_OFN1077_n17766));
   in01f01 FE_OFC2355_FE_OFN1077_n17766 (.o(FE_OFN25758_FE_OFN1077_n17766),
	.a(FE_OFN1077_n17766));
   in01f01 FE_OFC2354_FE_OFN1077_n17766 (.o(FE_OFN25757_FE_OFN1077_n17766),
	.a(FE_OFN1077_n17766));
   in01f02 FE_OFC2353_FE_OFN1077_n17766 (.o(FE_OFN25756_FE_OFN1077_n17766),
	.a(FE_OFN1077_n17766));
   in01f01 FE_OFC2352_FE_OFN1077_n17766 (.o(FE_OFN25755_FE_OFN1077_n17766),
	.a(FE_OFN1077_n17766));
   in01f01 FE_OFC2351_FE_OFN1077_n17766 (.o(FE_OFN25754_FE_OFN1077_n17766),
	.a(FE_OFN1077_n17766));
   in01f01 FE_OFC2350_FE_OFN24796_n20854 (.o(FE_OFN25753_FE_OFN24796_n20854),
	.a(FE_OFN25745_FE_OFN24796_n20854));
   in01f01 FE_OFC2348_FE_OFN24796_n20854 (.o(FE_OFN25751_FE_OFN24796_n20854),
	.a(FE_OFN25745_FE_OFN24796_n20854));
   in01f03 FE_OFC2347_FE_OFN24796_n20854 (.o(FE_OFN25750_FE_OFN24796_n20854),
	.a(FE_OFN25744_FE_OFN24796_n20854));
   in01f02 FE_OFC2346_FE_OFN24796_n20854 (.o(FE_OFN25749_FE_OFN24796_n20854),
	.a(FE_OFN25744_FE_OFN24796_n20854));
   in01f03 FE_OFC2345_FE_OFN24796_n20854 (.o(FE_OFN25748_FE_OFN24796_n20854),
	.a(FE_OFN25743_FE_OFN24796_n20854));
   in01f03 FE_OFC2344_FE_OFN24796_n20854 (.o(FE_OFN25747_FE_OFN24796_n20854),
	.a(FE_OFN25743_FE_OFN24796_n20854));
   in01f01 FE_OFC2342_FE_OFN24796_n20854 (.o(FE_OFN25745_FE_OFN24796_n20854),
	.a(FE_OFN24796_n20854));
   in01f02 FE_OFC2341_FE_OFN24796_n20854 (.o(FE_OFN25744_FE_OFN24796_n20854),
	.a(FE_OFN24796_n20854));
   in01f02 FE_OFC2340_FE_OFN24796_n20854 (.o(FE_OFN25743_FE_OFN24796_n20854),
	.a(FE_OFN24796_n20854));
   in01f10 FE_OFC2339_FE_OFN25605_n21944 (.o(FE_OFN25742_FE_OFN25605_n21944),
	.a(FE_OFN25738_FE_OFN25605_n21944));
   in01f02 FE_OFC2338_FE_OFN25605_n21944 (.o(FE_OFN25741_FE_OFN25605_n21944),
	.a(FE_OFN25737_FE_OFN25605_n21944));
   in01f01 FE_OFC2337_FE_OFN25605_n21944 (.o(FE_OFN25740_FE_OFN25605_n21944),
	.a(FE_OFN25736_FE_OFN25605_n21944));
   in01f01 FE_OFC2336_FE_OFN25605_n21944 (.o(FE_OFN25739_FE_OFN25605_n21944),
	.a(FE_OFN25735_FE_OFN25605_n21944));
   in01f10 FE_OFC2335_FE_OFN25605_n21944 (.o(FE_OFN25738_FE_OFN25605_n21944),
	.a(FE_OFN25605_n21944));
   in01f01 FE_OFC2334_FE_OFN25605_n21944 (.o(FE_OFN25737_FE_OFN25605_n21944),
	.a(FE_OFN25605_n21944));
   in01f01 FE_OFC2333_FE_OFN25605_n21944 (.o(FE_OFN25736_FE_OFN25605_n21944),
	.a(FE_OFN25605_n21944));
   in01f01 FE_OFC2332_FE_OFN25605_n21944 (.o(FE_OFN25735_FE_OFN25605_n21944),
	.a(FE_OFN25605_n21944));
   in01f02 FE_OFC2331_dataOut_E_8 (.o(dataOut_E_8_),
	.a(FE_OFN25734_dataOut_E_8));
   in01f01 FE_OFC2330_dataOut_E_8 (.o(FE_OFN25734_dataOut_E_8),
	.a(FE_OFN25733_dataOut_E_8));
   in01f02 FE_OFC2329_dataOut_P_9 (.o(dataOut_P_9_),
	.a(FE_OFN25732_dataOut_P_9));
   in01f02 FE_OFC2328_dataOut_P_9 (.o(FE_OFN25732_dataOut_P_9),
	.a(FE_OFN25731_dataOut_P_9));
   in01f02 FE_OFC2327_dataOut_W_9 (.o(dataOut_W_9_),
	.a(FE_OFN25730_dataOut_W_9));
   in01f01 FE_OFC2326_dataOut_W_9 (.o(FE_OFN25730_dataOut_W_9),
	.a(FE_OFN25729_dataOut_W_9));
   in01f02 FE_OFC2325_dataOut_P_31 (.o(dataOut_P_31_),
	.a(FE_OFN25728_dataOut_P_31));
   in01f02 FE_OFC2324_dataOut_P_31 (.o(FE_OFN25728_dataOut_P_31),
	.a(FE_OFN25727_dataOut_P_31));
   in01f02 FE_OFC2323_dataOut_E_37 (.o(dataOut_E_37_),
	.a(FE_OFN25726_dataOut_E_37));
   in01f01 FE_OFC2322_dataOut_E_37 (.o(FE_OFN25726_dataOut_E_37),
	.a(FE_OFN25725_dataOut_E_37));
   in01f02 FE_OFC2321_dataOut_W_31 (.o(dataOut_W_31_),
	.a(FE_OFN25724_dataOut_W_31));
   in01f02 FE_OFC2320_dataOut_W_31 (.o(FE_OFN25724_dataOut_W_31),
	.a(FE_OFN25723_dataOut_W_31));
   in01f02 FE_OFC2319_dataOut_N_31 (.o(dataOut_N_31_),
	.a(FE_OFN25722_dataOut_N_31));
   in01f02 FE_OFC2318_dataOut_N_31 (.o(FE_OFN25722_dataOut_N_31),
	.a(FE_OFN25721_dataOut_N_31));
   in01f02 FE_OFC2317_dataOut_E_22 (.o(dataOut_E_22_),
	.a(FE_OFN25720_dataOut_E_22));
   in01f01 FE_OFC2316_dataOut_E_22 (.o(FE_OFN25720_dataOut_E_22),
	.a(FE_OFN25719_dataOut_E_22));
   in01f01 FE_OFC2315_dataOut_P_37 (.o(dataOut_P_37_),
	.a(FE_OFN25718_dataOut_P_37));
   in01f01 FE_OFC2314_dataOut_P_37 (.o(FE_OFN25718_dataOut_P_37),
	.a(FE_OFN25717_dataOut_P_37));
   in01f01 FE_OFC2313_dataOut_W_37 (.o(dataOut_W_37_),
	.a(FE_OFN25716_dataOut_W_37));
   in01f01 FE_OFC2312_dataOut_W_37 (.o(FE_OFN25716_dataOut_W_37),
	.a(FE_OFN25715_dataOut_W_37));
   in01f01 FE_OFC2311_dataOut_W_48 (.o(dataOut_W_48_),
	.a(FE_OFN25714_dataOut_W_48));
   in01f01 FE_OFC2310_dataOut_W_48 (.o(FE_OFN25714_dataOut_W_48),
	.a(FE_OFN25713_dataOut_W_48));
   in01f01 FE_OFC2309_dataOut_P_49 (.o(dataOut_P_49_),
	.a(FE_OFN25712_dataOut_P_49));
   in01f01 FE_OFC2308_dataOut_P_49 (.o(FE_OFN25712_dataOut_P_49),
	.a(FE_OFN25711_dataOut_P_49));
   in01f01 FE_OFC2307_dataOut_W_49 (.o(dataOut_W_49_),
	.a(FE_OFN25710_dataOut_W_49));
   in01f01 FE_OFC2306_dataOut_W_49 (.o(FE_OFN25710_dataOut_W_49),
	.a(FE_OFN25709_dataOut_W_49));
   in01f01 FE_OFC2305_dataOut_P_35 (.o(dataOut_P_35_),
	.a(FE_OFN25708_dataOut_P_35));
   in01f01 FE_OFC2304_dataOut_P_35 (.o(FE_OFN25708_dataOut_P_35),
	.a(FE_OFN25707_dataOut_P_35));
   in01f01 FE_OFC2303_dataOut_N_35 (.o(dataOut_N_35_),
	.a(FE_OFN25706_dataOut_N_35));
   in01f01 FE_OFC2302_dataOut_N_35 (.o(FE_OFN25706_dataOut_N_35),
	.a(FE_OFN25705_dataOut_N_35));
   in01f01 FE_OFC2301_dataOut_N_37 (.o(dataOut_N_37_),
	.a(FE_OFN25704_dataOut_N_37));
   in01f01 FE_OFC2300_dataOut_N_37 (.o(FE_OFN25704_dataOut_N_37),
	.a(FE_OFN25703_dataOut_N_37));
   in01f02 FE_OFC2299_dataOut_W_35 (.o(dataOut_W_35_),
	.a(FE_OFN25702_dataOut_W_35));
   in01f01 FE_OFC2298_dataOut_W_35 (.o(FE_OFN25702_dataOut_W_35),
	.a(FE_OFN25701_dataOut_W_35));
   in01f01 FE_OFC2297_dataOut_P_48 (.o(dataOut_P_48_),
	.a(FE_OFN25700_dataOut_P_48));
   in01f01 FE_OFC2296_dataOut_P_48 (.o(FE_OFN25700_dataOut_P_48),
	.a(FE_OFN25699_dataOut_P_48));
   in01f02 FE_OFC2295_dataOut_E_39 (.o(dataOut_E_39_),
	.a(FE_OFN25698_dataOut_E_39));
   in01f02 FE_OFC2294_dataOut_E_39 (.o(FE_OFN25698_dataOut_E_39),
	.a(FE_OFN25697_dataOut_E_39));
   in01f20 FE_OFC2293_n18151 (.o(FE_OFN25607_n18151),
	.a(FE_RN_37));
   in01f20 FE_OFC2292_n18151 (.o(n17788),
	.a(n18151));
   in01f01 FE_OFC2291_n19372 (.o(FE_OFN25696_n19372),
	.a(n19372));
   in01f10 FE_OFC2290_n19372 (.o(n24001),
	.a(n19372));
   in01f10 FE_OFC2289_n17814 (.o(FE_OFN25682_n17814),
	.a(n24244));
   in01f20 FE_OFC2288_n17814 (.o(FE_OFN25681_n17814),
	.a(n24244));
   in01f02 FE_OFC2287_n17814 (.o(FE_OFN25680_n17814),
	.a(n24244));
   in01f01 FE_OFC2286_n17814 (.o(FE_OFN25679_n17814),
	.a(n24244));
   in01f01 FE_OFC2285_n17814 (.o(FE_OFN25678_n17814),
	.a(n24244));
   in01f02 FE_OFC2284_n17814 (.o(FE_OFN25677_n17814),
	.a(n24244));
   in01f10 FE_OFC2283_n17814 (.o(n20056),
	.a(n24244));
   in01f08 FE_OFC2282_n17814 (.o(n24060),
	.a(n24244));
   in01f20 FE_OFC2281_n17814 (.o(n19705),
	.a(n24244));
   in01f04 FE_OFC2280_n17814 (.o(n20012),
	.a(n24244));
   in01f20 FE_OFC2279_n17814 (.o(n24244),
	.a(n17814));
   in01f01 FE_OFC2278_n22902 (.o(n25096),
	.a(FE_OFN428_n22902));
   in01f06 FE_OFC2277_n22902 (.o(FE_OFN428_n22902),
	.a(n22902));
   in01f40 FE_OFC2276_proc_input_NIB_head_ptr_f_0 (.o(n20508),
	.a(proc_input_NIB_head_ptr_f_0_));
   in01f01 FE_OFC2273_n19503 (.o(FE_OFN25693_n19503),
	.a(FE_OFN25690_n19503));
   in01f01 FE_OFC2272_n19503 (.o(FE_OFN25692_n19503),
	.a(FE_OFN24798_n19503));
   in01f01 FE_OFC2271_n19503 (.o(FE_OFN25691_n19503),
	.a(n19656));
   in01f01 FE_OFC2269_n19503 (.o(FE_OFN25689_n19503),
	.a(n21746));
   in01f10 FE_OFC2264_n19508 (.o(n17741),
	.a(FE_OFN25606_n19508));
   in01f40 FE_OFC2263_n19508 (.o(n21749),
	.a(FE_OFN25606_n19508));
   in01f10 FE_OFC2262_n19508 (.o(n17744),
	.a(FE_RN_53));
   in01f08 FE_OFC2261_n19508 (.o(n17743),
	.a(FE_RN_53));
   in01f20 FE_OFC2260_n19508 (.o(FE_OFN25606_n19508),
	.a(n19508));
   in01f01 FE_OFC2258_n19500 (.o(FE_OFN25687_n19500),
	.a(FE_OFN25675_n17777));
   in01f01 FE_OFC2256_n19500 (.o(FE_OFN25685_n19500),
	.a(FE_OFN25675_n17777));
   in01f02 FE_OFC2255_n19500 (.o(n17777),
	.a(FE_OFN25675_n17777));
   in01f10 FE_OFC2252_n19547 (.o(FE_OFN25673_n18033),
	.a(n19547));
   in01f01 FE_OFC2248_n21340 (.o(n21341),
	.a(n21340));
   in01f01 FE_OFC2247_n22903 (.o(proc_input_control_N52),
	.a(n22903));
   in01f04 FE_OFC2246_dataOut_P_2 (.o(dataOut_P_2_),
	.a(FE_OFN1073_dataOut_P_2));
   in01f03 FE_OFC2245_dataOut_W_2 (.o(dataOut_W_2_),
	.a(FE_OFN1051_dataOut_W_2));
   in01f02 FE_OFC2244_n24601 (.o(FE_OFN499_n24601),
	.a(FE_OFN498_n24601));
   in01f02 FE_OFC2243_n24630 (.o(FE_OFN211_n24630),
	.a(FE_OFN210_n24630));
   in01f02 FE_OFC2242_dataOut_N_27 (.o(dataOut_N_27_),
	.a(FE_OFN596_dataOut_N_27));
   in01f02 FE_OFC2241_n20239 (.o(n20258),
	.a(n20239));
   in01f02 FE_OFC2240_dataOut_S_26 (.o(dataOut_S_26_),
	.a(FE_OFN702_dataOut_S_26));
   in01f04 FE_OFC2239_dataOut_W_19 (.o(dataOut_W_19_),
	.a(FE_OFN792_dataOut_W_19));
   in01f04 FE_OFC2238_dataOut_N_19 (.o(dataOut_N_19_),
	.a(FE_OFN325_dataOut_N_19));
   in01f04 FE_OFC2237_dataOut_E_6 (.o(dataOut_E_6_),
	.a(FE_OFN656_dataOut_E_6));
   in01f04 FE_OFC2236_east_input_valid (.o(n19456),
	.a(east_input_valid));
   in01f04 FE_OFC2235_dataOut_S_6 (.o(dataOut_S_6_),
	.a(FE_OFN730_dataOut_S_6));
   in01f04 FE_OFC2234_dataOut_P_19 (.o(dataOut_P_19_),
	.a(FE_OFN866_dataOut_P_19));
   in01f04 FE_OFC2233_dataOut_S_17 (.o(dataOut_S_17_),
	.a(FE_OFN718_dataOut_S_17));
   in01f02 FE_OFC2232_dataOut_N_11 (.o(dataOut_N_11_),
	.a(FE_OFN335_dataOut_N_11));
   in01f02 FE_OFC2231_n20292 (.o(n20293),
	.a(n20292));
   in01f03 FE_OFC2230_dataOut_P_17 (.o(dataOut_P_17_),
	.a(FE_OFN868_dataOut_P_17));
   in01f03 FE_OFC2229_dataOut_E_33 (.o(dataOut_E_33_),
	.a(FE_OFN622_dataOut_E_33));
   in01f02 FE_OFC2228_n19884 (.o(n18479),
	.a(n19884));
   in01f03 FE_OFC2227_dataOut_E_19 (.o(dataOut_E_19_),
	.a(FE_OFN642_dataOut_E_19));
   in01f04 FE_OFC2226_dataOut_S_33 (.o(dataOut_S_33_),
	.a(FE_OFN694_dataOut_S_33));
   in01f02 FE_OFC2225_dataOut_S_19 (.o(dataOut_S_19_),
	.a(FE_OFN716_dataOut_S_19));
   in01f02 FE_OFC2224_dataOut_N_10 (.o(dataOut_N_10_),
	.a(FE_OFN337_dataOut_N_10));
   in01f04 FE_OFC2223_dataOut_P_11 (.o(dataOut_P_11_),
	.a(FE_OFN876_dataOut_P_11));
   in01f04 FE_OFC2222_dataOut_W_6 (.o(dataOut_W_6_),
	.a(FE_OFN806_dataOut_W_6));
   in01f02 FE_OFC2221_dataOut_E_11 (.o(dataOut_E_11_),
	.a(FE_OFN652_dataOut_E_11));
   in01f02 FE_OFC2220_n20469 (.o(n18285),
	.a(n20469));
   in01f04 FE_OFC2219_dataOut_N_6 (.o(dataOut_N_6_),
	.a(FE_OFN339_dataOut_N_6));
   in01f03 FE_OFC2218_dataOut_W_11 (.o(dataOut_W_11_),
	.a(FE_OFN802_dataOut_W_11));
   in01f04 FE_OFC2217_dataOut_S_5 (.o(dataOut_S_5_),
	.a(FE_OFN1021_dataOut_S_5));
   in01f04 FE_OFC2216_dataOut_S_11 (.o(dataOut_S_11_),
	.a(FE_OFN726_dataOut_S_11));
   in01f04 FE_OFC2215_dataOut_E_5 (.o(dataOut_E_5_),
	.a(FE_OFN999_dataOut_E_5));
   in01f03 FE_OFC2214_dataOut_N_5 (.o(dataOut_N_5_),
	.a(FE_OFN975_dataOut_N_5));
   in01f03 FE_OFC2213_dataOut_N_17 (.o(dataOut_N_17_),
	.a(FE_OFN327_dataOut_N_17));
   in01f03 FE_OFC2212_dataOut_P_5 (.o(dataOut_P_5_),
	.a(FE_OFN1067_dataOut_P_5));
   in01f02 FE_OFC2211_dataOut_N_2 (.o(dataOut_N_2_),
	.a(FE_OFN981_dataOut_N_2));
   in01f03 FE_OFC2210_dataOut_W_33 (.o(dataOut_W_33_),
	.a(FE_OFN770_dataOut_W_33));
   in01f03 FE_OFC2209_dataOut_P_4 (.o(dataOut_P_4_),
	.a(FE_OFN1069_dataOut_P_4));
   in01f04 FE_OFC2208_dataOut_S_13 (.o(dataOut_S_13_),
	.a(FE_OFN724_dataOut_S_13));
   in01f04 FE_OFC2207_dataOut_W_17 (.o(dataOut_W_17_),
	.a(FE_OFN794_dataOut_W_17));
   in01f01 FE_OFC2206_n24760 (.o(east_output_space_N46),
	.a(n24760));
   in01f03 FE_OFC2205_dataOut_W_5 (.o(dataOut_W_5_),
	.a(FE_OFN1045_dataOut_W_5));
   in01f04 FE_OFC2204_dataOut_S_2 (.o(dataOut_S_2_),
	.a(FE_OFN1027_dataOut_S_2));
   in01f04 FE_OFC2203_dataOut_E_2 (.o(dataOut_E_2_),
	.a(FE_OFN1005_dataOut_E_2));
   in01f20 FE_OFC2199_n19508 (.o(n17742),
	.a(FE_RN_53));
   in01f01 FE_OFC2196_n21435 (.o(n21437),
	.a(n21435));
   in01f04 FE_OFC2195_n25474 (.o(FE_OFN25684_n25474),
	.a(n25474));
   in01f01 FE_OFC2194_n25474 (.o(n25483),
	.a(n25474));
   in01f01 FE_OFC2193_n21333 (.o(n23614),
	.a(n21333));
   in01f02 FE_OFC2192_n20927 (.o(n22844),
	.a(n20927));
   in01f02 FE_OFC2191_n24704 (.o(FE_OFN231_n24704),
	.a(FE_OFN230_n24704));
   in01f08 FE_OFC2184_n20506 (.o(FE_OFN24800_n20506),
	.a(n20506));
   in01f40 FE_OFC2183_n20506 (.o(FE_OFN24799_n20506),
	.a(n20506));
   in01f06 FE_OFC2182_n20506 (.o(n19400),
	.a(n20506));
   in01f02 FE_OFC2169_east_input_NIB_storage_data_f_3__43 (.o(n19260),
	.a(east_input_NIB_storage_data_f_3__43_));
   in01f02 FE_OFC2168_east_input_NIB_storage_data_f_0__26 (.o(n19918),
	.a(east_input_NIB_storage_data_f_0__26_));
   in01f02 FE_OFC2167_proc_input_NIB_storage_data_f_15__25 (.o(n18426),
	.a(proc_input_NIB_storage_data_f_15__25_));
   in01f04 FE_OFC2165_dataOut_E_13 (.o(dataOut_E_13_),
	.a(FE_OFN650_dataOut_E_13));
   in01f02 FE_OFC2164_east_input_NIB_storage_data_f_2__32 (.o(n19302),
	.a(east_input_NIB_storage_data_f_2__32_));
   in01f01 FE_OFC2163_north_input_NIB_storage_data_f_0__22 (.o(n19890),
	.a(north_input_NIB_storage_data_f_0__22_));
   in01f03 FE_OFC2162_dataOut_S_4 (.o(dataOut_S_4_),
	.a(FE_OFN1023_dataOut_S_4));
   in01f02 FE_OFC2161_north_input_NIB_storage_data_f_2__31 (.o(n19104),
	.a(north_input_NIB_storage_data_f_2__31_));
   in01f02 FE_OFC2160_east_input_NIB_storage_data_f_3__26 (.o(n19917),
	.a(east_input_NIB_storage_data_f_3__26_));
   in01f02 FE_OFC2159_south_input_NIB_storage_data_f_2__29 (.o(n18603),
	.a(south_input_NIB_storage_data_f_2__29_));
   in01f01 FE_OFC2158_n20753 (.o(n20756),
	.a(n20753));
   in01f02 FE_OFC2157_n19139 (.o(n19142),
	.a(n19139));
   in01f02 FE_OFC2156_east_input_NIB_storage_data_f_2__34 (.o(n19309),
	.a(east_input_NIB_storage_data_f_2__34_));
   in01f01 FE_OFC2155_north_input_NIB_storage_data_f_3__22 (.o(n19891),
	.a(north_input_NIB_storage_data_f_3__22_));
   in01f03 FE_OFC2154_n18133 (.o(n18132),
	.a(n18133));
   in01f01 FE_OFC2153_n20791 (.o(n20792),
	.a(n20791));
   in01f02 FE_OFC2152_n24978 (.o(n18013),
	.a(n24978));
   in01f01 FE_OFC2151_dataOut_S_15 (.o(dataOut_S_15_),
	.a(FE_OFN722_dataOut_S_15));
   in01f02 FE_OFC2150_dataOut_N_42 (.o(dataOut_N_42_),
	.a(FE_OFN291_dataOut_N_42));
   in01f02 FE_OFC2149_proc_input_NIB_storage_data_f_3__28 (.o(n17911),
	.a(proc_input_NIB_storage_data_f_3__28_));
   in01f02 FE_OFC2148_n18141 (.o(n18140),
	.a(n18141));
   in01f02 FE_OFC2147_proc_input_NIB_storage_data_f_3__23 (.o(n17909),
	.a(proc_input_NIB_storage_data_f_3__23_));
   in01f02 FE_OFC2146_dataOut_W_42 (.o(dataOut_W_42_),
	.a(FE_OFN756_dataOut_W_42));
   in01f02 FE_OFC2145_dataOut_P_36 (.o(dataOut_P_36_),
	.a(FE_OFN838_dataOut_P_36));
   in01f02 FE_OFC2144_dataOut_S_42 (.o(dataOut_S_42_),
	.a(FE_OFN680_dataOut_S_42));
   in01f02 FE_OFC2143_proc_input_NIB_storage_data_f_4__53 (.o(n17739),
	.a(proc_input_NIB_storage_data_f_4__53_));
   in01f02 FE_OFC2142_dataOut_S_36 (.o(dataOut_S_36_),
	.a(FE_OFN688_dataOut_S_36));
   in01f02 FE_OFC2141_dataOut_N_15 (.o(dataOut_N_15_),
	.a(FE_OFN331_dataOut_N_15));
   in01f02 FE_OFC2140_dataOut_E_36 (.o(dataOut_E_36_),
	.a(FE_OFN616_dataOut_E_36));
   in01f03 FE_OFC2139_n23559 (.o(FE_OFN130_n23559),
	.a(FE_OFN129_n23559));
   in01f01 FE_OFC2138_n22519 (.o(n22520),
	.a(n22519));
   in01f01 FE_OFC2137_n22533 (.o(n22534),
	.a(n22533));
   in01f01 FE_OFC2136_n20748 (.o(n20749),
	.a(n20748));
   in01f04 FE_OFC2135_n24579 (.o(FE_OFN495_n24579),
	.a(FE_OFN494_n24579));
   in01f01 FE_OFC2134_n20422 (.o(FE_OFN25676_n20422),
	.a(n20377));
   in01m08 FE_OFC2133_n20422 (.o(n20377),
	.a(n20422));
   in01f20 FE_OFC2132_n19530 (.o(FE_OFN25602_n19530),
	.a(FE_RN_18));
   in01f10 FE_OFC2130_n19530 (.o(FE_OFN191_n24454),
	.a(FE_RN_18));
   in01f10 FE_OFC2129_n19530 (.o(FE_OFN25604_n19530),
	.a(FE_RN_18));
   in01f04 FE_OFC2125_n23576 (.o(FE_OFN923_n23576),
	.a(FE_OFN922_n23576));
   in01f10 FE_OFC2121_myChipID_f_4 (.o(FE_OFN53_n19355),
	.a(myChipID_f_4_));
   in01f10 FE_OFC2120_n19655 (.o(n19709),
	.a(n19688));
   in01f20 FE_OFC2119_n19655 (.o(n21768),
	.a(FE_OFN24806_n19655));
   in01f10 FE_OFC2118_n19655 (.o(n17754),
	.a(FE_OFN25671_n19655));
   in01f08 FE_OFC2117_n19655 (.o(n19707),
	.a(FE_OFN25671_n19655));
   in01f06 FE_OFC2116_n19655 (.o(n19688),
	.a(n19655));
   in01f20 FE_OFC2115_n19655 (.o(FE_OFN24806_n19655),
	.a(n19655));
   in01f10 FE_OFC2114_n19655 (.o(FE_OFN25671_n19655),
	.a(n19655));
   in01f02 FE_OFC2108_dataOut_P_42 (.o(dataOut_P_42_),
	.a(FE_OFN830_dataOut_P_42));
   in01f02 FE_OFC2107_dataOut_N_36 (.o(dataOut_N_36_),
	.a(FE_OFN299_dataOut_N_36));
   in01f02 FE_OFC2106_west_input_NIB_storage_data_f_2__32 (.o(n18952),
	.a(west_input_NIB_storage_data_f_2__32_));
   in01f02 FE_OFC2105_dataOut_W_36 (.o(dataOut_W_36_),
	.a(FE_OFN764_dataOut_W_36));
   in01f02 FE_OFC2104_dataOut_E_42 (.o(dataOut_E_42_),
	.a(FE_OFN608_dataOut_E_42));
   in01f02 FE_OFC2103_dataOut_E_17 (.o(dataOut_E_17_),
	.a(FE_OFN644_dataOut_E_17));
   in01f02 FE_OFC2102_north_input_NIB_storage_data_f_2__41 (.o(n19074),
	.a(north_input_NIB_storage_data_f_2__41_));
   in01f06 FE_OFC2101_n22827 (.o(n19324),
	.a(n22827));
   in01f04 FE_OFC2100_dataOut_N_25 (.o(dataOut_N_25_),
	.a(FE_OFN313_dataOut_N_25));
   in01f01 FE_OFC2099_n23544 (.o(n23545),
	.a(n23544));
   in01f02 FE_OFC2097_dataOut_P_10 (.o(dataOut_P_10_),
	.a(FE_OFN878_dataOut_P_10));
   in01f02 FE_OFC2096_dataOut_E_23 (.o(dataOut_E_23_),
	.a(FE_OFN634_dataOut_E_23));
   in01f02 FE_OFC2095_dataOut_W_10 (.o(dataOut_W_10_),
	.a(FE_OFN804_dataOut_W_10));
   in01f02 FE_OFC2094_n18393 (.o(n18392),
	.a(n18393));
   in01f03 FE_OFC2093_n18096 (.o(n18097),
	.a(n18096));
   in01f02 FE_OFC2092_dataOut_S_23 (.o(dataOut_S_23_),
	.a(FE_OFN708_dataOut_S_23));
   in01f04 FE_OFC2091_dataOut_P_33 (.o(dataOut_P_33_),
	.a(FE_OFN844_dataOut_P_33));
   in01f04 FE_OFC2090_dataOut_N_33 (.o(dataOut_N_33_),
	.a(FE_OFN305_dataOut_N_33));
   in01f03 FE_OFC2089_dataOut_N_4 (.o(dataOut_N_4_),
	.a(FE_OFN977_dataOut_N_4));
   in01f02 FE_OFC2088_dataOut_N_23 (.o(dataOut_N_23_),
	.a(FE_OFN317_dataOut_N_23));
   in01f10 FE_OFC2087_n19421 (.o(n22874),
	.a(n19421));
   in01f02 FE_OFC2086_dataOut_S_43 (.o(dataOut_S_43_),
	.a(FE_OFN678_dataOut_S_43));
   in01f02 FE_OFC2085_dataOut_N_43 (.o(dataOut_N_43_),
	.a(FE_OFN289_dataOut_N_43));
   in01f02 FE_OFC2084_n22773 (.o(FE_OFN25672_n22773),
	.a(FE_OFN111_n22773));
   in01f02 FE_OFC2083_n22773 (.o(FE_OFN525_n24731),
	.a(FE_OFN111_n22773));
   in01f01 FE_OFC2082_n22773 (.o(n24731),
	.a(FE_OFN111_n22773));
   in01f01 FE_OFC2081_n22773 (.o(FE_OFN112_n22773),
	.a(FE_OFN111_n22773));
   in01f08 FE_OFC2080_n22773 (.o(FE_OFN111_n22773),
	.a(n22773));
   in01f03 FE_OFC2079_n24732 (.o(FE_OFN528_n24732),
	.a(FE_OFN527_n24732));
   in01f02 FE_OFC2078_dataOut_E_43 (.o(dataOut_E_43_),
	.a(FE_OFN353_dataOut_E_43));
   in01f02 FE_OFC2077_dataOut_E_4 (.o(dataOut_E_4_),
	.a(FE_OFN1001_dataOut_E_4));
   in01f06 FE_OFC2076_n24739 (.o(FE_OFN239_n24739),
	.a(FE_OFN238_n24739));
   in01f02 FE_OFC2075_dataOut_P_23 (.o(dataOut_P_23_),
	.a(FE_OFN858_dataOut_P_23));
   in01f04 FE_OFC2074_dataOut_P_13 (.o(dataOut_P_13_),
	.a(FE_OFN874_dataOut_P_13));
   in01f02 FE_OFC2073_dataOut_P_43 (.o(dataOut_P_43_),
	.a(FE_OFN828_dataOut_P_43));
   in01f04 FE_OFC2072_n24751 (.o(FE_OFN546_n24751),
	.a(FE_OFN545_n24751));
   in01f03 FE_OFC2071_dataOut_S_20 (.o(dataOut_S_20_),
	.a(FE_OFN714_dataOut_S_20));
   in01f06 FE_OFC2070_n25017 (.o(n25077),
	.a(n25017));
   in01f08 FE_OFC2069_n18963 (.o(n18470),
	.a(n18963));
   in01f08 FE_OFC2068_n19064 (.o(n23036),
	.a(n19064));
   in01f02 FE_OFC2067_dataOut_S_25 (.o(dataOut_S_25_),
	.a(FE_OFN704_dataOut_S_25));
   in01f03 FE_OFC2066_dataOut_S_12 (.o(dataOut_S_12_),
	.a(FE_OFN1013_dataOut_S_12));
   in01f02 FE_OFC2065_east_input_control_header_last_f (.o(n19449),
	.a(east_input_control_header_last_f));
   in01f04 FE_OFC2064_dataOut_N_13 (.o(dataOut_N_13_),
	.a(FE_OFN333_dataOut_N_13));
   in01f01 FE_OFC2063_n20928 (.o(n22846),
	.a(n20928));
   in01f01 FE_OFC2062_n21293 (.o(n22293),
	.a(n21293));
   in01f01 FE_OFC2061_n22766 (.o(FE_OFN424_n22766),
	.a(FE_OFN423_n22766));
   in01f03 FE_OFC2060_dataOut_E_14 (.o(dataOut_E_14_),
	.a(FE_OFN989_dataOut_E_14));
   in01f06 FE_OFC2059_n24719 (.o(FE_OFN233_n24719),
	.a(FE_OFN232_n24719));
   in01f04 FE_OFC2058_n24584 (.o(FE_OFN201_n24584),
	.a(FE_OFN200_n24584));
   in01f06 FE_OFC2057_n21907 (.o(FE_OFN100_n21907),
	.a(FE_OFN99_n21907));
   in01f03 FE_OFC2056_n23148 (.o(FE_OFN116_n23148),
	.a(FE_OFN115_n23148));
   in01f02 FE_OFC2055_dataOut_W_23 (.o(dataOut_W_23_),
	.a(FE_OFN784_dataOut_W_23));
   in01f04 FE_OFC2041_n24027 (.o(FE_OFN153_n24027),
	.a(FE_OFN152_n24027));
   in01f04 FE_OFC2040_n24636 (.o(FE_OFN215_n24636),
	.a(FE_OFN214_n24636));
   in01f10 FE_OFC2039_n23992 (.o(n19354),
	.a(n23992));
   in01f20 FE_OFC2036_n21747 (.o(FE_OFN165_n24129),
	.a(FE_RN_48));
   in01f10 FE_OFC2035_n21747 (.o(FE_OFN156_n24129),
	.a(FE_RN_48));
   in01f20 FE_OFC2032_proc_input_NIB_head_ptr_f_3 (.o(n19496),
	.a(proc_input_NIB_head_ptr_f_3_));
   in01f01 FE_OFC2030_n20137 (.o(n20140),
	.a(n20137));
   in01f10 FE_OFC2027_n19482 (.o(FE_OFN94_n21695),
	.a(n21695));
   in01f06 FE_OFC2026_n19482 (.o(n21695),
	.a(n19482));
   in01f03 FE_OFC2025_n24710 (.o(FE_OFN937_n24710),
	.a(FE_OFN934_n24710));
   in01f03 FE_OFC1999_dataOut_W_4 (.o(dataOut_W_4_),
	.a(FE_OFN1047_dataOut_W_4));
   in01f01 FE_OFC1998_dataOut_S_37 (.o(dataOut_S_37_),
	.a(FE_OFN686_dataOut_S_37));
   in01f03 FE_OFC1997_dataOut_S_10 (.o(dataOut_S_10_),
	.a(FE_OFN728_dataOut_S_10));
   in01f01 FE_OFC1996_dataOut_S_35 (.o(dataOut_S_35_),
	.a(FE_OFN690_dataOut_S_35));
   in01f02 FE_OFC1995_dataOut_N_29 (.o(dataOut_N_29_),
	.a(FE_OFN309_dataOut_N_29));
   in01f02 FE_OFC1994_n18604 (.o(n25071),
	.a(n18604));
   in01f01 FE_OFC1993_dataOut_W_46 (.o(dataOut_W_46_),
	.a(FE_OFN748_dataOut_W_46));
   in01f01 FE_OFC1992_dataOut_S_49 (.o(dataOut_S_49_),
	.a(FE_OFN666_dataOut_S_49));
   in01f02 FE_OFC1991_dataOut_S_1 (.o(dataOut_S_1_),
	.a(FE_OFN732_dataOut_S_1));
   in01f10 FE_OFC1990_myChipID_f_10 (.o(n19387),
	.a(myChipID_f_10_));
   in01f02 FE_OFC1989_dataOut_S_7 (.o(dataOut_S_7_),
	.a(FE_OFN1019_dataOut_S_7));
   in01f03 FE_OFC1988_n24011 (.o(FE_OFN485_n24011),
	.a(FE_OFN484_n24011));
   in01f01 FE_OFC1987_dataOut_S_40 (.o(dataOut_S_40_),
	.a(FE_OFN361_dataOut_S_40));
   in01f01 FE_OFC1986_dataOut_N_40 (.o(dataOut_N_40_),
	.a(FE_OFN1_dataOut_N_40));
   in01f01 FE_OFC1985_dataOut_P_40 (.o(dataOut_P_40_),
	.a(FE_OFN365_dataOut_P_40));
   in01f02 FE_OFC1984_dataOut_S_22 (.o(dataOut_S_22_),
	.a(FE_OFN710_dataOut_S_22));
   in01f02 FE_OFC1983_dataOut_S_31 (.o(dataOut_S_31_),
	.a(FE_OFN1007_dataOut_S_31));
   in01f02 FE_OFC1982_dataOut_S_16 (.o(dataOut_S_16_),
	.a(FE_OFN720_dataOut_S_16));
   in01f01 FE_OFC1981_dataOut_W_40 (.o(dataOut_W_40_),
	.a(FE_OFN363_dataOut_W_40));
   in01f02 FE_OFC1980_dataOut_E_40 (.o(dataOut_E_40_),
	.a(FE_OFN355_dataOut_E_40));
   in01f04 FE_OFC1979_n25499 (.o(FE_OFN25652_n25499),
	.a(n25499));
   in01f02 FE_OFC1978_n25499 (.o(FE_OFN25651_n25499),
	.a(n25499));
   in01f06 FE_OFC1977_n25499 (.o(FE_OFN266_n25499),
	.a(n25499));
   in01f02 FE_OFC1976_dataOut_N_28 (.o(dataOut_N_28_),
	.a(FE_OFN311_dataOut_N_28));
   in01f01 FE_OFC1975_dataOut_S_8 (.o(dataOut_S_8_),
	.a(FE_OFN1017_dataOut_S_8));
   in01f02 FE_OFC1974_dataOut_E_24 (.o(dataOut_E_24_),
	.a(FE_OFN632_dataOut_E_24));
   in01f02 FE_OFC1973_dataOut_E_28 (.o(dataOut_E_28_),
	.a(FE_OFN626_dataOut_E_28));
   in01f02 FE_OFC1972_dataOut_P_29 (.o(dataOut_P_29_),
	.a(FE_OFN846_dataOut_P_29));
   in01f02 FE_OFC1971_dataOut_W_38 (.o(dataOut_W_38_),
	.a(FE_OFN760_dataOut_W_38));
   in01f02 FE_OFC1970_dataOut_E_29 (.o(dataOut_E_29_),
	.a(FE_OFN624_dataOut_E_29));
   in01f02 FE_OFC1969_dataOut_P_24 (.o(dataOut_P_24_),
	.a(FE_OFN856_dataOut_P_24));
   in01f02 FE_OFC1968_dataOut_P_28 (.o(dataOut_P_28_),
	.a(FE_OFN848_dataOut_P_28));
   in01f02 FE_OFC1967_dataOut_S_24 (.o(dataOut_S_24_),
	.a(FE_OFN706_dataOut_S_24));
   in01f02 FE_OFC1966_dataOut_P_38 (.o(dataOut_P_38_),
	.a(FE_OFN834_dataOut_P_38));
   in01f02 FE_OFC1965_dataOut_W_24 (.o(dataOut_W_24_),
	.a(FE_OFN782_dataOut_W_24));
   in01f02 FE_OFC1964_dataOut_S_38 (.o(dataOut_S_38_),
	.a(FE_OFN684_dataOut_S_38));
   in01f02 FE_OFC1963_dataOut_W_28 (.o(dataOut_W_28_),
	.a(FE_OFN774_dataOut_W_28));
   in01f06 FE_OFC1962_n24729 (.o(FE_OFN235_n24729),
	.a(FE_OFN234_n24729));
   in01f04 FE_OFC1961_n24645 (.o(FE_OFN219_n24645),
	.a(FE_OFN218_n24645));
   in01f03 FE_OFC1960_n23536 (.o(FE_OFN128_n23536),
	.a(FE_OFN127_n23536));
   in01f02 FE_OFC1957_dataOut_S_28 (.o(dataOut_S_28_),
	.a(FE_OFN698_dataOut_S_28));
   in01f02 FE_OFC1956_dataOut_S_29 (.o(dataOut_S_29_),
	.a(FE_OFN696_dataOut_S_29));
   in01f03 FE_OFC1954_n24036 (.o(FE_OFN155_n24036),
	.a(FE_OFN154_n24036));
   in01f02 FE_OFC1953_dataOut_N_38 (.o(dataOut_N_38_),
	.a(FE_OFN295_dataOut_N_38));
   in01f03 FE_OFC1952_dataOut_N_24 (.o(dataOut_N_24_),
	.a(FE_OFN315_dataOut_N_24));
   in01f02 FE_OFC1951_dataOut_W_39 (.o(dataOut_W_39_),
	.a(FE_OFN758_dataOut_W_39));
   in01f02 FE_OFC1950_dataOut_N_39 (.o(dataOut_N_39_),
	.a(FE_OFN293_dataOut_N_39));
   in01f02 FE_OFC1948_dataOut_S_39 (.o(dataOut_S_39_),
	.a(FE_OFN682_dataOut_S_39));
   in01f02 FE_OFC1947_dataOut_P_39 (.o(dataOut_P_39_),
	.a(FE_OFN832_dataOut_P_39));
   in01f02 FE_OFC1946_dataOut_E_38 (.o(dataOut_E_38_),
	.a(FE_OFN612_dataOut_E_38));
   in01f02 FE_OFC1945_dataOut_W_34 (.o(dataOut_W_34_),
	.a(FE_OFN768_dataOut_W_34));
   in01f02 FE_OFC1944_dataOut_N_34 (.o(dataOut_N_34_),
	.a(FE_OFN303_dataOut_N_34));
   in01f02 FE_OFC1943_dataOut_P_34 (.o(dataOut_P_34_),
	.a(FE_OFN842_dataOut_P_34));
   in01f02 FE_OFC1942_dataOut_S_34 (.o(dataOut_S_34_),
	.a(FE_OFN692_dataOut_S_34));
   in01f02 FE_OFC1935_dataOut_E_34 (.o(dataOut_E_34_),
	.a(FE_OFN620_dataOut_E_34));
   in01f01 FE_OFC1932_n19482 (.o(n17773),
	.a(n21695));
   in01f04 FE_OFC1917_n18762 (.o(FE_OFN25648_n18762),
	.a(n18762));
   in01f01 FE_OFC1916_n18762 (.o(n24142),
	.a(n18762));
   in01f20 FE_OFC1915_n18762 (.o(n21806),
	.a(n18762));
   in01f08 FE_OFC1914_n18762 (.o(n24208),
	.a(n18762));
   in01f01 FE_OFC1913_n18762 (.o(n24321),
	.a(n18762));
   in01f04 FE_OFC1912_n25979 (.o(n25971),
	.a(n25979));
   in01f40 FE_OFC1911_n18960 (.o(FE_OFN24763_n18960),
	.a(n21829));
   in01f10 FE_OFC1910_n18960 (.o(n24466),
	.a(FE_OFN24762_n18960));
   in01f10 FE_OFC1909_n18960 (.o(FE_OFN24764_n18960),
	.a(FE_OFN24762_n18960));
   in01f20 FE_OFC1908_n18960 (.o(n18995),
	.a(n18960));
   in01f20 FE_OFC1907_n18960 (.o(n21829),
	.a(n18960));
   in01f10 FE_OFC1906_n18960 (.o(FE_OFN24762_n18960),
	.a(n18960));
   in01f06 FE_OFC1903_reset (.o(FE_OFN25647_reset),
	.a(FE_OFN25646_reset));
   in01f01 FE_OFC1902_reset (.o(FE_OFN25646_reset),
	.a(reset));
   in01f02 FE_OFC1901_reset (.o(FE_OFN571_n25463),
	.a(reset));
   in01f01 FE_OFC1900_reset (.o(FE_OFN574_n25463),
	.a(reset));
   in01f01 FE_OFC1899_reset (.o(FE_OFN25597_reset),
	.a(reset));
   in01f01 FE_OFC1898_reset (.o(n25463),
	.a(reset));
   in01f06 FE_OFC1897_n21748 (.o(FE_OFN25645_n21748),
	.a(n21748));
   in01f20 FE_OFC1896_n21748 (.o(FE_OFN170_n24343),
	.a(n21748));
   in01f08 FE_OFC1895_n21748 (.o(FE_OFN168_n24343),
	.a(n21748));
   in01f08 FE_OFC1894_n21748 (.o(FE_OFN167_n24343),
	.a(n21748));
   in01f08 FE_OFC1893_n21748 (.o(n24343),
	.a(n21748));
   in01f10 FE_OFC1892_n21748 (.o(FE_OFN169_n24343),
	.a(n21748));
   in01f20 FE_OFC1891_n19073 (.o(FE_OFN96_n21865),
	.a(n24365));
   in01f06 FE_OFC1890_n19073 (.o(FE_OFN24774_n19073),
	.a(n24365));
   in01f10 FE_OFC1889_n19073 (.o(n21865),
	.a(n24365));
   in01f20 FE_OFC1886_n19073 (.o(n24365),
	.a(n19073));
   in01f20 FE_OFC1885_n19073 (.o(FE_OFN24776_n19073),
	.a(FE_RN_11));
   in01f08 FE_OFC1884_n19073 (.o(FE_OFN97_n21865),
	.a(n19073));
   in01f10 FE_OFC1875_n19225 (.o(FE_OFN48_n19193),
	.a(n19225));
   in01f06 FE_OFC1874_n19225 (.o(n25428),
	.a(n19225));
   in01f10 FE_OFC1873_n19225 (.o(n19193),
	.a(n19225));
   in01f08 FE_OFC1872_n19225 (.o(FE_OFN51_n19193),
	.a(n19225));
   in01f01 FE_OFC1870_n23253 (.o(n7838),
	.a(n23253));
   in01f04 FE_OFC1869_n18139 (.o(n24971),
	.a(n18139));
   in01f01 FE_OFC1868_east_output_space_valid_f (.o(n22371),
	.a(east_output_space_valid_f));
   in01f01 FE_OFC1867_proc_input_NIB_storage_data_f_10__47 (.o(n17847),
	.a(proc_input_NIB_storage_data_f_10__47_));
   in01f02 FE_OFC1866_n18058 (.o(n25104),
	.a(n18058));
   in01f01 FE_OFC1865_n20919 (.o(n22830),
	.a(n20919));
   in01f01 FE_OFC1864_n23587 (.o(n21616),
	.a(n23587));
   in01f02 FE_OFC1863_n25062 (.o(FE_OFN25642_n25062),
	.a(n25062));
   in01f02 FE_OFC1862_n25062 (.o(n25392),
	.a(n25062));
   in01f04 FE_OFC1854_n25384 (.o(n25403),
	.a(n25384));
   in01f06 FE_OFC1853_n19230 (.o(FE_OFN25638_n19230),
	.a(n19230));
   in01f01 FE_OFC1852_n19230 (.o(n22845),
	.a(n19230));
   in01f01 FE_OFC1851_n25434 (.o(west_output_space_N46),
	.a(n25434));
   in01f02 FE_OFC1850_n20503 (.o(n19954),
	.a(n20503));
   in01f04 FE_OFC1849_n18552 (.o(n20226),
	.a(n18552));
   in01f02 FE_OFC1831_n18455 (.o(n18454),
	.a(n18455));
   in01f02 FE_OFC1830_n17872 (.o(n18032),
	.a(n17872));
   in01f02 FE_OFC1829_n19796 (.o(n19797),
	.a(n19796));
   in01f02 FE_OFC1828_n25092 (.o(n25093),
	.a(n25092));
   in01f08 FE_OFC1827_n17868 (.o(n25087),
	.a(n17868));
   in01f01 FE_OFC1826_east_output_space_N44 (.o(n22382),
	.a(east_output_space_N44));
   in01f01 FE_OFC1825_proc_output_space_N44 (.o(n22074),
	.a(proc_output_space_N44));
   in01f10 FE_OFC1824_n23540 (.o(n19386),
	.a(n23540));
   in01f01 FE_OFC1822_n19915 (.o(n19921),
	.a(n19915));
   in01f08 FE_OFC1821_n20933 (.o(n20934),
	.a(FE_OFN1092_n20934));
   in01f06 FE_OFC1820_n20933 (.o(n17771),
	.a(FE_OFN1092_n20934));
   in01f06 FE_OFC1819_n20933 (.o(FE_OFN1092_n20934),
	.a(n20933));
   in01f02 FE_OFC1818_n20356 (.o(n19445),
	.a(n20356));
   in01f06 FE_OFC1817_n19056 (.o(FE_OFN563_n25120),
	.a(n19056));
   in01f04 FE_OFC1816_myLocY_f_2 (.o(FE_OFN67_n19548),
	.a(myLocY_f_2_));
   in01f20 FE_OFC1805_south_input_NIB_head_ptr_f_1 (.o(FE_OFN15_south_input_NIB_head_ptr_f_1),
	.a(south_input_NIB_head_ptr_f_1_));
   in01f08 FE_OFC1802_n19505 (.o(n18121),
	.a(n19505));
   in01f10 FE_OFC1800_n18815 (.o(n18127),
	.a(n18837));
   in01f20 FE_OFC1799_n18815 (.o(FE_OFN27_n18974),
	.a(n18837));
   in01f20 FE_OFC1798_n18815 (.o(FE_OFN26_n18974),
	.a(n18974));
   in01f20 FE_OFC1797_n18815 (.o(n19980),
	.a(n18815));
   in01f20 FE_OFC1796_n18815 (.o(n18837),
	.a(n18815));
   in01f10 FE_OFC1795_n18815 (.o(n18974),
	.a(n18815));
   in01f06 FE_OFC1794_n18815 (.o(FE_OFN30_n18974),
	.a(n18815));
   in01f01 FE_OFC1793_n19165 (.o(FE_OFN25630_n19165),
	.a(n19165));
   in01f06 FE_OFC1792_n19165 (.o(n23342),
	.a(n19165));
   in01f02 FE_OFC1791_n21910 (.o(FE_OFN25629_n21910),
	.a(FE_OFN912_n23246));
   in01f06 FE_OFC1790_n21910 (.o(FE_OFN25628_n21910),
	.a(FE_OFN912_n23246));
   in01f03 FE_OFC1789_n21910 (.o(FE_OFN25627_n21910),
	.a(FE_OFN912_n23246));
   in01f02 FE_OFC1788_n21910 (.o(FE_OFN25626_n21910),
	.a(FE_OFN912_n23246));
   in01f03 FE_OFC1787_n21910 (.o(FE_OFN913_n23246),
	.a(FE_OFN912_n23246));
   in01f02 FE_OFC1786_n21910 (.o(FE_OFN914_n23246),
	.a(FE_OFN912_n23246));
   in01f02 FE_OFC1785_n21910 (.o(n21911),
	.a(FE_OFN912_n23246));
   in01f08 FE_OFC1784_n21910 (.o(FE_OFN912_n23246),
	.a(n21910));
   in01f08 FE_OFC1782_n19003 (.o(FE_OFN25624_n19003),
	.a(n19003));
   in01f01 FE_OFC1781_n19003 (.o(n22882),
	.a(n19003));
   in01f08 FE_OFC1776_n23186 (.o(n18730),
	.a(n23186));
   in01f01 FE_OFC1772_n19123 (.o(FE_OFN25623_n19123),
	.a(n19123));
   in01f04 FE_OFC1771_n19123 (.o(n22837),
	.a(n19123));
   in01f02 FE_OFC1770_n23789 (.o(FE_OFN25622_n23789),
	.a(FE_OFN580_n25547));
   in01f03 FE_OFC1769_n23789 (.o(FE_OFN25621_n23789),
	.a(FE_OFN580_n25547));
   in01f02 FE_OFC1768_n23789 (.o(FE_OFN25620_n23789),
	.a(FE_OFN580_n25547));
   in01f02 FE_OFC1767_n23789 (.o(FE_OFN25619_n23789),
	.a(FE_OFN580_n25547));
   in01f03 FE_OFC1766_n23789 (.o(FE_OFN25618_n23789),
	.a(FE_OFN580_n25547));
   in01f04 FE_OFC1765_n23789 (.o(n17765),
	.a(FE_OFN580_n25547));
   in01f03 FE_OFC1764_n23789 (.o(n25547),
	.a(FE_OFN580_n25547));
   in01f08 FE_OFC1763_n23789 (.o(FE_OFN580_n25547),
	.a(n23789));
   in01f01 FE_OFC1762_n25287 (.o(n21218),
	.a(n25287));
   in01f10 FE_OFC1761_north_input_NIB_head_ptr_f_1 (.o(FE_OFN25617_north_input_NIB_head_ptr_f_1),
	.a(north_input_NIB_head_ptr_f_1_));
   in01f01 FE_OFC1760_north_input_NIB_head_ptr_f_1 (.o(n25430),
	.a(north_input_NIB_head_ptr_f_1_));
   in01f20 FE_OFC1759_n19932 (.o(FE_OFN24780_n19932),
	.a(n19924));
   in01f10 FE_OFC1758_n19932 (.o(FE_OFN24779_n19932),
	.a(n19924));
   in01f20 FE_OFC1757_n19932 (.o(FE_OFN24778_n19932),
	.a(n19924));
   in01f10 FE_OFC1756_n19932 (.o(FE_OFN24777_n19932),
	.a(FE_OFN24787_n19932));
   in01f20 FE_OFC1755_n19932 (.o(n19924),
	.a(n19932));
   in01f06 FE_OFC1754_n19932 (.o(n21858),
	.a(n19932));
   in01f08 FE_OFC1753_n19932 (.o(FE_OFN24787_n19932),
	.a(n19932));
   in01f02 FE_OFC1752_n19007 (.o(FE_OFN25616_n19007),
	.a(n19007));
   in01f04 FE_OFC1751_n19007 (.o(FE_OFN25615_n19007),
	.a(n19007));
   in01f01 FE_OFC1750_n19007 (.o(n22828),
	.a(n19007));
   in01f10 FE_OFC1749_n24002 (.o(n18935),
	.a(n24002));
   in01f10 FE_OFC1748_n22866 (.o(n19378),
	.a(n22866));
   in01f02 FE_OFC1747_n19237 (.o(FE_OFN25614_n19237),
	.a(n19237));
   in01f01 FE_OFC1746_n19237 (.o(n23324),
	.a(n19237));
   in01f04 FE_OFC1743_n20334 (.o(n19736),
	.a(n20334));
   in01f01 FE_OFC1742_n17934 (.o(FE_OFN25613_n17934),
	.a(n17934));
   in01f10 FE_OFC1741_n17934 (.o(FE_OFN24792_n17934),
	.a(n17934));
   in01f20 FE_OFC1740_n17934 (.o(n18145),
	.a(n17934));
   in01f20 FE_OFC1739_n17934 (.o(FE_OFN24793_n17934),
	.a(n17934));
   in01f20 FE_OFC1727_n21745 (.o(FE_OFN188_n24453),
	.a(n21745));
   in01f20 FE_OFC1726_n19507 (.o(n18385),
	.a(n19507));
   in01f10 FE_OFC1716_n25140 (.o(n17785),
	.a(n25140));
   in01f10 FE_OFC1708_n23739 (.o(FE_OFN582_n25619),
	.a(n25619));
   in01f02 FE_OFC1707_n23739 (.o(n17763),
	.a(n23739));
   in01f08 FE_OFC1706_n23739 (.o(n25619),
	.a(n23739));
   in01f06 FE_OFC1704_n20437 (.o(n17813),
	.a(n20437));
   in01f08 FE_OFC1703_n22097 (.o(FE_OFN465_n23476),
	.a(n22098));
   in01f08 FE_OFC1702_n22097 (.o(FE_OFN101_n22098),
	.a(n22098));
   in01f06 FE_OFC1701_n22097 (.o(n22098),
	.a(n22097));
   in01f20 FE_OFC1700_n18377 (.o(FE_OFN25609_n18377),
	.a(n18377));
   in01f10 FE_OFC1699_n18377 (.o(n17811),
	.a(n18377));
   in01f10 FE_OFC1688_n21944 (.o(FE_OFN25605_n21944),
	.a(n21945));
   in01f06 FE_OFC1687_n21944 (.o(FE_OFN453_n23262),
	.a(n21945));
   in01f01 FE_OFC1686_n21944 (.o(FE_OFN452_n23262),
	.a(n21945));
   in01f06 FE_OFC1685_n21944 (.o(n21945),
	.a(n21944));
   in01f03 FE_OFC1661_reset (.o(FE_OFN25601_reset),
	.a(FE_OFN25596_reset));
   in01f06 FE_OFC1660_reset (.o(FE_OFN25600_reset),
	.a(FE_OFN25596_reset));
   in01f02 FE_OFC1659_reset (.o(FE_OFN25599_reset),
	.a(reset));
   in01f10 FE_OFC1658_reset (.o(FE_OFN25598_reset),
	.a(reset));
   in01f10 FE_OFC1656_reset (.o(FE_OFN25596_reset),
	.a(reset));
   in01f02 FE_OFC1654_reset (.o(n25433),
	.a(reset));
   in01f02 FE_OFC1653_n20163 (.o(n20164),
	.a(n20163));
   in01f02 FE_OFC1652_south_input_NIB_storage_data_f_2__34 (.o(n18352),
	.a(south_input_NIB_storage_data_f_2__34_));
   in01f01 FE_OFC1651_proc_input_NIB_storage_data_f_10__30 (.o(n17929),
	.a(proc_input_NIB_storage_data_f_10__30_));
   in01f01 FE_OFC1650_n20107 (.o(n20108),
	.a(n20107));
   in01f06 FE_OFC1649_n19020 (.o(FE_OFN565_n25385),
	.a(n19020));
   in01f03 FE_OFC1648_north_input_NIB_storage_data_f_2__40 (.o(n19078),
	.a(north_input_NIB_storage_data_f_2__40_));
   in01f01 FE_OFC1647_n24726 (.o(n24727),
	.a(n24726));
   in01f02 FE_OFC1646_east_input_NIB_storage_data_f_3__53 (.o(n19375),
	.a(east_input_NIB_storage_data_f_3__53_));
   in01f04 FE_OFC1645_n20501 (.o(FE_OFN902_n18421),
	.a(FE_OFN79_n20501));
   in01f01 FE_OFC1644_n20501 (.o(FE_OFN78_n20501),
	.a(FE_OFN79_n20501));
   in01f10 FE_OFC1643_n20501 (.o(FE_OFN79_n20501),
	.a(n20501));
   in01f01 FE_OFC1642_n18646 (.o(n18647),
	.a(n18646));
   in01f10 FE_OFC1641_n19871 (.o(n17774),
	.a(n19871));
   in01f03 FE_OFC1640_north_input_NIB_storage_data_f_1__40 (.o(n19079),
	.a(north_input_NIB_storage_data_f_1__40_));
   in01f03 FE_OFC1639_proc_input_NIB_storage_data_f_10__51 (.o(n17927),
	.a(proc_input_NIB_storage_data_f_10__51_));
   in01f02 FE_OFC1638_proc_input_NIB_storage_data_f_3__53 (.o(n17933),
	.a(proc_input_NIB_storage_data_f_3__53_));
   in01f01 FE_OFC1637_n22604 (.o(n22605),
	.a(n22604));
   in01f02 FE_OFC1636_proc_input_NIB_storage_data_f_3__49 (.o(n17849),
	.a(proc_input_NIB_storage_data_f_3__49_));
   in01f03 FE_OFC1635_proc_input_NIB_storage_data_f_3__51 (.o(n17907),
	.a(proc_input_NIB_storage_data_f_3__51_));
   in01f03 FE_OFC1634_west_input_NIB_storage_data_f_2__54 (.o(n18893),
	.a(west_input_NIB_storage_data_f_2__54_));
   in01f10 FE_OFC1633_myChipID_f_13 (.o(n19617),
	.a(myChipID_f_13_));
   in01f01 FE_OFC1632_n21336 (.o(n21337),
	.a(n21336));
   in01f01 FE_OFC1631_n23054 (.o(n5618),
	.a(n23054));
   in01f01 FE_OFC1630_n23558 (.o(north_output_space_N46),
	.a(n23558));
   in01f01 FE_OFC1629_n25614 (.o(n4343),
	.a(n25614));
   in01f01 FE_OFC1628_n23130 (.o(n4913),
	.a(n23130));
   in01f01 FE_OFC1627_n24482 (.o(n24483),
	.a(n24482));
   in01f01 FE_OFC1626_n21166 (.o(n21167),
	.a(n21166));
   in01f01 FE_OFC1625_n24374 (.o(n24375),
	.a(n24374));
   in01f01 FE_OFC1624_n21132 (.o(n21133),
	.a(n21132));
   in01f01 FE_OFC1623_n22412 (.o(n10778),
	.a(n22412));
   in01f01 FE_OFC1622_n24490 (.o(n24491),
	.a(n24490));
   in01f01 FE_OFC1621_n20963 (.o(n20964),
	.a(n20963));
   in01f04 FE_OFC1620_n22945 (.o(FE_OFN24862_n22945),
	.a(FE_OFN24861_n22945));
   in01f06 FE_OFC1619_n22945 (.o(FE_OFN24861_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1618_n22945 (.o(FE_OFN24860_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1617_n22945 (.o(FE_OFN24859_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1616_n22945 (.o(FE_OFN24858_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1615_n22945 (.o(FE_OFN24857_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1614_n22945 (.o(FE_OFN24856_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1613_n22945 (.o(FE_OFN24855_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1612_n22945 (.o(FE_OFN24854_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1611_n22945 (.o(FE_OFN24853_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1610_n22945 (.o(FE_OFN24852_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1609_n22945 (.o(FE_OFN24851_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1608_n22945 (.o(FE_OFN24850_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1607_n22945 (.o(FE_OFN24849_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1606_n22945 (.o(FE_OFN24848_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1605_n22945 (.o(FE_OFN24847_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1604_n22945 (.o(FE_OFN24846_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1603_n22945 (.o(FE_OFN24845_n22945),
	.a(FE_OFN431_n22945));
   in01m03 FE_OFC1602_n22945 (.o(FE_OFN24844_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1601_n22945 (.o(FE_OFN24843_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1600_n22945 (.o(FE_OFN24842_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1599_n22945 (.o(FE_OFN24841_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1598_n22945 (.o(FE_OFN24840_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1597_n22945 (.o(FE_OFN24839_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1596_n22945 (.o(FE_OFN24838_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1595_n22945 (.o(FE_OFN24837_n22945),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1594_n22945 (.o(n22946),
	.a(FE_OFN431_n22945));
   in01f01 FE_OFC1593_n22945 (.o(FE_OFN433_n22945),
	.a(FE_OFN431_n22945));
   in01f06 FE_OFC1592_n22945 (.o(FE_OFN431_n22945),
	.a(n22945));
   in01f01 FE_OFC1591_n22902 (.o(FE_OFN947_n25096),
	.a(FE_OFN428_n22902));
   in01f01 FE_OFC1589_n22902 (.o(FE_OFN946_n25096),
	.a(FE_OFN428_n22902));
   in01f01 FE_OFC1586_n22517 (.o(FE_OFN24836_n22517),
	.a(FE_OFN105_n22517));
   in01f01 FE_OFC1585_n22517 (.o(FE_OFN24835_n22517),
	.a(FE_OFN105_n22517));
   in01f01 FE_OFC1584_n22517 (.o(FE_OFN24834_n22517),
	.a(FE_OFN105_n22517));
   in01f01 FE_OFC1583_n22517 (.o(FE_OFN386_n17783),
	.a(FE_OFN105_n22517));
   in01f01 FE_OFC1582_n22517 (.o(FE_OFN387_n17783),
	.a(FE_OFN105_n22517));
   in01f01 FE_OFC1581_n22517 (.o(n17783),
	.a(FE_OFN105_n22517));
   in01f01 FE_OFC1580_n22517 (.o(FE_OFN106_n22517),
	.a(FE_OFN105_n22517));
   in01f10 FE_OFC1579_n22517 (.o(FE_OFN105_n22517),
	.a(n22517));
   in01f01 FE_OFC1578_n24438 (.o(n24439),
	.a(n24438));
   in01f01 FE_OFC1577_n24558 (.o(n24559),
	.a(n24558));
   in01f01 FE_OFC1576_n22219 (.o(n22220),
	.a(n22219));
   in01f01 FE_OFC1575_n24673 (.o(n24674),
	.a(n24673));
   in01f01 FE_OFC1574_n21136 (.o(n21137),
	.a(n21136));
   in01f01 FE_OFC1573_n24717 (.o(n24718),
	.a(n24717));
   in01f02 FE_OFC1572_east_input_NIB_storage_data_f_1__38 (.o(n24905),
	.a(east_input_NIB_storage_data_f_1__38_));
   in01f01 FE_OFC1571_n25232 (.o(FE_OFN24833_n25232),
	.a(n24970));
   in01f01 FE_OFC1570_n25232 (.o(FE_OFN24832_n25232),
	.a(n24970));
   in01f02 FE_OFC1569_n25232 (.o(FE_OFN24831_n25232),
	.a(n24970));
   in01f08 FE_OFC1568_n25232 (.o(n24970),
	.a(n25232));
   in01f01 FE_OFC1567_n24617 (.o(n24618),
	.a(n24617));
   in01f01 FE_OFC1566_n21397 (.o(n21398),
	.a(n21397));
   in01f01 FE_OFC1565_n24430 (.o(n24431),
	.a(n24430));
   in01f02 FE_OFC1564_n25499 (.o(FE_OFN24830_n25499),
	.a(FE_OFN266_n25499));
   in01f01 FE_OFC1563_n25499 (.o(FE_OFN24829_n25499),
	.a(FE_OFN266_n25499));
   in01f01 FE_OFC1562_n25499 (.o(FE_OFN24828_n25499),
	.a(FE_OFN266_n25499));
   in01f01 FE_OFC1561_n25499 (.o(FE_OFN24827_n25499),
	.a(FE_OFN266_n25499));
   in01f01 FE_OFC1560_n25499 (.o(FE_OFN24826_n25499),
	.a(FE_OFN266_n25499));
   in01f01 FE_OFC1559_n25499 (.o(FE_OFN24825_n25499),
	.a(FE_OFN266_n25499));
   in01f01 FE_OFC1558_n25499 (.o(FE_OFN559_n24969),
	.a(FE_OFN266_n25499));
   in01f01 FE_OFC1557_n25499 (.o(FE_OFN558_n24969),
	.a(FE_OFN266_n25499));
   in01f01 FE_OFC1556_n25499 (.o(FE_OFN557_n24969),
	.a(FE_OFN266_n25499));
   in01f06 FE_OFC1552_n20737 (.o(n21893),
	.a(n20737));
   in01f01 FE_OFC1551_n24402 (.o(n24403),
	.a(n24402));
   in01f01 FE_OFC1550_n24546 (.o(n24547),
	.a(n24546));
   in01f02 FE_OFC1549_east_input_NIB_storage_data_f_3__60 (.o(n19382),
	.a(east_input_NIB_storage_data_f_3__60_));
   in01f01 FE_OFC1548_n24648 (.o(n24649),
	.a(n24648));
   in01f02 FE_OFC1547_n24977 (.o(n17749),
	.a(n24977));
   in01f01 FE_OFC1546_n24410 (.o(n24411),
	.a(n24410));
   in01f02 FE_OFC1545_n21667 (.o(FE_OFN540_n24743),
	.a(FE_OFN93_n21667));
   in01f01 FE_OFC1544_n21667 (.o(FE_OFN539_n24743),
	.a(FE_OFN93_n21667));
   in01f01 FE_OFC1543_n21667 (.o(FE_OFN538_n24743),
	.a(FE_OFN93_n21667));
   in01f01 FE_OFC1542_n21667 (.o(FE_OFN537_n24743),
	.a(FE_OFN93_n21667));
   in01f01 FE_OFC1541_n21667 (.o(FE_OFN535_n24743),
	.a(FE_OFN93_n21667));
   in01f01 FE_OFC1540_n21667 (.o(FE_OFN534_n24743),
	.a(FE_OFN93_n21667));
   in01f01 FE_OFC1539_n21667 (.o(FE_OFN533_n24743),
	.a(FE_OFN93_n21667));
   in01f01 FE_OFC1538_n21667 (.o(n24743),
	.a(FE_OFN93_n21667));
   in01f01 FE_OFC1537_n21667 (.o(FE_OFN92_n21667),
	.a(FE_OFN93_n21667));
   in01f01 FE_OFC1536_n21667 (.o(FE_OFN536_n24743),
	.a(FE_OFN93_n21667));
   in01f10 FE_OFC1535_n21667 (.o(FE_OFN93_n21667),
	.a(n21667));
   in01f01 FE_OFC1534_n22231 (.o(n22232),
	.a(n22231));
   in01f01 FE_OFC1533_n24530 (.o(n24531),
	.a(n24530));
   in01f10 FE_OFC1532_myChipID_f_8 (.o(n19575),
	.a(myChipID_f_8_));
   in01f01 FE_OFC1531_n24196 (.o(n24197),
	.a(n24196));
   in01f01 FE_OFC1530_n23971 (.o(n23972),
	.a(n23971));
   in01f01 FE_OFC1529_n24265 (.o(n24266),
	.a(n24265));
   in01f01 FE_OFC1528_n24518 (.o(n24519),
	.a(n24518));
   in01f01 FE_OFC1527_n22365 (.o(n22366),
	.a(n22365));
   in01f01 FE_OFC1526_n24570 (.o(n24571),
	.a(n24570));
   in01f01 FE_OFC1525_n24699 (.o(n24700),
	.a(n24699));
   in01f01 FE_OFC1524_n20967 (.o(n20968),
	.a(n20967));
   in01f10 FE_OFC1523_myChipID_f_7 (.o(FE_OFN73_n19631),
	.a(myChipID_f_7_));
   in01f01 FE_OFC1522_n24708 (.o(n24709),
	.a(n24708));
   in01f02 FE_OFC1521_n22357 (.o(n22358),
	.a(n22357));
   in01f06 FE_OFC1520_n19059 (.o(FE_OFN366_n17753),
	.a(n25095));
   in01f02 FE_OFC1519_n19059 (.o(n17753),
	.a(n25095));
   in01f06 FE_OFC1518_n19059 (.o(n25095),
	.a(n19059));
   in01f01 FE_OFC1517_n24418 (.o(n24419),
	.a(n24418));
   in01f01 FE_OFC1516_n24174 (.o(n24175),
	.a(n24174));
   in01f01 FE_OFC1515_n24634 (.o(n24635),
	.a(n24634));
   in01f01 FE_OFC1514_n19916 (.o(n19920),
	.a(n19916));
   in01f01 FE_OFC1513_n22285 (.o(n22286),
	.a(n22285));
   in01f02 FE_OFC1512_n24681 (.o(n24682),
	.a(n24681));
   in01f01 FE_OFC1511_n22353 (.o(n22354),
	.a(n22353));
   in01f01 FE_OFC1510_n24550 (.o(n24551),
	.a(n24550));
   in01f03 FE_OFC1509_n23535 (.o(n17863),
	.a(n23535));
   in01f01 FE_OFC1508_n24498 (.o(n24499),
	.a(n24498));
   in01f01 FE_OFC1507_n24058 (.o(n24059),
	.a(n24058));
   in01f01 FE_OFC1506_n24309 (.o(n24310),
	.a(n24309));
   in01f01 FE_OFC1504_n24690 (.o(n24691),
	.a(n24690));
   in01f01 FE_OFC1503_n21836 (.o(n21837),
	.a(n21836));
   in01f02 FE_OFC1502_n24643 (.o(n24644),
	.a(n24643));
   in01f02 FE_OFC1501_n22616 (.o(n22617),
	.a(n22616));
   in01f01 FE_OFC1500_n24921 (.o(FE_OFN24824_n24921),
	.a(FE_OFN940_n24921));
   in01f01 FE_OFC1499_n24921 (.o(FE_OFN24823_n24921),
	.a(FE_OFN940_n24921));
   in01f01 FE_OFC1498_n24921 (.o(FE_OFN24822_n24921),
	.a(FE_OFN940_n24921));
   in01f01 FE_OFC1497_n24921 (.o(FE_OFN24821_n24921),
	.a(FE_OFN940_n24921));
   in01f01 FE_OFC1496_n24921 (.o(FE_OFN24820_n24921),
	.a(FE_OFN940_n24921));
   in01f01 FE_OFC1495_n24921 (.o(FE_OFN24819_n24921),
	.a(FE_OFN940_n24921));
   in01f01 FE_OFC1494_n24921 (.o(FE_OFN24818_n24921),
	.a(FE_OFN940_n24921));
   in01f01 FE_OFC1493_n24921 (.o(FE_OFN24817_n24921),
	.a(FE_OFN940_n24921));
   in01f01 FE_OFC1492_n24921 (.o(FE_OFN24816_n24921),
	.a(FE_OFN940_n24921));
   in01f01 FE_OFC1491_n24921 (.o(n25869),
	.a(FE_OFN940_n24921));
   in01f01 FE_OFC1490_n24921 (.o(FE_OFN942_n24921),
	.a(FE_OFN940_n24921));
   in01f06 FE_OFC1489_n24921 (.o(FE_OFN940_n24921),
	.a(n24921));
   in01f01 FE_OFC1488_n22600 (.o(n22601),
	.a(n22600));
   in01f01 FE_OFC1487_n24574 (.o(n24575),
	.a(n24574));
   in01f01 FE_OFC1486_n24566 (.o(n24567),
	.a(n24566));
   in01f01 FE_OFC1485_n24625 (.o(n24626),
	.a(n24625));
   in01f01 FE_OFC1484_n21880 (.o(n21881),
	.a(n21880));
   in01f06 FE_OFC1483_myLocY_f_6 (.o(FE_OFN65_n19542),
	.a(myLocY_f_6_));
   in01f02 FE_OFC1482_n19827 (.o(n18445),
	.a(n19827));
   in01f01 FE_OFC1481_n24562 (.o(n24563),
	.a(n24562));
   in01f02 FE_OFC1480_n24757 (.o(n24758),
	.a(n24757));
   in01f01 FE_OFC1479_n24510 (.o(n24511),
	.a(n24510));
   in01f01 FE_OFC1478_n24378 (.o(n24379),
	.a(n24378));
   in01f01 FE_OFC1477_n24406 (.o(n24407),
	.a(n24406));
   in01f01 FE_OFC1476_n24542 (.o(n24543),
	.a(n24542));
   in01f01 FE_OFC1475_n24478 (.o(n24479),
	.a(n24478));
   in01f01 FE_OFC1474_n22958 (.o(FE_OFN24815_n22958),
	.a(FE_OFN435_n22958));
   in01f01 FE_OFC1473_n22958 (.o(FE_OFN24814_n22958),
	.a(FE_OFN435_n22958));
   in01f01 FE_OFC1472_n22958 (.o(FE_OFN24813_n22958),
	.a(FE_OFN435_n22958));
   in01f01 FE_OFC1471_n22958 (.o(FE_OFN24812_n22958),
	.a(FE_OFN435_n22958));
   in01f01 FE_OFC1470_n22958 (.o(FE_OFN24811_n22958),
	.a(FE_OFN435_n22958));
   in01f01 FE_OFC1469_n22958 (.o(FE_OFN24810_n22958),
	.a(FE_OFN435_n22958));
   in01f01 FE_OFC1468_n22958 (.o(FE_OFN24809_n22958),
	.a(FE_OFN435_n22958));
   in01f01 FE_OFC1467_n22958 (.o(FE_OFN24808_n22958),
	.a(FE_OFN435_n22958));
   in01f01 FE_OFC1466_n22958 (.o(FE_OFN24807_n22958),
	.a(FE_OFN435_n22958));
   in01f01 FE_OFC1465_n22958 (.o(FE_OFN438_n22958),
	.a(FE_OFN435_n22958));
   in01f01 FE_OFC1464_n22958 (.o(n22959),
	.a(FE_OFN435_n22958));
   in01f06 FE_OFC1463_n22958 (.o(FE_OFN435_n22958),
	.a(n22958));
   in01f02 FE_OFC1462_n21374 (.o(n21375),
	.a(n21374));
   in01f01 FE_OFC1461_n24652 (.o(n24653),
	.a(n24652));
   in01f01 FE_OFC1460_n21844 (.o(n21845),
	.a(n21844));
   in01f01 FE_OFC1459_n24434 (.o(n24435),
	.a(n24434));
   in01f01 FE_OFC1458_n24609 (.o(n24610),
	.a(n24609));
   in01f01 FE_OFC1447_n24747 (.o(n24748),
	.a(n24747));
   in01f01 FE_OFC1446_n24554 (.o(n24555),
	.a(n24554));
   in01f01 FE_OFC1445_n24526 (.o(n24527),
	.a(n24526));
   in01f02 FE_OFC1444_n25973 (.o(n25980),
	.a(n25973));
   in01f01 FE_OFC1443_n22433 (.o(n22434),
	.a(n22433));
   in01f01 FE_OFC1442_n24016 (.o(n24017),
	.a(n24016));
   in01f01 FE_OFC1441_n21876 (.o(n21877),
	.a(n21876));
   in01f01 FE_OFC1440_n24336 (.o(n24337),
	.a(n24336));
   in01f01 FE_OFC1439_n24582 (.o(n24583),
	.a(n24582));
   in01f01 FE_OFC1429_n24105 (.o(n24106),
	.a(n24105));
   in01f02 FE_OFC1428_n21324 (.o(n21325),
	.a(n21324));
   in01f10 FE_OFC1401_n22139 (.o(FE_OFN103_n22140),
	.a(n22140));
   in01f08 FE_OFC1400_n22139 (.o(n23453),
	.a(n22140));
   in01f06 FE_OFC1399_n22139 (.o(n22140),
	.a(n22139));
   in01f02 FE_OFC1398_n22139 (.o(FE_OFN104_n22140),
	.a(n22139));
   in01f10 FE_OFC1397_n20858 (.o(FE_OFN381_n17772),
	.a(n17772));
   in01m06 FE_OFC1396_n20858 (.o(FE_OFN382_n17772),
	.a(n17772));
   in01f03 FE_OFC1395_n20858 (.o(FE_OFN380_n17772),
	.a(n20858));
   in01f02 FE_OFC1394_n20858 (.o(n17772),
	.a(n20858));
   in01f10 FE_OFC1384_n22084 (.o(n22085),
	.a(FE_OFN416_n22085));
   in01f08 FE_OFC1383_n22084 (.o(n23471),
	.a(FE_OFN416_n22085));
   in01f06 FE_OFC1382_n22084 (.o(FE_OFN416_n22085),
	.a(n22084));
   in01f10 FE_OFC1381_n22778 (.o(FE_OFN1085_n22923),
	.a(n22779));
   in01f06 FE_OFC1380_n22778 (.o(FE_OFN1086_n22923),
	.a(n22779));
   in01f02 FE_OFC1379_n22778 (.o(n22923),
	.a(n22779));
   in01f06 FE_OFC1378_n22778 (.o(n22779),
	.a(n22778));
   in01f01 FE_OFC1377_n25977 (.o(n22271),
	.a(n25977));
   in01f04 FE_OFC1376_n20854 (.o(FE_OFN24796_n20854),
	.a(n20855));
   in01f01 FE_OFC1375_n20854 (.o(FE_OFN24795_n20854),
	.a(n20855));
   in01f01 FE_OFC1374_n20854 (.o(FE_OFN24794_n20854),
	.a(n20855));
   in01f01 FE_OFC1373_n20854 (.o(FE_OFN1102_n25965),
	.a(n20855));
   in01f01 FE_OFC1372_n20854 (.o(FE_OFN1090_n20855),
	.a(n20855));
   in01f01 FE_OFC1371_n20854 (.o(FE_OFN1101_n25965),
	.a(n20855));
   in01f01 FE_OFC1370_n20854 (.o(FE_OFN1089_n20855),
	.a(n20855));
   in01f01 FE_OFC1369_n20854 (.o(n25965),
	.a(n20855));
   in01f01 FE_OFC1368_n20854 (.o(FE_OFN1083_n20854),
	.a(n20855));
   in01m03 FE_OFC1367_n20854 (.o(FE_OFN1084_n20854),
	.a(n20855));
   in01f06 FE_OFC1366_n20854 (.o(n20855),
	.a(n20854));
   in01f03 FE_OFC1365_validIn_P (.o(n25978),
	.a(validIn_P));
   in01f10 FE_OFC1364_n23089 (.o(FE_OFN1077_n17766),
	.a(n23090));
   in01f01 FE_OFC1363_n23089 (.o(FE_OFN1076_n17766),
	.a(n23090));
   in01f01 FE_OFC1362_n23089 (.o(FE_OFN1075_n17766),
	.a(n23090));
   in01f01 FE_OFC1361_n23089 (.o(FE_OFN1074_n17766),
	.a(n23090));
   in01m03 FE_OFC1360_n23089 (.o(n17766),
	.a(n23090));
   in01f08 FE_OFC1359_n23089 (.o(n23090),
	.a(n23089));
   in01f20 FE_OFC1350_east_input_NIB_head_ptr_f_1 (.o(n18442),
	.a(east_input_NIB_head_ptr_f_1_));
   in01f10 FE_OFC1349_n20995 (.o(n17769),
	.a(n20996));
   in01f10 FE_OFC1348_n20995 (.o(FE_OFN896_n17769),
	.a(n20996));
   in01f06 FE_OFC1347_n20995 (.o(n20996),
	.a(n20995));
   in01f06 FE_OFC1346_n23101 (.o(FE_OFN369_n17761),
	.a(n23102));
   in01f10 FE_OFC1345_n23101 (.o(FE_OFN368_n17761),
	.a(n23102));
   in01f01 FE_OFC1344_n23101 (.o(n17761),
	.a(n23102));
   in01f01 FE_OFC1343_n23101 (.o(FE_OFN114_n23102),
	.a(n23102));
   in01f01 FE_OFC1342_n23101 (.o(FE_OFN113_n23102),
	.a(n23102));
   in01f01 FE_OFC1341_n23101 (.o(FE_OFN370_n17761),
	.a(n23102));
   in01f08 FE_OFC1340_n23101 (.o(n23102),
	.a(n23101));
   in01f01 FE_OFC1318_n19932 (.o(n20507),
	.a(FE_OFN24777_n19932));
   in01f20 FE_OFC1305_n19075 (.o(FE_OFN24773_n19075),
	.a(FE_OFN265_n25427));
   in01f03 FE_OFC1304_n19075 (.o(FE_OFN24772_n19075),
	.a(FE_OFN265_n25427));
   in01f08 FE_OFC1303_n19075 (.o(FE_OFN24771_n19075),
	.a(FE_OFN265_n25427));
   in01f10 FE_OFC1302_n19075 (.o(FE_OFN24770_n19075),
	.a(FE_OFN265_n25427));
   in01f10 FE_OFC1301_n19075 (.o(FE_OFN24769_n19075),
	.a(n19192));
   in01f08 FE_OFC1300_n19075 (.o(FE_OFN24768_n19075),
	.a(n19192));
   in01f20 FE_OFC1299_n19075 (.o(FE_OFN265_n25427),
	.a(n19075));
   in01f01 FE_OFC1298_n19075 (.o(FE_OFN264_n25427),
	.a(n19075));
   in01f01 FE_OFC1297_n19075 (.o(n19159),
	.a(n19075));
   in01f01 FE_OFC1296_n19075 (.o(n21864),
	.a(n19075));
   in01f01 FE_OFC1295_n19075 (.o(n25427),
	.a(n19075));
   in01f10 FE_OFC1294_n19075 (.o(n19192),
	.a(n19075));
   in01f06 FE_OFC1293_n21069 (.o(FE_OFN24767_n21069),
	.a(n21070));
   in01f08 FE_OFC1292_n21069 (.o(FE_OFN24766_n21069),
	.a(n21070));
   in01f01 FE_OFC1291_n21069 (.o(FE_OFN1100_n25937),
	.a(n21070));
   in01f01 FE_OFC1290_n21069 (.o(FE_OFN1098_n25937),
	.a(n21070));
   in01f01 FE_OFC1289_n21069 (.o(FE_OFN1099_n25937),
	.a(n21070));
   in01f01 FE_OFC1288_n21069 (.o(n25937),
	.a(n21070));
   in01f06 FE_OFC1287_n21069 (.o(n21070),
	.a(n21069));
   in01f10 FE_OFC1276_n20971 (.o(FE_OFN84_n20972),
	.a(n20972));
   in01f06 FE_OFC1275_n20971 (.o(n25905),
	.a(n20972));
   in01f06 FE_OFC1274_n20971 (.o(n20972),
	.a(n20971));
   in01f10 FE_OFC1273_n23045 (.o(n17767),
	.a(n23046));
   in01f08 FE_OFC1272_n23045 (.o(FE_OFN1081_n17767),
	.a(n23046));
   in01f01 FE_OFC1271_n23045 (.o(FE_OFN1080_n17767),
	.a(n23046));
   in01f01 FE_OFC1270_n23045 (.o(FE_OFN907_n23046),
	.a(n23046));
   in01f08 FE_OFC1269_n23045 (.o(n23046),
	.a(n23045));
   in01f06 FE_OFC1268_n23761 (.o(FE_OFN374_n17762),
	.a(n25571));
   in01f10 FE_OFC1267_n23761 (.o(FE_OFN373_n17762),
	.a(n25571));
   in01f01 FE_OFC1266_n23761 (.o(n17762),
	.a(n25571));
   in01f08 FE_OFC1265_n23761 (.o(n25571),
	.a(n23761));
   in01f01 FE_OFC1262_n23520 (.o(FE_OFN122_n23520),
	.a(n23520));
   in01f02 FE_OFC1256_n23735 (.o(n23788),
	.a(n23735));
   in01f06 FE_OFC1229_n21914 (.o(n23236),
	.a(n21915));
   in01f10 FE_OFC1228_n21914 (.o(FE_OFN448_n23236),
	.a(n21915));
   in01f06 FE_OFC1227_n21914 (.o(n21915),
	.a(n21914));
   in01f02 FE_OFC1226_n21051 (.o(n18632),
	.a(n21051));
   in01f02 FE_OFC1223_n21944 (.o(n23262),
	.a(FE_OFN452_n23262));
   in01f20 FE_OFC1211_north_input_NIB_head_ptr_f_0 (.o(n25109),
	.a(north_input_NIB_head_ptr_f_0_));
   in01f20 FE_OFC1210_n18683 (.o(FE_OFN24742_n18683),
	.a(n18683));
   in01f10 FE_OFC1209_n18683 (.o(FE_OFN24741_n18683),
	.a(n18683));
   in01f10 FE_OFC1208_n18683 (.o(n18060),
	.a(FE_RN_40));
   in01f20 FE_OFC1207_n18683 (.o(n17756),
	.a(FE_RN_40));
   in01f20 FE_OFC1206_n18683 (.o(n18061),
	.a(FE_RN_40));
   in01f08 FE_OFC1205_n21052 (.o(n21053),
	.a(n25945));
   in01f06 FE_OFC1204_n21052 (.o(n25945),
	.a(n21052));
   in01f20 FE_OFC1200_n20152 (.o(n20403),
	.a(n20152));
   in01f01 FE_OFC1198_n24998 (.o(FE_OFN945_n24998),
	.a(n24998));
   in01f20 FE_OFC1193_east_input_NIB_head_ptr_f_0 (.o(n18391),
	.a(east_input_NIB_head_ptr_f_0_));
   in01f08 FE_OFC1178_n20655 (.o(FE_OFN1087_n20656),
	.a(n20656));
   in01f02 FE_OFC1177_n20655 (.o(n25842),
	.a(n20656));
   in01f06 FE_OFC1176_n20655 (.o(n20656),
	.a(n20655));
   in01f01 FE_OFC1172_n21910 (.o(n23246),
	.a(FE_OFN25626_n21910));
   in01f10 FE_OFC1170_n23050 (.o(n23051),
	.a(FE_OFN440_n23051));
   in01m06 FE_OFC1169_n23050 (.o(FE_OFN442_n23051),
	.a(FE_OFN440_n23051));
   in01f08 FE_OFC1168_n23050 (.o(FE_OFN440_n23051),
	.a(n23050));
   in01f08 FE_OFC1162_n21219 (.o(FE_OFN88_n21220),
	.a(n21220));
   in01f08 FE_OFC1161_n21219 (.o(n25848),
	.a(n21220));
   in01f06 FE_OFC1160_n21219 (.o(n21220),
	.a(n21219));
   in01f06 FE_OFC1151_n21174 (.o(FE_OFN86_n21175),
	.a(n21175));
   in01f08 FE_OFC1150_n21174 (.o(n25836),
	.a(n21175));
   in01f06 FE_OFC1149_n21174 (.o(n21175),
	.a(n21174));
   in01f08 FE_OFC1148_n23737 (.o(FE_OFN272_n25595),
	.a(n25595));
   in01f10 FE_OFC1147_n23737 (.o(n17764),
	.a(n25595));
   in01f08 FE_OFC1146_n23737 (.o(n25595),
	.a(n23737));
   in01f02 FE_OFC1135_n20796 (.o(n17770),
	.a(n20797));
   in01f04 FE_OFC1134_n20796 (.o(FE_OFN899_n17770),
	.a(n20797));
   in01f06 FE_OFC1133_n20796 (.o(n20797),
	.a(n20796));
   in01f02 FE_OFC1128_n19306 (.o(FE_OFN24733_n19306),
	.a(FE_RN_69));
   in01f02 FE_OFC1126_n19306 (.o(n21857),
	.a(FE_OCPN25906_n19306));
   in01f02 FE_OFC1125_n19306 (.o(FE_OFN61_n19435),
	.a(FE_OCPN25906_n19306));
   in01f02 FE_OFC1124_n19306 (.o(FE_OFN59_n19435),
	.a(FE_OFN24737_n19306));
   in01f01 FE_OFC1123_n19306 (.o(FE_OFN58_n19435),
	.a(FE_OFN24732_n19306));
   in01f02 FE_OFC1122_n19306 (.o(n19933),
	.a(FE_OCPN25907_n19306));
   in01f06 FE_OFC1121_n19306 (.o(FE_OFN60_n19435),
	.a(FE_OCPN25907_n19306));
   in01f06 FE_OFC1120_n19306 (.o(n19435),
	.a(FE_OFN24735_n19306));
   in01f10 FE_OFC1119_n20814 (.o(FE_OFN952_n25916),
	.a(FE_OFN83_n20814));
   in01f06 FE_OFC1118_n20814 (.o(FE_OFN403_n20815),
	.a(FE_OFN83_n20814));
   in01f01 FE_OFC1117_n20814 (.o(n25916),
	.a(FE_OFN83_n20814));
   in01f01 FE_OFC1116_n20814 (.o(n20815),
	.a(FE_OFN83_n20814));
   in01f01 FE_OFC1115_n20814 (.o(FE_OFN82_n20814),
	.a(FE_OFN83_n20814));
   in01f01 FE_OFC1114_n20814 (.o(FE_OFN953_n25916),
	.a(FE_OFN83_n20814));
   in01f06 FE_OFC1113_n20814 (.o(FE_OFN83_n20814),
	.a(n20814));
   in01f10 FE_OFC1112_n22273 (.o(FE_OFN585_n25643),
	.a(n25643));
   in01f06 FE_OFC1111_n22273 (.o(n17768),
	.a(n25643));
   in01f02 FE_OFC1110_n22273 (.o(FE_OFN584_n25643),
	.a(n25643));
   in01f06 FE_OFC1109_n22273 (.o(n25643),
	.a(n22273));
   in01f40 FE_OFC1105_n18131 (.o(n24342),
	.a(n18131));
   in01f01 FE_OFC1104_n24728 (.o(FE_OFN24730_n),
	.a(FE_OFN24729_n));
   in01f01 FE_OFC1103_n24728 (.o(FE_OFN24729_n),
	.a(FE_OFN524_n24728));
   in01f01 FE_OFC1072_dataOut_P_2 (.o(FE_OFN1073_dataOut_P_2),
	.a(FE_OFN1072_dataOut_P_2));
   in01f02 FE_OFC1071_dataOut_P_3 (.o(dataOut_P_3_),
	.a(FE_OFN1071_dataOut_P_3));
   in01f02 FE_OFC1070_dataOut_P_3 (.o(FE_OFN1071_dataOut_P_3),
	.a(FE_OFN1070_dataOut_P_3));
   in01f02 FE_OFC1068_dataOut_P_4 (.o(FE_OFN1069_dataOut_P_4),
	.a(FE_OFN1068_dataOut_P_4));
   in01f02 FE_OFC1066_dataOut_P_5 (.o(FE_OFN1067_dataOut_P_5),
	.a(FE_OFN1066_dataOut_P_5));
   in01f02 FE_OFC1065_dataOut_P_7 (.o(dataOut_P_7_),
	.a(FE_OFN1065_dataOut_P_7));
   in01f02 FE_OFC1064_dataOut_P_7 (.o(FE_OFN1065_dataOut_P_7),
	.a(FE_OFN1064_dataOut_P_7));
   in01f02 FE_OFC1063_dataOut_P_8 (.o(dataOut_P_8_),
	.a(FE_OFN1063_dataOut_P_8));
   in01f02 FE_OFC1062_dataOut_P_8 (.o(FE_OFN1063_dataOut_P_8),
	.a(FE_OFN1062_dataOut_P_8));
   in01f02 FE_OFC1059_dataOut_P_12 (.o(dataOut_P_12_),
	.a(FE_OFN1059_dataOut_P_12));
   in01f02 FE_OFC1058_dataOut_P_12 (.o(FE_OFN1059_dataOut_P_12),
	.a(FE_OFN1058_dataOut_P_12));
   in01f02 FE_OFC1057_dataOut_P_14 (.o(dataOut_P_14_),
	.a(FE_OFN1057_dataOut_P_14));
   in01f02 FE_OFC1056_dataOut_P_14 (.o(FE_OFN1057_dataOut_P_14),
	.a(FE_OFN1056_dataOut_P_14));
   in01f02 FE_OFC1055_dataOut_P_18 (.o(dataOut_P_18_),
	.a(FE_OFN1055_dataOut_P_18));
   in01f02 FE_OFC1054_dataOut_P_18 (.o(FE_OFN1055_dataOut_P_18),
	.a(FE_OFN1054_dataOut_P_18));
   in01f02 FE_OFC1050_dataOut_W_2 (.o(FE_OFN1051_dataOut_W_2),
	.a(FE_OFN1050_dataOut_W_2));
   in01f02 FE_OFC1049_dataOut_W_3 (.o(dataOut_W_3_),
	.a(FE_OFN1049_dataOut_W_3));
   in01f02 FE_OFC1048_dataOut_W_3 (.o(FE_OFN1049_dataOut_W_3),
	.a(FE_OFN1048_dataOut_W_3));
   in01f01 FE_OFC1046_dataOut_W_4 (.o(FE_OFN1047_dataOut_W_4),
	.a(FE_OFN1046_dataOut_W_4));
   in01f02 FE_OFC1044_dataOut_W_5 (.o(FE_OFN1045_dataOut_W_5),
	.a(FE_OFN1044_dataOut_W_5));
   in01f02 FE_OFC1043_dataOut_W_7 (.o(dataOut_W_7_),
	.a(FE_OFN1043_dataOut_W_7));
   in01f02 FE_OFC1042_dataOut_W_7 (.o(FE_OFN1043_dataOut_W_7),
	.a(FE_OFN1042_dataOut_W_7));
   in01f02 FE_OFC1041_dataOut_W_8 (.o(dataOut_W_8_),
	.a(FE_OFN1041_dataOut_W_8));
   in01f02 FE_OFC1040_dataOut_W_8 (.o(FE_OFN1041_dataOut_W_8),
	.a(FE_OFN1040_dataOut_W_8));
   in01f02 FE_OFC1037_dataOut_W_12 (.o(dataOut_W_12_),
	.a(FE_OFN1037_dataOut_W_12));
   in01f02 FE_OFC1036_dataOut_W_12 (.o(FE_OFN1037_dataOut_W_12),
	.a(FE_OFN1036_dataOut_W_12));
   in01f02 FE_OFC1035_dataOut_W_14 (.o(dataOut_W_14_),
	.a(FE_OFN1035_dataOut_W_14));
   in01f02 FE_OFC1034_dataOut_W_14 (.o(FE_OFN1035_dataOut_W_14),
	.a(FE_OFN1034_dataOut_W_14));
   in01f01 FE_OFC1033_dataOut_W_18 (.o(dataOut_W_18_),
	.a(FE_OFN1033_dataOut_W_18));
   in01f02 FE_OFC1032_dataOut_W_18 (.o(FE_OFN1033_dataOut_W_18),
	.a(FE_OFN1032_dataOut_W_18));
   in01f02 FE_OFC1026_dataOut_S_2 (.o(FE_OFN1027_dataOut_S_2),
	.a(FE_OFN1026_dataOut_S_2));
   in01f02 FE_OFC1025_dataOut_S_3 (.o(dataOut_S_3_),
	.a(FE_OFN1025_dataOut_S_3));
   in01f02 FE_OFC1024_dataOut_S_3 (.o(FE_OFN1025_dataOut_S_3),
	.a(FE_OFN1024_dataOut_S_3));
   in01f01 FE_OFC1022_dataOut_S_4 (.o(FE_OFN1023_dataOut_S_4),
	.a(FE_OFN1022_dataOut_S_4));
   in01f02 FE_OFC1020_dataOut_S_5 (.o(FE_OFN1021_dataOut_S_5),
	.a(FE_OFN1020_dataOut_S_5));
   in01f01 FE_OFC1018_dataOut_S_7 (.o(FE_OFN1019_dataOut_S_7),
	.a(FE_OFN1018_dataOut_S_7));
   in01f01 FE_OFC1016_dataOut_S_8 (.o(FE_OFN1017_dataOut_S_8),
	.a(FE_OFN1016_dataOut_S_8));
   in01f02 FE_OFC1015_dataOut_S_9 (.o(dataOut_S_9_),
	.a(FE_OFN1015_dataOut_S_9));
   in01f01 FE_OFC1014_dataOut_S_9 (.o(FE_OFN1015_dataOut_S_9),
	.a(FE_OFN1014_dataOut_S_9));
   in01f01 FE_OFC1012_dataOut_S_12 (.o(FE_OFN1013_dataOut_S_12),
	.a(FE_OFN1012_dataOut_S_12));
   in01f02 FE_OFC1011_dataOut_S_14 (.o(dataOut_S_14_),
	.a(FE_OFN1011_dataOut_S_14));
   in01f02 FE_OFC1010_dataOut_S_14 (.o(FE_OFN1011_dataOut_S_14),
	.a(FE_OFN1010_dataOut_S_14));
   in01f01 FE_OFC1009_dataOut_S_18 (.o(dataOut_S_18_),
	.a(FE_OFN1009_dataOut_S_18));
   in01f02 FE_OFC1008_dataOut_S_18 (.o(FE_OFN1009_dataOut_S_18),
	.a(FE_OFN1008_dataOut_S_18));
   in01f01 FE_OFC1006_dataOut_S_31 (.o(FE_OFN1007_dataOut_S_31),
	.a(FE_OFN1006_dataOut_S_31));
   in01f02 FE_OFC1004_dataOut_E_2 (.o(FE_OFN1005_dataOut_E_2),
	.a(FE_OFN1004_dataOut_E_2));
   in01f02 FE_OFC1003_dataOut_E_3 (.o(dataOut_E_3_),
	.a(FE_OFN1003_dataOut_E_3));
   in01f02 FE_OFC1002_dataOut_E_3 (.o(FE_OFN1003_dataOut_E_3),
	.a(FE_OFN1002_dataOut_E_3));
   in01f01 FE_OFC1000_dataOut_E_4 (.o(FE_OFN1001_dataOut_E_4),
	.a(FE_OFN1000_dataOut_E_4));
   in01f02 FE_OFC998_dataOut_E_5 (.o(FE_OFN999_dataOut_E_5),
	.a(FE_OFN998_dataOut_E_5));
   in01f02 FE_OFC997_dataOut_E_7 (.o(dataOut_E_7_),
	.a(FE_OFN997_dataOut_E_7));
   in01f02 FE_OFC996_dataOut_E_7 (.o(FE_OFN997_dataOut_E_7),
	.a(FE_OFN996_dataOut_E_7));
   in01f02 FE_OFC993_dataOut_E_9 (.o(dataOut_E_9_),
	.a(FE_OFN993_dataOut_E_9));
   in01f02 FE_OFC992_dataOut_E_9 (.o(FE_OFN993_dataOut_E_9),
	.a(FE_OFN992_dataOut_E_9));
   in01f01 FE_OFC991_dataOut_E_12 (.o(dataOut_E_12_),
	.a(FE_OFN991_dataOut_E_12));
   in01f02 FE_OFC990_dataOut_E_12 (.o(FE_OFN991_dataOut_E_12),
	.a(FE_OFN990_dataOut_E_12));
   in01f01 FE_OFC988_dataOut_E_14 (.o(FE_OFN989_dataOut_E_14),
	.a(FE_OFN988_dataOut_E_14));
   in01f01 FE_OFC987_dataOut_E_18 (.o(dataOut_E_18_),
	.a(FE_OFN987_dataOut_E_18));
   in01f02 FE_OFC986_dataOut_E_18 (.o(FE_OFN987_dataOut_E_18),
	.a(FE_OFN986_dataOut_E_18));
   in01f01 FE_OFC980_dataOut_N_2 (.o(FE_OFN981_dataOut_N_2),
	.a(FE_OFN980_dataOut_N_2));
   in01f02 FE_OFC979_dataOut_N_3 (.o(dataOut_N_3_),
	.a(FE_OFN979_dataOut_N_3));
   in01f02 FE_OFC978_dataOut_N_3 (.o(FE_OFN979_dataOut_N_3),
	.a(FE_OFN978_dataOut_N_3));
   in01f01 FE_OFC976_dataOut_N_4 (.o(FE_OFN977_dataOut_N_4),
	.a(FE_OFN976_dataOut_N_4));
   in01f02 FE_OFC974_dataOut_N_5 (.o(FE_OFN975_dataOut_N_5),
	.a(FE_OFN974_dataOut_N_5));
   in01f02 FE_OFC973_dataOut_N_7 (.o(dataOut_N_7_),
	.a(FE_OFN973_dataOut_N_7));
   in01f02 FE_OFC972_dataOut_N_7 (.o(FE_OFN973_dataOut_N_7),
	.a(FE_OFN972_dataOut_N_7));
   in01f01 FE_OFC971_dataOut_N_8 (.o(dataOut_N_8_),
	.a(FE_OFN971_dataOut_N_8));
   in01f02 FE_OFC970_dataOut_N_8 (.o(FE_OFN971_dataOut_N_8),
	.a(FE_OFN970_dataOut_N_8));
   in01f02 FE_OFC969_dataOut_N_9 (.o(dataOut_N_9_),
	.a(FE_OFN969_dataOut_N_9));
   in01f02 FE_OFC968_dataOut_N_9 (.o(FE_OFN969_dataOut_N_9),
	.a(FE_OFN968_dataOut_N_9));
   in01f02 FE_OFC967_dataOut_N_12 (.o(dataOut_N_12_),
	.a(FE_OFN967_dataOut_N_12));
   in01f01 FE_OFC966_dataOut_N_12 (.o(FE_OFN967_dataOut_N_12),
	.a(FE_OFN966_dataOut_N_12));
   in01f02 FE_OFC965_dataOut_N_14 (.o(dataOut_N_14_),
	.a(FE_OFN965_dataOut_N_14));
   in01f02 FE_OFC964_dataOut_N_14 (.o(FE_OFN965_dataOut_N_14),
	.a(FE_OFN964_dataOut_N_14));
   in01f01 FE_OFC963_dataOut_N_18 (.o(dataOut_N_18_),
	.a(FE_OFN963_dataOut_N_18));
   in01f02 FE_OFC962_dataOut_N_18 (.o(FE_OFN963_dataOut_N_18),
	.a(FE_OFN962_dataOut_N_18));
   in01f02 FE_OFC959_n25972 (.o(FE_OFN959_n25972),
	.a(FE_OFN958_n25972));
   in01f01 FE_OFC958_n25972 (.o(FE_OFN958_n25972),
	.a(n25972));
   in01f01 FE_OFC951_n25881 (.o(FE_OFN951_n25881),
	.a(FE_OFN950_n25881));
   in01f01 FE_OFC950_n25881 (.o(FE_OFN950_n25881),
	.a(n25881));
   in01f03 FE_OFC943_n24921 (.o(FE_OFN943_n24921),
	.a(FE_OFN941_n24921));
   in01f01 FE_OFC941_n24921 (.o(FE_OFN941_n24921),
	.a(n24921));
   in01f01 FE_OFC934_n24710 (.o(FE_OFN934_n24710),
	.a(n24710));
   in01f02 FE_OFC922_n23576 (.o(FE_OFN922_n23576),
	.a(n23576));
   in01f01 FE_OFC906_n21586 (.o(FE_OFN906_n21586),
	.a(FE_OFN905_n21586));
   in01f01 FE_OFC905_n21586 (.o(FE_OFN905_n21586),
	.a(n21586));
   in01f01 FE_OFC904_n20750 (.o(FE_OFN904_n20750),
	.a(FE_OFN903_n20750));
   in01f01 FE_OFC903_n20750 (.o(FE_OFN903_n20750),
	.a(n20750));
   in01f01 FE_OFC884_dataOut_P_0 (.o(dataOut_P_0_),
	.a(FE_OFN884_dataOut_P_0));
   in01f02 FE_OFC883_dataOut_P_0 (.o(FE_OFN884_dataOut_P_0),
	.a(FE_OFN883_dataOut_P_0));
   in01f02 FE_OFC882_dataOut_P_1 (.o(dataOut_P_1_),
	.a(FE_OFN882_dataOut_P_1));
   in01f02 FE_OFC881_dataOut_P_1 (.o(FE_OFN882_dataOut_P_1),
	.a(FE_OFN881_dataOut_P_1));
   in01f02 FE_OFC880_dataOut_P_6 (.o(dataOut_P_6_),
	.a(FE_OFN880_dataOut_P_6));
   in01f02 FE_OFC879_dataOut_P_6 (.o(FE_OFN880_dataOut_P_6),
	.a(FE_OFN879_dataOut_P_6));
   in01f01 FE_OFC877_dataOut_P_10 (.o(FE_OFN878_dataOut_P_10),
	.a(FE_OFN877_dataOut_P_10));
   in01f02 FE_OFC875_dataOut_P_11 (.o(FE_OFN876_dataOut_P_11),
	.a(FE_OFN875_dataOut_P_11));
   in01f02 FE_OFC873_dataOut_P_13 (.o(FE_OFN874_dataOut_P_13),
	.a(FE_OFN873_dataOut_P_13));
   in01f02 FE_OFC872_dataOut_P_15 (.o(dataOut_P_15_),
	.a(FE_OFN872_dataOut_P_15));
   in01f02 FE_OFC871_dataOut_P_15 (.o(FE_OFN872_dataOut_P_15),
	.a(FE_OFN871_dataOut_P_15));
   in01f01 FE_OFC870_dataOut_P_16 (.o(dataOut_P_16_),
	.a(FE_OFN870_dataOut_P_16));
   in01f02 FE_OFC869_dataOut_P_16 (.o(FE_OFN870_dataOut_P_16),
	.a(FE_OFN869_dataOut_P_16));
   in01f02 FE_OFC867_dataOut_P_17 (.o(FE_OFN868_dataOut_P_17),
	.a(FE_OFN867_dataOut_P_17));
   in01f02 FE_OFC865_dataOut_P_19 (.o(FE_OFN866_dataOut_P_19),
	.a(FE_OFN865_dataOut_P_19));
   in01f02 FE_OFC864_dataOut_P_20 (.o(dataOut_P_20_),
	.a(FE_OFN864_dataOut_P_20));
   in01f02 FE_OFC863_dataOut_P_20 (.o(FE_OFN864_dataOut_P_20),
	.a(FE_OFN863_dataOut_P_20));
   in01f02 FE_OFC862_dataOut_P_21 (.o(dataOut_P_21_),
	.a(FE_OFN862_dataOut_P_21));
   in01f02 FE_OFC861_dataOut_P_21 (.o(FE_OFN862_dataOut_P_21),
	.a(FE_OFN861_dataOut_P_21));
   in01f01 FE_OFC857_dataOut_P_23 (.o(FE_OFN858_dataOut_P_23),
	.a(FE_OFN857_dataOut_P_23));
   in01f01 FE_OFC855_dataOut_P_24 (.o(FE_OFN856_dataOut_P_24),
	.a(FE_OFN855_dataOut_P_24));
   in01f02 FE_OFC854_dataOut_P_25 (.o(dataOut_P_25_),
	.a(FE_OFN854_dataOut_P_25));
   in01f02 FE_OFC853_dataOut_P_25 (.o(FE_OFN854_dataOut_P_25),
	.a(FE_OFN853_dataOut_P_25));
   in01f01 FE_OFC847_dataOut_P_28 (.o(FE_OFN848_dataOut_P_28),
	.a(FE_OFN847_dataOut_P_28));
   in01f01 FE_OFC845_dataOut_P_29 (.o(FE_OFN846_dataOut_P_29),
	.a(FE_OFN845_dataOut_P_29));
   in01f02 FE_OFC843_dataOut_P_33 (.o(FE_OFN844_dataOut_P_33),
	.a(FE_OFN843_dataOut_P_33));
   in01f01 FE_OFC841_dataOut_P_34 (.o(FE_OFN842_dataOut_P_34),
	.a(FE_OFN841_dataOut_P_34));
   in01f01 FE_OFC837_dataOut_P_36 (.o(FE_OFN838_dataOut_P_36),
	.a(FE_OFN837_dataOut_P_36));
   in01f01 FE_OFC833_dataOut_P_38 (.o(FE_OFN834_dataOut_P_38),
	.a(FE_OFN833_dataOut_P_38));
   in01f01 FE_OFC831_dataOut_P_39 (.o(FE_OFN832_dataOut_P_39),
	.a(FE_OFN831_dataOut_P_39));
   in01f01 FE_OFC829_dataOut_P_42 (.o(FE_OFN830_dataOut_P_42),
	.a(FE_OFN829_dataOut_P_42));
   in01f01 FE_OFC827_dataOut_P_43 (.o(FE_OFN828_dataOut_P_43),
	.a(FE_OFN827_dataOut_P_43));
   in01f02 FE_OFC810_dataOut_W_0 (.o(dataOut_W_0_),
	.a(FE_OFN810_dataOut_W_0));
   in01f02 FE_OFC809_dataOut_W_0 (.o(FE_OFN810_dataOut_W_0),
	.a(FE_OFN809_dataOut_W_0));
   in01f02 FE_OFC808_dataOut_W_1 (.o(dataOut_W_1_),
	.a(FE_OFN808_dataOut_W_1));
   in01f02 FE_OFC807_dataOut_W_1 (.o(FE_OFN808_dataOut_W_1),
	.a(FE_OFN807_dataOut_W_1));
   in01f02 FE_OFC805_dataOut_W_6 (.o(FE_OFN806_dataOut_W_6),
	.a(FE_OFN805_dataOut_W_6));
   in01f01 FE_OFC803_dataOut_W_10 (.o(FE_OFN804_dataOut_W_10),
	.a(FE_OFN803_dataOut_W_10));
   in01f02 FE_OFC801_dataOut_W_11 (.o(FE_OFN802_dataOut_W_11),
	.a(FE_OFN801_dataOut_W_11));
   in01f02 FE_OFC800_dataOut_W_13 (.o(dataOut_W_13_),
	.a(FE_OFN800_dataOut_W_13));
   in01f02 FE_OFC799_dataOut_W_13 (.o(FE_OFN800_dataOut_W_13),
	.a(FE_OFN799_dataOut_W_13));
   in01f01 FE_OFC798_dataOut_W_15 (.o(dataOut_W_15_),
	.a(FE_OFN798_dataOut_W_15));
   in01f02 FE_OFC797_dataOut_W_15 (.o(FE_OFN798_dataOut_W_15),
	.a(FE_OFN797_dataOut_W_15));
   in01f02 FE_OFC796_dataOut_W_16 (.o(dataOut_W_16_),
	.a(FE_OFN796_dataOut_W_16));
   in01f02 FE_OFC795_dataOut_W_16 (.o(FE_OFN796_dataOut_W_16),
	.a(FE_OFN795_dataOut_W_16));
   in01f02 FE_OFC793_dataOut_W_17 (.o(FE_OFN794_dataOut_W_17),
	.a(FE_OFN793_dataOut_W_17));
   in01f02 FE_OFC791_dataOut_W_19 (.o(FE_OFN792_dataOut_W_19),
	.a(FE_OFN791_dataOut_W_19));
   in01f02 FE_OFC790_dataOut_W_20 (.o(dataOut_W_20_),
	.a(FE_OFN790_dataOut_W_20));
   in01f02 FE_OFC789_dataOut_W_20 (.o(FE_OFN790_dataOut_W_20),
	.a(FE_OFN789_dataOut_W_20));
   in01f02 FE_OFC788_dataOut_W_21 (.o(dataOut_W_21_),
	.a(FE_OFN788_dataOut_W_21));
   in01f02 FE_OFC787_dataOut_W_21 (.o(FE_OFN788_dataOut_W_21),
	.a(FE_OFN787_dataOut_W_21));
   in01f01 FE_OFC783_dataOut_W_23 (.o(FE_OFN784_dataOut_W_23),
	.a(FE_OFN783_dataOut_W_23));
   in01f01 FE_OFC781_dataOut_W_24 (.o(FE_OFN782_dataOut_W_24),
	.a(FE_OFN781_dataOut_W_24));
   in01f02 FE_OFC780_dataOut_W_25 (.o(dataOut_W_25_),
	.a(FE_OFN780_dataOut_W_25));
   in01f02 FE_OFC779_dataOut_W_25 (.o(FE_OFN780_dataOut_W_25),
	.a(FE_OFN779_dataOut_W_25));
   in01f01 FE_OFC776_dataOut_W_27 (.o(dataOut_W_27_),
	.a(FE_OFN776_dataOut_W_27));
   in01f01 FE_OFC775_dataOut_W_27 (.o(FE_OFN776_dataOut_W_27),
	.a(FE_OFN775_dataOut_W_27));
   in01f01 FE_OFC773_dataOut_W_28 (.o(FE_OFN774_dataOut_W_28),
	.a(FE_OFN773_dataOut_W_28));
   in01f01 FE_OFC769_dataOut_W_33 (.o(FE_OFN770_dataOut_W_33),
	.a(FE_OFN769_dataOut_W_33));
   in01f01 FE_OFC767_dataOut_W_34 (.o(FE_OFN768_dataOut_W_34),
	.a(FE_OFN767_dataOut_W_34));
   in01f01 FE_OFC763_dataOut_W_36 (.o(FE_OFN764_dataOut_W_36),
	.a(FE_OFN763_dataOut_W_36));
   in01f01 FE_OFC759_dataOut_W_38 (.o(FE_OFN760_dataOut_W_38),
	.a(FE_OFN759_dataOut_W_38));
   in01f01 FE_OFC757_dataOut_W_39 (.o(FE_OFN758_dataOut_W_39),
	.a(FE_OFN757_dataOut_W_39));
   in01f01 FE_OFC755_dataOut_W_42 (.o(FE_OFN756_dataOut_W_42),
	.a(FE_OFN755_dataOut_W_42));
   in01f01 FE_OFC747_dataOut_W_46 (.o(FE_OFN748_dataOut_W_46),
	.a(FE_OFN747_dataOut_W_46));
   in01f02 FE_OFC734_dataOut_S_0 (.o(dataOut_S_0_),
	.a(FE_OFN734_dataOut_S_0));
   in01f02 FE_OFC733_dataOut_S_0 (.o(FE_OFN734_dataOut_S_0),
	.a(FE_OFN733_dataOut_S_0));
   in01f01 FE_OFC731_dataOut_S_1 (.o(FE_OFN732_dataOut_S_1),
	.a(FE_OFN731_dataOut_S_1));
   in01f02 FE_OFC729_dataOut_S_6 (.o(FE_OFN730_dataOut_S_6),
	.a(FE_OFN729_dataOut_S_6));
   in01f01 FE_OFC727_dataOut_S_10 (.o(FE_OFN728_dataOut_S_10),
	.a(FE_OFN727_dataOut_S_10));
   in01f02 FE_OFC725_dataOut_S_11 (.o(FE_OFN726_dataOut_S_11),
	.a(FE_OFN725_dataOut_S_11));
   in01f02 FE_OFC723_dataOut_S_13 (.o(FE_OFN724_dataOut_S_13),
	.a(FE_OFN723_dataOut_S_13));
   in01f01 FE_OFC721_dataOut_S_15 (.o(FE_OFN722_dataOut_S_15),
	.a(FE_OFN721_dataOut_S_15));
   in01f01 FE_OFC719_dataOut_S_16 (.o(FE_OFN720_dataOut_S_16),
	.a(FE_OFN719_dataOut_S_16));
   in01f02 FE_OFC717_dataOut_S_17 (.o(FE_OFN718_dataOut_S_17),
	.a(FE_OFN717_dataOut_S_17));
   in01f01 FE_OFC715_dataOut_S_19 (.o(FE_OFN716_dataOut_S_19),
	.a(FE_OFN715_dataOut_S_19));
   in01f01 FE_OFC713_dataOut_S_20 (.o(FE_OFN714_dataOut_S_20),
	.a(FE_OFN713_dataOut_S_20));
   in01f02 FE_OFC712_dataOut_S_21 (.o(dataOut_S_21_),
	.a(FE_OFN712_dataOut_S_21));
   in01f02 FE_OFC711_dataOut_S_21 (.o(FE_OFN712_dataOut_S_21),
	.a(FE_OFN711_dataOut_S_21));
   in01f01 FE_OFC709_dataOut_S_22 (.o(FE_OFN710_dataOut_S_22),
	.a(FE_OFN709_dataOut_S_22));
   in01f01 FE_OFC707_dataOut_S_23 (.o(FE_OFN708_dataOut_S_23),
	.a(FE_OFN707_dataOut_S_23));
   in01f01 FE_OFC705_dataOut_S_24 (.o(FE_OFN706_dataOut_S_24),
	.a(FE_OFN705_dataOut_S_24));
   in01f01 FE_OFC703_dataOut_S_25 (.o(FE_OFN704_dataOut_S_25),
	.a(FE_OFN703_dataOut_S_25));
   in01f01 FE_OFC701_dataOut_S_26 (.o(FE_OFN702_dataOut_S_26),
	.a(FE_OFN701_dataOut_S_26));
   in01f01 FE_OFC700_dataOut_S_27 (.o(dataOut_S_27_),
	.a(FE_OFN700_dataOut_S_27));
   in01f02 FE_OFC699_dataOut_S_27 (.o(FE_OFN700_dataOut_S_27),
	.a(FE_OFN699_dataOut_S_27));
   in01f01 FE_OFC697_dataOut_S_28 (.o(FE_OFN698_dataOut_S_28),
	.a(FE_OFN697_dataOut_S_28));
   in01f01 FE_OFC695_dataOut_S_29 (.o(FE_OFN696_dataOut_S_29),
	.a(FE_OFN695_dataOut_S_29));
   in01f02 FE_OFC693_dataOut_S_33 (.o(FE_OFN694_dataOut_S_33),
	.a(FE_OFN693_dataOut_S_33));
   in01f01 FE_OFC691_dataOut_S_34 (.o(FE_OFN692_dataOut_S_34),
	.a(FE_OFN691_dataOut_S_34));
   in01f01 FE_OFC689_dataOut_S_35 (.o(FE_OFN690_dataOut_S_35),
	.a(FE_OFN689_dataOut_S_35));
   in01f01 FE_OFC687_dataOut_S_36 (.o(FE_OFN688_dataOut_S_36),
	.a(FE_OFN687_dataOut_S_36));
   in01f01 FE_OFC685_dataOut_S_37 (.o(FE_OFN686_dataOut_S_37),
	.a(FE_OFN685_dataOut_S_37));
   in01f01 FE_OFC683_dataOut_S_38 (.o(FE_OFN684_dataOut_S_38),
	.a(FE_OFN683_dataOut_S_38));
   in01f01 FE_OFC681_dataOut_S_39 (.o(FE_OFN682_dataOut_S_39),
	.a(FE_OFN681_dataOut_S_39));
   in01f01 FE_OFC679_dataOut_S_42 (.o(FE_OFN680_dataOut_S_42),
	.a(FE_OFN679_dataOut_S_42));
   in01f01 FE_OFC677_dataOut_S_43 (.o(FE_OFN678_dataOut_S_43),
	.a(FE_OFN677_dataOut_S_43));
   in01f01 FE_OFC665_dataOut_S_49 (.o(FE_OFN666_dataOut_S_49),
	.a(FE_OFN665_dataOut_S_49));
   in01f02 FE_OFC660_dataOut_E_0 (.o(dataOut_E_0_),
	.a(FE_OFN660_dataOut_E_0));
   in01f01 FE_OFC659_dataOut_E_0 (.o(FE_OFN660_dataOut_E_0),
	.a(FE_OFN659_dataOut_E_0));
   in01f02 FE_OFC655_dataOut_E_6 (.o(FE_OFN656_dataOut_E_6),
	.a(FE_OFN655_dataOut_E_6));
   in01f02 FE_OFC654_dataOut_E_10 (.o(dataOut_E_10_),
	.a(FE_OFN654_dataOut_E_10));
   in01f02 FE_OFC653_dataOut_E_10 (.o(FE_OFN654_dataOut_E_10),
	.a(FE_OFN653_dataOut_E_10));
   in01f01 FE_OFC651_dataOut_E_11 (.o(FE_OFN652_dataOut_E_11),
	.a(FE_OFN651_dataOut_E_11));
   in01f02 FE_OFC649_dataOut_E_13 (.o(FE_OFN650_dataOut_E_13),
	.a(FE_OFN649_dataOut_E_13));
   in01f02 FE_OFC648_dataOut_E_15 (.o(dataOut_E_15_),
	.a(FE_OFN648_dataOut_E_15));
   in01f02 FE_OFC647_dataOut_E_15 (.o(FE_OFN648_dataOut_E_15),
	.a(FE_OFN647_dataOut_E_15));
   in01f01 FE_OFC643_dataOut_E_17 (.o(FE_OFN644_dataOut_E_17),
	.a(FE_OFN643_dataOut_E_17));
   in01f02 FE_OFC641_dataOut_E_19 (.o(FE_OFN642_dataOut_E_19),
	.a(FE_OFN641_dataOut_E_19));
   in01f02 FE_OFC640_dataOut_E_20 (.o(dataOut_E_20_),
	.a(FE_OFN640_dataOut_E_20));
   in01f02 FE_OFC639_dataOut_E_20 (.o(FE_OFN640_dataOut_E_20),
	.a(FE_OFN639_dataOut_E_20));
   in01f02 FE_OFC638_dataOut_E_21 (.o(dataOut_E_21_),
	.a(FE_OFN638_dataOut_E_21));
   in01f02 FE_OFC637_dataOut_E_21 (.o(FE_OFN638_dataOut_E_21),
	.a(FE_OFN637_dataOut_E_21));
   in01f01 FE_OFC633_dataOut_E_23 (.o(FE_OFN634_dataOut_E_23),
	.a(FE_OFN633_dataOut_E_23));
   in01f01 FE_OFC631_dataOut_E_24 (.o(FE_OFN632_dataOut_E_24),
	.a(FE_OFN631_dataOut_E_24));
   in01f01 FE_OFC628_dataOut_E_27 (.o(dataOut_E_27_),
	.a(FE_OFN628_dataOut_E_27));
   in01f01 FE_OFC627_dataOut_E_27 (.o(FE_OFN628_dataOut_E_27),
	.a(FE_OFN627_dataOut_E_27));
   in01f01 FE_OFC625_dataOut_E_28 (.o(FE_OFN626_dataOut_E_28),
	.a(FE_OFN625_dataOut_E_28));
   in01f01 FE_OFC623_dataOut_E_29 (.o(FE_OFN624_dataOut_E_29),
	.a(FE_OFN623_dataOut_E_29));
   in01f02 FE_OFC621_dataOut_E_33 (.o(FE_OFN622_dataOut_E_33),
	.a(FE_OFN621_dataOut_E_33));
   in01f01 FE_OFC619_dataOut_E_34 (.o(FE_OFN620_dataOut_E_34),
	.a(FE_OFN619_dataOut_E_34));
   in01f01 FE_OFC615_dataOut_E_36 (.o(FE_OFN616_dataOut_E_36),
	.a(FE_OFN615_dataOut_E_36));
   in01f01 FE_OFC611_dataOut_E_38 (.o(FE_OFN612_dataOut_E_38),
	.a(FE_OFN611_dataOut_E_38));
   in01f01 FE_OFC607_dataOut_E_42 (.o(FE_OFN608_dataOut_E_42),
	.a(FE_OFN607_dataOut_E_42));
   in01f01 FE_OFC595_dataOut_N_27 (.o(FE_OFN596_dataOut_N_27),
	.a(FE_OFN595_dataOut_N_27));
   in01f01 FE_OFC579_n25511 (.o(FE_OFN579_n25511),
	.a(FE_OFN578_n25511));
   in01f01 FE_OFC578_n25511 (.o(FE_OFN578_n25511),
	.a(n25511));
   in01f04 FE_OFC577_n25498 (.o(FE_OFN577_n25498),
	.a(FE_OFN576_n25498));
   in01f02 FE_OFC576_n25498 (.o(FE_OFN576_n25498),
	.a(n25498));
   in01f06 FE_OFC575_n25463 (.o(FE_OFN575_n25463),
	.a(FE_OFN572_n25463));
   in01f01 FE_OFC573_n25463 (.o(FE_OFN573_n25463),
	.a(reset));
   in01f02 FE_OFC572_n25463 (.o(FE_OFN572_n25463),
	.a(FE_OFN25598_reset));
   in01f01 FE_OFC570_n25395 (.o(FE_OFN570_n25395),
	.a(FE_OFN567_n25395));
   in01f01 FE_OFC569_n25395 (.o(FE_OFN569_n25395),
	.a(FE_OFN566_n25395));
   in01f01 FE_OFC567_n25395 (.o(FE_OFN567_n25395),
	.a(FE_OFN25891_n25395));
   in01f01 FE_OFC566_n25395 (.o(FE_OFN566_n25395),
	.a(FE_OFN25891_n25395));
   in01f01 FE_OFC556_n24761 (.o(FE_OFN556_n24761),
	.a(FE_OFN554_n24761));
   in01f04 FE_OFC555_n24761 (.o(FE_OFN555_n24761),
	.a(FE_OFN553_n24761));
   in01f01 FE_OFC554_n24761 (.o(FE_OFN554_n24761),
	.a(n24761));
   in01f01 FE_OFC553_n24761 (.o(FE_OFN553_n24761),
	.a(n24761));
   in01f02 FE_OFC545_n24751 (.o(FE_OFN545_n24751),
	.a(n24751));
   in01f02 FE_OFC530_n24733 (.o(FE_OFN530_n24733),
	.a(FE_OFN529_n24733));
   in01f02 FE_OFC529_n24733 (.o(FE_OFN529_n24733),
	.a(n24733));
   in01f02 FE_OFC527_n24732 (.o(FE_OFN527_n24732),
	.a(n24732));
   in01f03 FE_OFC526_n24731 (.o(FE_OFN526_n24731),
	.a(FE_OFN25672_n22773));
   in01f04 FE_OFC524_n24728 (.o(FE_OFN524_n24728),
	.a(FE_OFN522_n24728));
   in01f01 FE_OFC523_n24728 (.o(FE_OFN523_n24728),
	.a(FE_OFN522_n24728));
   in01f01 FE_OFC522_n24728 (.o(FE_OFN522_n24728),
	.a(n24728));
   in01f02 FE_OFC521_n24723 (.o(FE_OFN521_n24723),
	.a(FE_OFN520_n24723));
   in01f01 FE_OFC520_n24723 (.o(FE_OFN520_n24723),
	.a(n24723));
   in01f02 FE_OFC517_n24712 (.o(FE_OFN517_n24712),
	.a(FE_OFN516_n24712));
   in01f01 FE_OFC516_n24712 (.o(FE_OFN516_n24712),
	.a(n24712));
   in01f02 FE_OFC515_n24702 (.o(FE_OFN515_n24702),
	.a(FE_OFN514_n24702));
   in01f02 FE_OFC514_n24702 (.o(FE_OFN514_n24702),
	.a(n24702));
   in01f02 FE_OFC513_n24695 (.o(FE_OFN513_n24695),
	.a(FE_OFN512_n24695));
   in01f01 FE_OFC512_n24695 (.o(FE_OFN512_n24695),
	.a(n24695));
   in01f01 FE_OFC498_n24601 (.o(FE_OFN498_n24601),
	.a(n24601));
   in01f02 FE_OFC497_n24586 (.o(FE_OFN497_n24586),
	.a(FE_OFN496_n24586));
   in01f01 FE_OFC496_n24586 (.o(FE_OFN496_n24586),
	.a(n24586));
   in01f02 FE_OFC494_n24579 (.o(FE_OFN494_n24579),
	.a(n24579));
   in01f02 FE_OFC493_n24577 (.o(FE_OFN493_n24577),
	.a(FE_OFN492_n24577));
   in01f01 FE_OFC492_n24577 (.o(FE_OFN492_n24577),
	.a(n24577));
   in01f02 FE_OFC491_n24022 (.o(FE_OFN491_n24022),
	.a(FE_OFN490_n24022));
   in01f02 FE_OFC490_n24022 (.o(FE_OFN490_n24022),
	.a(n24022));
   in01f02 FE_OFC487_n24013 (.o(FE_OFN487_n24013),
	.a(FE_OFN486_n24013));
   in01f01 FE_OFC486_n24013 (.o(FE_OFN486_n24013),
	.a(n24013));
   in01f02 FE_OFC484_n24011 (.o(FE_OFN484_n24011),
	.a(n24011));
   in01f01 FE_OFC483_n23987 (.o(FE_OFN483_n23987),
	.a(FE_OFN482_n23987));
   in01f02 FE_OFC482_n23987 (.o(FE_OFN482_n23987),
	.a(n23987));
   in01f02 FE_OFC479_n23631 (.o(FE_OFN479_n23631),
	.a(FE_OFN478_n23631));
   in01f01 FE_OFC478_n23631 (.o(FE_OFN478_n23631),
	.a(n23631));
   in01f02 FE_OFC477_n23578 (.o(FE_OFN477_n23578),
	.a(FE_OFN476_n23578));
   in01f02 FE_OFC476_n23578 (.o(FE_OFN476_n23578),
	.a(n23578));
   in01f02 FE_OFC473_n23560 (.o(FE_OFN473_n23560),
	.a(FE_OFN472_n23560));
   in01f01 FE_OFC472_n23560 (.o(FE_OFN472_n23560),
	.a(n23560));
   in01f01 FE_OFC437_n22958 (.o(FE_OFN437_n22958),
	.a(FE_OFN435_n22958));
   in01f04 FE_OFC436_n22958 (.o(FE_OFN436_n22958),
	.a(FE_OFN434_n22958));
   in01f01 FE_OFC434_n22958 (.o(FE_OFN434_n22958),
	.a(n22958));
   in01f04 FE_OFC432_n22945 (.o(FE_OFN432_n22945),
	.a(FE_OFN430_n22945));
   in01f01 FE_OFC430_n22945 (.o(FE_OFN430_n22945),
	.a(FE_OFN24860_n22945));
   in01f01 FE_OFC427_n22778 (.o(FE_OFN427_n22778),
	.a(FE_OFN425_n22778));
   in01f01 FE_OFC426_n22778 (.o(FE_OFN426_n22778),
	.a(FE_OFN425_n22778));
   in01f01 FE_OFC425_n22778 (.o(FE_OFN425_n22778),
	.a(n22778));
   in01f01 FE_OFC423_n22766 (.o(FE_OFN423_n22766),
	.a(n22766));
   in01f01 FE_OFC418_n22535 (.o(FE_OFN418_n22535),
	.a(FE_OFN417_n22535));
   in01f01 FE_OFC417_n22535 (.o(FE_OFN417_n22535),
	.a(n22535));
   in01f03 FE_OFC412_n21671 (.o(FE_OFN412_n21671),
	.a(FE_OFN411_n21671));
   in01f02 FE_OFC411_n21671 (.o(FE_OFN411_n21671),
	.a(n21671));
   in01f01 FE_OFC408_n21421 (.o(FE_OFN408_n21421),
	.a(FE_OFN407_n21421));
   in01f01 FE_OFC407_n21421 (.o(FE_OFN407_n21421),
	.a(n21421));
   in01f02 FE_OFC396_n19493 (.o(FE_OFN396_n19493),
	.a(FE_OFN395_n19493));
   in01f01 FE_OFC395_n19493 (.o(FE_OFN395_n19493),
	.a(n19493));
   in01f01 FE_OFC394_n19446 (.o(FE_OFN394_n19446),
	.a(FE_OFN391_n19446));
   in01f02 FE_OFC393_n19446 (.o(FE_OFN393_n19446),
	.a(FE_OFN390_n19446));
   in01f01 FE_OFC391_n19446 (.o(FE_OFN391_n19446),
	.a(FE_OFN25878_n19446));
   in01f01 FE_OFC390_n19446 (.o(FE_OFN390_n19446),
	.a(FE_OFN25880_n19446));
   in01f06 FE_OFC389_n17786 (.o(FE_OFN389_n17786),
	.a(FE_OFN388_n17786));
   in01f02 FE_OFC388_n17786 (.o(FE_OFN388_n17786),
	.a(n17786));
   in01f01 FE_OFC364_dataOut_P_40 (.o(FE_OFN365_dataOut_P_40),
	.a(FE_OFN364_dataOut_P_40));
   in01f01 FE_OFC362_dataOut_W_40 (.o(FE_OFN363_dataOut_W_40),
	.a(FE_OFN362_dataOut_W_40));
   in01f01 FE_OFC360_dataOut_S_40 (.o(FE_OFN361_dataOut_S_40),
	.a(FE_OFN360_dataOut_S_40));
   in01f01 FE_OFC354_dataOut_E_40 (.o(FE_OFN355_dataOut_E_40),
	.a(FE_OFN354_dataOut_E_40));
   in01f01 FE_OFC352_dataOut_E_43 (.o(FE_OFN353_dataOut_E_43),
	.a(FE_OFN352_dataOut_E_43));
   in01f02 FE_OFC343_dataOut_N_0 (.o(dataOut_N_0_),
	.a(FE_OFN343_dataOut_N_0));
   in01f02 FE_OFC342_dataOut_N_0 (.o(FE_OFN343_dataOut_N_0),
	.a(FE_OFN342_dataOut_N_0));
   in01f02 FE_OFC341_dataOut_N_1 (.o(dataOut_N_1_),
	.a(FE_OFN341_dataOut_N_1));
   in01f02 FE_OFC340_dataOut_N_1 (.o(FE_OFN341_dataOut_N_1),
	.a(FE_OFN340_dataOut_N_1));
   in01f02 FE_OFC338_dataOut_N_6 (.o(FE_OFN339_dataOut_N_6),
	.a(FE_OFN338_dataOut_N_6));
   in01f01 FE_OFC336_dataOut_N_10 (.o(FE_OFN337_dataOut_N_10),
	.a(FE_OFN336_dataOut_N_10));
   in01f02 FE_OFC334_dataOut_N_11 (.o(FE_OFN335_dataOut_N_11),
	.a(FE_OFN334_dataOut_N_11));
   in01f02 FE_OFC332_dataOut_N_13 (.o(FE_OFN333_dataOut_N_13),
	.a(FE_OFN332_dataOut_N_13));
   in01f01 FE_OFC330_dataOut_N_15 (.o(FE_OFN331_dataOut_N_15),
	.a(FE_OFN330_dataOut_N_15));
   in01f02 FE_OFC329_dataOut_N_16 (.o(dataOut_N_16_),
	.a(FE_OFN329_dataOut_N_16));
   in01f02 FE_OFC328_dataOut_N_16 (.o(FE_OFN329_dataOut_N_16),
	.a(FE_OFN328_dataOut_N_16));
   in01f02 FE_OFC326_dataOut_N_17 (.o(FE_OFN327_dataOut_N_17),
	.a(FE_OFN326_dataOut_N_17));
   in01f02 FE_OFC324_dataOut_N_19 (.o(FE_OFN325_dataOut_N_19),
	.a(FE_OFN324_dataOut_N_19));
   in01f02 FE_OFC323_dataOut_N_20 (.o(dataOut_N_20_),
	.a(FE_OFN323_dataOut_N_20));
   in01f01 FE_OFC322_dataOut_N_20 (.o(FE_OFN323_dataOut_N_20),
	.a(FE_OFN322_dataOut_N_20));
   in01f01 FE_OFC321_dataOut_N_21 (.o(dataOut_N_21_),
	.a(FE_OFN321_dataOut_N_21));
   in01f02 FE_OFC320_dataOut_N_21 (.o(FE_OFN321_dataOut_N_21),
	.a(FE_OFN320_dataOut_N_21));
   in01f01 FE_OFC316_dataOut_N_23 (.o(FE_OFN317_dataOut_N_23),
	.a(FE_OFN316_dataOut_N_23));
   in01f01 FE_OFC314_dataOut_N_24 (.o(FE_OFN315_dataOut_N_24),
	.a(FE_OFN314_dataOut_N_24));
   in01f01 FE_OFC312_dataOut_N_25 (.o(FE_OFN313_dataOut_N_25),
	.a(FE_OFN312_dataOut_N_25));
   in01f01 FE_OFC310_dataOut_N_28 (.o(FE_OFN311_dataOut_N_28),
	.a(FE_OFN310_dataOut_N_28));
   in01f01 FE_OFC308_dataOut_N_29 (.o(FE_OFN309_dataOut_N_29),
	.a(FE_OFN308_dataOut_N_29));
   in01f02 FE_OFC304_dataOut_N_33 (.o(FE_OFN305_dataOut_N_33),
	.a(FE_OFN304_dataOut_N_33));
   in01f01 FE_OFC302_dataOut_N_34 (.o(FE_OFN303_dataOut_N_34),
	.a(FE_OFN302_dataOut_N_34));
   in01f01 FE_OFC298_dataOut_N_36 (.o(FE_OFN299_dataOut_N_36),
	.a(FE_OFN298_dataOut_N_36));
   in01f01 FE_OFC294_dataOut_N_38 (.o(FE_OFN295_dataOut_N_38),
	.a(FE_OFN294_dataOut_N_38));
   in01f01 FE_OFC292_dataOut_N_39 (.o(FE_OFN293_dataOut_N_39),
	.a(FE_OFN292_dataOut_N_39));
   in01f01 FE_OFC290_dataOut_N_42 (.o(FE_OFN291_dataOut_N_42),
	.a(FE_OFN290_dataOut_N_42));
   in01f01 FE_OFC288_dataOut_N_43 (.o(FE_OFN289_dataOut_N_43),
	.a(FE_OFN288_dataOut_N_43));
   in01f04 FE_OFC269_n25506 (.o(FE_OFN269_n25506),
	.a(FE_OFN268_n25506));
   in01f02 FE_OFC268_n25506 (.o(FE_OFN268_n25506),
	.a(n25506));
   in01f01 FE_OFC262_n25301 (.o(FE_OFN262_n25301),
	.a(FE_OFN261_n25301));
   in01f01 FE_OFC261_n25301 (.o(FE_OFN261_n25301),
	.a(n25301));
   in01f01 FE_OFC260_n25295 (.o(FE_OFN260_n25295),
	.a(FE_OFN258_n25295));
   in01f04 FE_OFC259_n25295 (.o(FE_OFN259_n25295),
	.a(FE_OFN258_n25295));
   in01f02 FE_OFC258_n25295 (.o(FE_OFN258_n25295),
	.a(n25295));
   in01f02 FE_OFC257_n25294 (.o(FE_OFN257_n25294),
	.a(FE_OFN256_n25294));
   in01f01 FE_OFC256_n25294 (.o(FE_OFN256_n25294),
	.a(n25294));
   in01f01 FE_OFC255_n25247 (.o(FE_OFN255_n25247),
	.a(FE_OFN254_n25247));
   in01f01 FE_OFC254_n25247 (.o(FE_OFN254_n25247),
	.a(n25247));
   in01f01 FE_OFC253_n25241 (.o(FE_OFN253_n25241),
	.a(FE_OFN252_n25241));
   in01f01 FE_OFC252_n25241 (.o(FE_OFN252_n25241),
	.a(n25241));
   in01f01 FE_OFC251_n25152 (.o(FE_OFN251_n25152),
	.a(FE_OFN249_n25152));
   in01f01 FE_OFC250_n25152 (.o(FE_OFN250_n25152),
	.a(FE_OFN248_n25152));
   in01f01 FE_OFC249_n25152 (.o(FE_OFN249_n25152),
	.a(n25152));
   in01f01 FE_OFC248_n25152 (.o(FE_OFN248_n25152),
	.a(n25152));
   in01f08 FE_OFC247_n24982 (.o(FE_OFN247_n24982),
	.a(FE_OFN246_n24982));
   in01f02 FE_OFC246_n24982 (.o(FE_OFN246_n24982),
	.a(n24982));
   in01f02 FE_OFC242_n24744 (.o(FE_OFN242_n24744),
	.a(FE_OFN241_n24744));
   in01f02 FE_OFC241_n24744 (.o(FE_OFN241_n24744),
	.a(n24744));
   in01f02 FE_OFC238_n24739 (.o(FE_OFN238_n24739),
	.a(n24739));
   in01f02 FE_OFC237_n24730 (.o(FE_OFN237_n24730),
	.a(FE_OFN236_n24730));
   in01f02 FE_OFC236_n24730 (.o(FE_OFN236_n24730),
	.a(n24730));
   in01f02 FE_OFC234_n24729 (.o(FE_OFN234_n24729),
	.a(n24729));
   in01f02 FE_OFC232_n24719 (.o(FE_OFN232_n24719),
	.a(n24719));
   in01f01 FE_OFC230_n24704 (.o(FE_OFN230_n24704),
	.a(n24704));
   in01f02 FE_OFC229_n24684 (.o(FE_OFN229_n24684),
	.a(FE_OFN228_n24684));
   in01f02 FE_OFC228_n24684 (.o(FE_OFN228_n24684),
	.a(n24684));
   in01f02 FE_OFC227_n24677 (.o(FE_OFN227_n24677),
	.a(FE_OFN226_n24677));
   in01f01 FE_OFC226_n24677 (.o(FE_OFN226_n24677),
	.a(n24677));
   in01f02 FE_OFC223_n24664 (.o(FE_OFN223_n24664),
	.a(FE_OFN222_n24664));
   in01f01 FE_OFC222_n24664 (.o(FE_OFN222_n24664),
	.a(n24664));
   in01f03 FE_OFC221_n24662 (.o(FE_OFN221_n24662),
	.a(FE_OFN220_n24662));
   in01f02 FE_OFC220_n24662 (.o(FE_OFN220_n24662),
	.a(n24662));
   in01f02 FE_OFC218_n24645 (.o(FE_OFN218_n24645),
	.a(n24645));
   in01f02 FE_OFC217_n24637 (.o(FE_OFN217_n24637),
	.a(FE_OFN216_n24637));
   in01f01 FE_OFC216_n24637 (.o(FE_OFN216_n24637),
	.a(n24637));
   in01f02 FE_OFC214_n24636 (.o(FE_OFN214_n24636),
	.a(n24636));
   in01f01 FE_OFC210_n24630 (.o(FE_OFN210_n24630),
	.a(n24630));
   in01f02 FE_OFC207_n24619 (.o(FE_OFN207_n24619),
	.a(FE_OFN206_n24619));
   in01f01 FE_OFC206_n24619 (.o(FE_OFN206_n24619),
	.a(n24619));
   in01f02 FE_OFC203_n24600 (.o(FE_OFN203_n24600),
	.a(FE_OFN202_n24600));
   in01f02 FE_OFC202_n24600 (.o(FE_OFN202_n24600),
	.a(n24600));
   in01f02 FE_OFC200_n24584 (.o(FE_OFN200_n24584),
	.a(n24584));
   in01f01 FE_OFC154_n24036 (.o(FE_OFN154_n24036),
	.a(n24036));
   in01f02 FE_OFC152_n24027 (.o(FE_OFN152_n24027),
	.a(n24027));
   in01f02 FE_OFC151_n24019 (.o(FE_OFN151_n24019),
	.a(FE_OFN150_n24019));
   in01f02 FE_OFC150_n24019 (.o(FE_OFN150_n24019),
	.a(n24019));
   in01f02 FE_OFC146_n24010 (.o(FE_OFN146_n24010),
	.a(FE_OFN145_n24010));
   in01f02 FE_OFC145_n24010 (.o(FE_OFN145_n24010),
	.a(n24010));
   in01f01 FE_OFC143_n23991 (.o(FE_OFN143_n23991),
	.a(n23991));
   in01f01 FE_OFC141_n23964 (.o(FE_OFN141_n23964),
	.a(n23964));
   in01f02 FE_OFC140_n23959 (.o(FE_OFN140_n23959),
	.a(FE_OFN139_n23959));
   in01f01 FE_OFC139_n23959 (.o(FE_OFN139_n23959),
	.a(n23959));
   in01f02 FE_OFC138_n23948 (.o(FE_OFN138_n23948),
	.a(FE_OFN137_n23948));
   in01f01 FE_OFC137_n23948 (.o(FE_OFN137_n23948),
	.a(n23948));
   in01f02 FE_OFC136_n23623 (.o(FE_OFN136_n23623),
	.a(FE_OFN135_n23623));
   in01f02 FE_OFC135_n23623 (.o(FE_OFN135_n23623),
	.a(n23623));
   in01f02 FE_OFC134_n23594 (.o(FE_OFN134_n23594),
	.a(FE_OFN133_n23594));
   in01f01 FE_OFC133_n23594 (.o(FE_OFN133_n23594),
	.a(n23594));
   in01f01 FE_OFC129_n23559 (.o(FE_OFN129_n23559),
	.a(n23559));
   in01f02 FE_OFC127_n23536 (.o(FE_OFN127_n23536),
	.a(n23536));
   in01f02 FE_OFC120_n23482 (.o(FE_OFN120_n23482),
	.a(FE_OFN119_n23482));
   in01f01 FE_OFC119_n23482 (.o(FE_OFN119_n23482),
	.a(n23482));
   in01f01 FE_OFC115_n23148 (.o(FE_OFN115_n23148),
	.a(n23148));
   in01f06 FE_OFC110_n22771 (.o(FE_OFN110_n22771),
	.a(FE_OFN109_n22771));
   in01f02 FE_OFC109_n22771 (.o(FE_OFN109_n22771),
	.a(n22771));
   in01f01 FE_OFC108_n22518 (.o(FE_OFN108_n22518),
	.a(FE_OFN107_n22518));
   in01f01 FE_OFC107_n22518 (.o(FE_OFN107_n22518),
	.a(n22518));
   in01f02 FE_OFC99_n21907 (.o(FE_OFN99_n21907),
	.a(n21907));
   in01f02 FE_OFC91_n21590 (.o(FE_OFN91_n21590),
	.a(FE_OFN90_n21590));
   in01f01 FE_OFC90_n21590 (.o(FE_OFN90_n21590),
	.a(n21590));
   in01f02 FE_OFC63_n19518 (.o(FE_OFN63_n19518),
	.a(FE_OFN62_n19518));
   in01f01 FE_OFC62_n19518 (.o(FE_OFN62_n19518),
	.a(n19518));
   in01f03 FE_OFC47_n19056 (.o(FE_OFN47_n19056),
	.a(FE_OFN46_n19056));
   in01f01 FE_OFC46_n19056 (.o(FE_OFN46_n19056),
	.a(n19056));
   in01f02 FE_OFC45_n19054 (.o(FE_OFN45_n19054),
	.a(FE_OFN43_n19054));
   in01f04 FE_OFC44_n19054 (.o(FE_OFN44_n19054),
	.a(FE_OFN43_n19054));
   in01f01 FE_OFC43_n19054 (.o(FE_OFN43_n19054),
	.a(n19054));
   in01f04 FE_OFC42_n19022 (.o(FE_OFN42_n19022),
	.a(FE_OFN41_n19022));
   in01f01 FE_OFC41_n19022 (.o(FE_OFN41_n19022),
	.a(n19022));
   in01f02 FE_OFC35_n19017 (.o(FE_OFN35_n19017),
	.a(FE_OFN34_n19017));
   in01f01 FE_OFC34_n19017 (.o(FE_OFN34_n19017),
	.a(n19017));
   in01f01 FE_OFC25_n17787 (.o(FE_OFN25_n17787),
	.a(FE_OFN24_n17787));
   in01f01 FE_OFC24_n17787 (.o(FE_OFN24_n17787),
	.a(n17787));
   in01f01 FE_OFC8_reset (.o(FE_OFN8_reset),
	.a(FE_OFN3_reset));
   in01f06 FE_OFC5_reset (.o(FE_OFN5_reset),
	.a(FE_OFN2_reset));
   in01f01 FE_OFC4_reset (.o(FE_OFN4_reset),
	.a(FE_OFN2_reset));
   in01f01 FE_OFC3_reset (.o(FE_OFN3_reset),
	.a(reset));
   in01f01 FE_OFC2_reset (.o(FE_OFN2_reset),
	.a(reset));
   in01f01 FE_OFC0_dataOut_N_40 (.o(FE_OFN1_dataOut_N_40),
	.a(FE_OFN0_dataOut_N_40));
   ms00f80 myChipID_f_reg_0_ (.o(myChipID_f_0_),
	.ck(clk),
	.d(N20));
   ms00f80 myChipID_f_reg_1_ (.o(myChipID_f_1_),
	.ck(clk),
	.d(N21));
   ms00f80 myChipID_f_reg_2_ (.o(myChipID_f_2_),
	.ck(clk),
	.d(N22));
   ms00f80 myChipID_f_reg_3_ (.o(myChipID_f_3_),
	.ck(clk),
	.d(N23));
   ms00f80 myChipID_f_reg_4_ (.o(myChipID_f_4_),
	.ck(clk),
	.d(N24));
   ms00f80 myChipID_f_reg_5_ (.o(myChipID_f_5_),
	.ck(clk),
	.d(N25));
   ms00f80 myChipID_f_reg_6_ (.o(myChipID_f_6_),
	.ck(clk),
	.d(N26));
   ms00f80 myChipID_f_reg_7_ (.o(myChipID_f_7_),
	.ck(clk),
	.d(N27));
   ms00f80 myChipID_f_reg_8_ (.o(myChipID_f_8_),
	.ck(clk),
	.d(N28));
   ms00f80 myChipID_f_reg_9_ (.o(myChipID_f_9_),
	.ck(clk),
	.d(N29));
   ms00f80 myChipID_f_reg_10_ (.o(myChipID_f_10_),
	.ck(clk),
	.d(N30));
   ms00f80 myChipID_f_reg_11_ (.o(myChipID_f_11_),
	.ck(clk),
	.d(N31));
   ms00f80 myChipID_f_reg_12_ (.o(myChipID_f_12_),
	.ck(clk),
	.d(N32));
   ms00f80 myChipID_f_reg_13_ (.o(myChipID_f_13_),
	.ck(clk),
	.d(N33));
   ms00f80 myLocX_f_reg_0_ (.o(myLocX_f_0_),
	.ck(clk),
	.d(N12));
   ms00f80 myLocX_f_reg_1_ (.o(myLocX_f_1_),
	.ck(clk),
	.d(N13));
   ms00f80 myLocX_f_reg_2_ (.o(myLocX_f_2_),
	.ck(clk),
	.d(N14));
   ms00f80 myLocX_f_reg_3_ (.o(myLocX_f_3_),
	.ck(clk),
	.d(N15));
   ms00f80 myLocX_f_reg_4_ (.o(myLocX_f_4_),
	.ck(clk),
	.d(N16));
   ms00f80 myLocX_f_reg_5_ (.o(myLocX_f_5_),
	.ck(clk),
	.d(N17));
   ms00f80 myLocX_f_reg_6_ (.o(myLocX_f_6_),
	.ck(clk),
	.d(N18));
   ms00f80 myLocX_f_reg_7_ (.o(myLocX_f_7_),
	.ck(clk),
	.d(N19));
   ms00f80 myLocY_f_reg_0_ (.o(myLocY_f_0_),
	.ck(clk),
	.d(N4));
   ms00f80 myLocY_f_reg_1_ (.o(myLocY_f_1_),
	.ck(clk),
	.d(N5));
   ms00f80 myLocY_f_reg_2_ (.o(myLocY_f_2_),
	.ck(clk),
	.d(N6));
   ms00f80 myLocY_f_reg_3_ (.o(myLocY_f_3_),
	.ck(clk),
	.d(N7));
   ms00f80 myLocY_f_reg_4_ (.o(myLocY_f_4_),
	.ck(clk),
	.d(N8));
   ms00f80 myLocY_f_reg_5_ (.o(myLocY_f_5_),
	.ck(clk),
	.d(N9));
   ms00f80 myLocY_f_reg_6_ (.o(myLocY_f_6_),
	.ck(clk),
	.d(N10));
   ms00f80 myLocY_f_reg_7_ (.o(myLocY_f_7_),
	.ck(clk),
	.d(N11));
   ms00f80 north_input_NIB_tail_ptr_f_reg_0_ (.o(north_input_NIB_tail_ptr_f_0_),
	.ck(clk),
	.d(n13388));
   ms00f80 north_input_NIB_tail_ptr_f_reg_1_ (.o(north_input_NIB_tail_ptr_f_1_),
	.ck(clk),
	.d(n13383));
   ms00f80 north_input_NIB_storage_data_f_reg_3__0_ (.o(north_input_NIB_storage_data_f_3__0_),
	.ck(clk),
	.d(n13378));
   ms00f80 north_input_NIB_storage_data_f_reg_3__1_ (.o(north_input_NIB_storage_data_f_3__1_),
	.ck(clk),
	.d(n13373));
   ms00f80 north_input_NIB_storage_data_f_reg_3__2_ (.o(north_input_NIB_storage_data_f_3__2_),
	.ck(clk),
	.d(n13368));
   ms00f80 north_input_NIB_storage_data_f_reg_3__3_ (.o(north_input_NIB_storage_data_f_3__3_),
	.ck(clk),
	.d(n13363));
   ms00f80 north_input_NIB_storage_data_f_reg_3__4_ (.o(north_input_NIB_storage_data_f_3__4_),
	.ck(clk),
	.d(n13358));
   ms00f80 north_input_NIB_storage_data_f_reg_3__5_ (.o(north_input_NIB_storage_data_f_3__5_),
	.ck(clk),
	.d(n13353));
   ms00f80 north_input_NIB_storage_data_f_reg_3__6_ (.o(north_input_NIB_storage_data_f_3__6_),
	.ck(clk),
	.d(n13348));
   ms00f80 north_input_NIB_storage_data_f_reg_3__7_ (.o(north_input_NIB_storage_data_f_3__7_),
	.ck(clk),
	.d(n13343));
   ms00f80 north_input_NIB_storage_data_f_reg_3__8_ (.o(north_input_NIB_storage_data_f_3__8_),
	.ck(clk),
	.d(n13338));
   ms00f80 north_input_NIB_storage_data_f_reg_3__9_ (.o(north_input_NIB_storage_data_f_3__9_),
	.ck(clk),
	.d(n13333));
   ms00f80 north_input_NIB_storage_data_f_reg_3__10_ (.o(north_input_NIB_storage_data_f_3__10_),
	.ck(clk),
	.d(n13328));
   ms00f80 north_input_NIB_storage_data_f_reg_3__11_ (.o(north_input_NIB_storage_data_f_3__11_),
	.ck(clk),
	.d(n13323));
   ms00f80 north_input_NIB_storage_data_f_reg_3__12_ (.o(north_input_NIB_storage_data_f_3__12_),
	.ck(clk),
	.d(n13318));
   ms00f80 north_input_NIB_storage_data_f_reg_3__13_ (.o(north_input_NIB_storage_data_f_3__13_),
	.ck(clk),
	.d(n13313));
   ms00f80 north_input_NIB_storage_data_f_reg_3__14_ (.o(north_input_NIB_storage_data_f_3__14_),
	.ck(clk),
	.d(n13308));
   ms00f80 north_input_NIB_storage_data_f_reg_3__15_ (.o(north_input_NIB_storage_data_f_3__15_),
	.ck(clk),
	.d(n13303));
   ms00f80 north_input_NIB_storage_data_f_reg_3__16_ (.o(north_input_NIB_storage_data_f_3__16_),
	.ck(clk),
	.d(n13298));
   ms00f80 north_input_NIB_storage_data_f_reg_3__17_ (.o(north_input_NIB_storage_data_f_3__17_),
	.ck(clk),
	.d(n13293));
   ms00f80 north_input_NIB_storage_data_f_reg_3__18_ (.o(north_input_NIB_storage_data_f_3__18_),
	.ck(clk),
	.d(n13288));
   ms00f80 north_input_NIB_storage_data_f_reg_3__19_ (.o(north_input_NIB_storage_data_f_3__19_),
	.ck(clk),
	.d(n13283));
   ms00f80 north_input_NIB_storage_data_f_reg_3__20_ (.o(north_input_NIB_storage_data_f_3__20_),
	.ck(clk),
	.d(n13278));
   ms00f80 north_input_NIB_storage_data_f_reg_3__21_ (.o(north_input_NIB_storage_data_f_3__21_),
	.ck(clk),
	.d(n13273));
   ms00f80 north_input_NIB_storage_data_f_reg_3__22_ (.o(north_input_NIB_storage_data_f_3__22_),
	.ck(clk),
	.d(n13268));
   ms00f80 north_input_NIB_storage_data_f_reg_3__23_ (.o(north_input_NIB_storage_data_f_3__23_),
	.ck(clk),
	.d(n13263));
   ms00f80 north_input_NIB_storage_data_f_reg_3__24_ (.o(north_input_NIB_storage_data_f_3__24_),
	.ck(clk),
	.d(n13258));
   ms00f80 north_input_NIB_storage_data_f_reg_3__25_ (.o(north_input_NIB_storage_data_f_3__25_),
	.ck(clk),
	.d(n13253));
   ms00f80 north_input_NIB_storage_data_f_reg_3__26_ (.o(north_input_NIB_storage_data_f_3__26_),
	.ck(clk),
	.d(n13248));
   ms00f80 north_input_NIB_storage_data_f_reg_3__27_ (.o(north_input_NIB_storage_data_f_3__27_),
	.ck(clk),
	.d(n13243));
   ms00f80 north_input_NIB_storage_data_f_reg_3__28_ (.o(north_input_NIB_storage_data_f_3__28_),
	.ck(clk),
	.d(n13238));
   ms00f80 north_input_NIB_storage_data_f_reg_3__29_ (.o(north_input_NIB_storage_data_f_3__29_),
	.ck(clk),
	.d(n13233));
   ms00f80 north_input_NIB_storage_data_f_reg_3__30_ (.o(north_input_NIB_storage_data_f_3__30_),
	.ck(clk),
	.d(n13228));
   ms00f80 north_input_NIB_storage_data_f_reg_3__31_ (.o(north_input_NIB_storage_data_f_3__31_),
	.ck(clk),
	.d(n13223));
   ms00f80 north_input_NIB_storage_data_f_reg_3__32_ (.o(north_input_NIB_storage_data_f_3__32_),
	.ck(clk),
	.d(n13218));
   ms00f80 north_input_NIB_storage_data_f_reg_3__33_ (.o(north_input_NIB_storage_data_f_3__33_),
	.ck(clk),
	.d(n13213));
   ms00f80 north_input_NIB_storage_data_f_reg_3__34_ (.o(north_input_NIB_storage_data_f_3__34_),
	.ck(clk),
	.d(n13208));
   ms00f80 north_input_NIB_storage_data_f_reg_3__35_ (.o(north_input_NIB_storage_data_f_3__35_),
	.ck(clk),
	.d(n13203));
   ms00f80 north_input_NIB_storage_data_f_reg_3__36_ (.o(north_input_NIB_storage_data_f_3__36_),
	.ck(clk),
	.d(n13198));
   ms00f80 north_input_NIB_storage_data_f_reg_3__37_ (.o(north_input_NIB_storage_data_f_3__37_),
	.ck(clk),
	.d(n13193));
   ms00f80 north_input_NIB_storage_data_f_reg_3__38_ (.o(north_input_NIB_storage_data_f_3__38_),
	.ck(clk),
	.d(n13188));
   ms00f80 north_input_NIB_storage_data_f_reg_3__39_ (.o(north_input_NIB_storage_data_f_3__39_),
	.ck(clk),
	.d(n13183));
   ms00f80 north_input_NIB_storage_data_f_reg_3__40_ (.o(north_input_NIB_storage_data_f_3__40_),
	.ck(clk),
	.d(n13178));
   ms00f80 north_input_NIB_storage_data_f_reg_3__41_ (.o(north_input_NIB_storage_data_f_3__41_),
	.ck(clk),
	.d(n13173));
   ms00f80 north_input_NIB_storage_data_f_reg_3__42_ (.o(north_input_NIB_storage_data_f_3__42_),
	.ck(clk),
	.d(n13168));
   ms00f80 north_input_NIB_storage_data_f_reg_3__43_ (.o(north_input_NIB_storage_data_f_3__43_),
	.ck(clk),
	.d(n13163));
   ms00f80 north_input_NIB_storage_data_f_reg_3__44_ (.o(north_input_NIB_storage_data_f_3__44_),
	.ck(clk),
	.d(n13158));
   ms00f80 north_input_NIB_storage_data_f_reg_3__45_ (.o(north_input_NIB_storage_data_f_3__45_),
	.ck(clk),
	.d(n13153));
   ms00f80 north_input_NIB_storage_data_f_reg_3__46_ (.o(north_input_NIB_storage_data_f_3__46_),
	.ck(clk),
	.d(n13148));
   ms00f80 north_input_NIB_storage_data_f_reg_3__47_ (.o(north_input_NIB_storage_data_f_3__47_),
	.ck(clk),
	.d(n13143));
   ms00f80 north_input_NIB_storage_data_f_reg_3__48_ (.o(north_input_NIB_storage_data_f_3__48_),
	.ck(clk),
	.d(n13138));
   ms00f80 north_input_NIB_storage_data_f_reg_3__49_ (.o(north_input_NIB_storage_data_f_3__49_),
	.ck(clk),
	.d(n13133));
   ms00f80 north_input_NIB_storage_data_f_reg_3__50_ (.o(north_input_NIB_storage_data_f_3__50_),
	.ck(clk),
	.d(n13128));
   ms00f80 north_input_NIB_storage_data_f_reg_3__51_ (.o(north_input_NIB_storage_data_f_3__51_),
	.ck(clk),
	.d(n13123));
   ms00f80 north_input_NIB_storage_data_f_reg_3__52_ (.o(north_input_NIB_storage_data_f_3__52_),
	.ck(clk),
	.d(n13118));
   ms00f80 north_input_NIB_storage_data_f_reg_3__53_ (.o(north_input_NIB_storage_data_f_3__53_),
	.ck(clk),
	.d(n13113));
   ms00f80 north_input_NIB_storage_data_f_reg_3__54_ (.o(north_input_NIB_storage_data_f_3__54_),
	.ck(clk),
	.d(n13108));
   ms00f80 north_input_NIB_storage_data_f_reg_3__55_ (.o(north_input_NIB_storage_data_f_3__55_),
	.ck(clk),
	.d(n13103));
   ms00f80 north_input_NIB_storage_data_f_reg_3__56_ (.o(north_input_NIB_storage_data_f_3__56_),
	.ck(clk),
	.d(n13098));
   ms00f80 north_input_NIB_storage_data_f_reg_3__57_ (.o(north_input_NIB_storage_data_f_3__57_),
	.ck(clk),
	.d(n13093));
   ms00f80 north_input_NIB_storage_data_f_reg_3__58_ (.o(north_input_NIB_storage_data_f_3__58_),
	.ck(clk),
	.d(n13088));
   ms00f80 north_input_NIB_storage_data_f_reg_3__59_ (.o(north_input_NIB_storage_data_f_3__59_),
	.ck(clk),
	.d(n13083));
   ms00f80 north_input_NIB_storage_data_f_reg_3__60_ (.o(north_input_NIB_storage_data_f_3__60_),
	.ck(clk),
	.d(n13078));
   ms00f80 north_input_NIB_storage_data_f_reg_3__61_ (.o(north_input_NIB_storage_data_f_3__61_),
	.ck(clk),
	.d(n13073));
   ms00f80 north_input_NIB_storage_data_f_reg_3__62_ (.o(north_input_NIB_storage_data_f_3__62_),
	.ck(clk),
	.d(n13068));
   ms00f80 north_input_NIB_storage_data_f_reg_3__63_ (.o(north_input_NIB_storage_data_f_3__63_),
	.ck(clk),
	.d(n13063));
   ms00f80 north_input_NIB_storage_data_f_reg_2__0_ (.o(north_input_NIB_storage_data_f_2__0_),
	.ck(clk),
	.d(n13058));
   ms00f80 north_input_NIB_storage_data_f_reg_2__1_ (.o(north_input_NIB_storage_data_f_2__1_),
	.ck(clk),
	.d(n13053));
   ms00f80 north_input_NIB_storage_data_f_reg_2__2_ (.o(north_input_NIB_storage_data_f_2__2_),
	.ck(clk),
	.d(n13048));
   ms00f80 north_input_NIB_storage_data_f_reg_2__3_ (.o(north_input_NIB_storage_data_f_2__3_),
	.ck(clk),
	.d(n13043));
   ms00f80 north_input_NIB_storage_data_f_reg_2__4_ (.o(north_input_NIB_storage_data_f_2__4_),
	.ck(clk),
	.d(n13038));
   ms00f80 north_input_NIB_storage_data_f_reg_2__5_ (.o(north_input_NIB_storage_data_f_2__5_),
	.ck(clk),
	.d(n13033));
   ms00f80 north_input_NIB_storage_data_f_reg_2__6_ (.o(north_input_NIB_storage_data_f_2__6_),
	.ck(clk),
	.d(n13028));
   ms00f80 north_input_NIB_storage_data_f_reg_2__7_ (.o(north_input_NIB_storage_data_f_2__7_),
	.ck(clk),
	.d(n13023));
   ms00f80 north_input_NIB_storage_data_f_reg_2__8_ (.o(north_input_NIB_storage_data_f_2__8_),
	.ck(clk),
	.d(n13018));
   ms00f80 north_input_NIB_storage_data_f_reg_2__9_ (.o(north_input_NIB_storage_data_f_2__9_),
	.ck(clk),
	.d(n13013));
   ms00f80 north_input_NIB_storage_data_f_reg_2__10_ (.o(north_input_NIB_storage_data_f_2__10_),
	.ck(clk),
	.d(n13008));
   ms00f80 north_input_NIB_storage_data_f_reg_2__11_ (.o(north_input_NIB_storage_data_f_2__11_),
	.ck(clk),
	.d(n13003));
   ms00f80 north_input_NIB_storage_data_f_reg_2__12_ (.o(north_input_NIB_storage_data_f_2__12_),
	.ck(clk),
	.d(n12998));
   ms00f80 north_input_NIB_storage_data_f_reg_2__13_ (.o(north_input_NIB_storage_data_f_2__13_),
	.ck(clk),
	.d(n12993));
   ms00f80 north_input_NIB_storage_data_f_reg_2__14_ (.o(north_input_NIB_storage_data_f_2__14_),
	.ck(clk),
	.d(n12988));
   ms00f80 north_input_NIB_storage_data_f_reg_2__15_ (.o(north_input_NIB_storage_data_f_2__15_),
	.ck(clk),
	.d(n12983));
   ms00f80 north_input_NIB_storage_data_f_reg_2__16_ (.o(north_input_NIB_storage_data_f_2__16_),
	.ck(clk),
	.d(n12978));
   ms00f80 north_input_NIB_storage_data_f_reg_2__17_ (.o(north_input_NIB_storage_data_f_2__17_),
	.ck(clk),
	.d(n12973));
   ms00f80 north_input_NIB_storage_data_f_reg_2__18_ (.o(north_input_NIB_storage_data_f_2__18_),
	.ck(clk),
	.d(n12968));
   ms00f80 north_input_NIB_storage_data_f_reg_2__19_ (.o(north_input_NIB_storage_data_f_2__19_),
	.ck(clk),
	.d(n12963));
   ms00f80 north_input_NIB_storage_data_f_reg_2__20_ (.o(north_input_NIB_storage_data_f_2__20_),
	.ck(clk),
	.d(n12958));
   ms00f80 north_input_NIB_storage_data_f_reg_2__21_ (.o(north_input_NIB_storage_data_f_2__21_),
	.ck(clk),
	.d(n12953));
   ms00f80 north_input_NIB_storage_data_f_reg_2__22_ (.o(north_input_NIB_storage_data_f_2__22_),
	.ck(clk),
	.d(n12948));
   ms00f80 north_input_NIB_storage_data_f_reg_2__23_ (.o(north_input_NIB_storage_data_f_2__23_),
	.ck(clk),
	.d(n12943));
   ms00f80 north_input_NIB_storage_data_f_reg_2__24_ (.o(north_input_NIB_storage_data_f_2__24_),
	.ck(clk),
	.d(n12938));
   ms00f80 north_input_NIB_storage_data_f_reg_2__25_ (.o(north_input_NIB_storage_data_f_2__25_),
	.ck(clk),
	.d(n12933));
   ms00f80 north_input_NIB_storage_data_f_reg_2__26_ (.o(north_input_NIB_storage_data_f_2__26_),
	.ck(clk),
	.d(n12928));
   ms00f80 north_input_NIB_storage_data_f_reg_2__27_ (.o(north_input_NIB_storage_data_f_2__27_),
	.ck(clk),
	.d(n12923));
   ms00f80 north_input_NIB_storage_data_f_reg_2__28_ (.o(north_input_NIB_storage_data_f_2__28_),
	.ck(clk),
	.d(n12918));
   ms00f80 north_input_NIB_storage_data_f_reg_2__29_ (.o(north_input_NIB_storage_data_f_2__29_),
	.ck(clk),
	.d(n12913));
   ms00f80 north_input_NIB_storage_data_f_reg_2__30_ (.o(north_input_NIB_storage_data_f_2__30_),
	.ck(clk),
	.d(n12908));
   ms00f80 north_input_NIB_storage_data_f_reg_2__31_ (.o(north_input_NIB_storage_data_f_2__31_),
	.ck(clk),
	.d(n12903));
   ms00f80 north_input_NIB_storage_data_f_reg_2__32_ (.o(north_input_NIB_storage_data_f_2__32_),
	.ck(clk),
	.d(n12898));
   ms00f80 north_input_NIB_storage_data_f_reg_2__33_ (.o(north_input_NIB_storage_data_f_2__33_),
	.ck(clk),
	.d(n12893));
   ms00f80 north_input_NIB_storage_data_f_reg_2__34_ (.o(north_input_NIB_storage_data_f_2__34_),
	.ck(clk),
	.d(n12888));
   ms00f80 north_input_NIB_storage_data_f_reg_2__35_ (.o(north_input_NIB_storage_data_f_2__35_),
	.ck(clk),
	.d(n12883));
   ms00f80 north_input_NIB_storage_data_f_reg_2__36_ (.o(north_input_NIB_storage_data_f_2__36_),
	.ck(clk),
	.d(n12878));
   ms00f80 north_input_NIB_storage_data_f_reg_2__37_ (.o(north_input_NIB_storage_data_f_2__37_),
	.ck(clk),
	.d(n12873));
   ms00f80 north_input_NIB_storage_data_f_reg_2__38_ (.o(north_input_NIB_storage_data_f_2__38_),
	.ck(clk),
	.d(n12868));
   ms00f80 north_input_NIB_storage_data_f_reg_2__39_ (.o(north_input_NIB_storage_data_f_2__39_),
	.ck(clk),
	.d(n12863));
   ms00f80 north_input_NIB_storage_data_f_reg_2__40_ (.o(north_input_NIB_storage_data_f_2__40_),
	.ck(clk),
	.d(n12858));
   ms00f80 north_input_NIB_storage_data_f_reg_2__41_ (.o(north_input_NIB_storage_data_f_2__41_),
	.ck(clk),
	.d(n12853));
   ms00f80 north_input_NIB_storage_data_f_reg_2__42_ (.o(north_input_NIB_storage_data_f_2__42_),
	.ck(clk),
	.d(n12848));
   ms00f80 north_input_NIB_storage_data_f_reg_2__43_ (.o(north_input_NIB_storage_data_f_2__43_),
	.ck(clk),
	.d(n12843));
   ms00f80 north_input_NIB_storage_data_f_reg_2__44_ (.o(north_input_NIB_storage_data_f_2__44_),
	.ck(clk),
	.d(n12838));
   ms00f80 north_input_NIB_storage_data_f_reg_2__45_ (.o(north_input_NIB_storage_data_f_2__45_),
	.ck(clk),
	.d(n12833));
   ms00f80 north_input_NIB_storage_data_f_reg_2__46_ (.o(north_input_NIB_storage_data_f_2__46_),
	.ck(clk),
	.d(n12828));
   ms00f80 north_input_NIB_storage_data_f_reg_2__47_ (.o(north_input_NIB_storage_data_f_2__47_),
	.ck(clk),
	.d(n12823));
   ms00f80 north_input_NIB_storage_data_f_reg_2__48_ (.o(north_input_NIB_storage_data_f_2__48_),
	.ck(clk),
	.d(n12818));
   ms00f80 north_input_NIB_storage_data_f_reg_2__49_ (.o(north_input_NIB_storage_data_f_2__49_),
	.ck(clk),
	.d(n12813));
   ms00f80 north_input_NIB_storage_data_f_reg_2__50_ (.o(north_input_NIB_storage_data_f_2__50_),
	.ck(clk),
	.d(n12808));
   ms00f80 north_input_NIB_storage_data_f_reg_2__51_ (.o(north_input_NIB_storage_data_f_2__51_),
	.ck(clk),
	.d(n12803));
   ms00f80 north_input_NIB_storage_data_f_reg_2__52_ (.o(north_input_NIB_storage_data_f_2__52_),
	.ck(clk),
	.d(n12798));
   ms00f80 north_input_NIB_storage_data_f_reg_2__53_ (.o(north_input_NIB_storage_data_f_2__53_),
	.ck(clk),
	.d(n12793));
   ms00f80 north_input_NIB_storage_data_f_reg_2__54_ (.o(north_input_NIB_storage_data_f_2__54_),
	.ck(clk),
	.d(n12788));
   ms00f80 north_input_NIB_storage_data_f_reg_2__55_ (.o(north_input_NIB_storage_data_f_2__55_),
	.ck(clk),
	.d(n12783));
   ms00f80 north_input_NIB_storage_data_f_reg_2__56_ (.o(north_input_NIB_storage_data_f_2__56_),
	.ck(clk),
	.d(n12778));
   ms00f80 north_input_NIB_storage_data_f_reg_2__57_ (.o(north_input_NIB_storage_data_f_2__57_),
	.ck(clk),
	.d(n12773));
   ms00f80 north_input_NIB_storage_data_f_reg_2__58_ (.o(north_input_NIB_storage_data_f_2__58_),
	.ck(clk),
	.d(n12768));
   ms00f80 north_input_NIB_storage_data_f_reg_2__59_ (.o(north_input_NIB_storage_data_f_2__59_),
	.ck(clk),
	.d(n12763));
   ms00f80 north_input_NIB_storage_data_f_reg_2__60_ (.o(north_input_NIB_storage_data_f_2__60_),
	.ck(clk),
	.d(n12758));
   ms00f80 north_input_NIB_storage_data_f_reg_2__61_ (.o(north_input_NIB_storage_data_f_2__61_),
	.ck(clk),
	.d(n12753));
   ms00f80 north_input_NIB_storage_data_f_reg_2__62_ (.o(north_input_NIB_storage_data_f_2__62_),
	.ck(clk),
	.d(n12748));
   ms00f80 north_input_NIB_storage_data_f_reg_2__63_ (.o(north_input_NIB_storage_data_f_2__63_),
	.ck(clk),
	.d(n12743));
   ms00f80 north_input_NIB_storage_data_f_reg_1__0_ (.o(north_input_NIB_storage_data_f_1__0_),
	.ck(clk),
	.d(n12738));
   ms00f80 north_input_NIB_storage_data_f_reg_1__1_ (.o(north_input_NIB_storage_data_f_1__1_),
	.ck(clk),
	.d(n12733));
   ms00f80 north_input_NIB_storage_data_f_reg_1__2_ (.o(north_input_NIB_storage_data_f_1__2_),
	.ck(clk),
	.d(n12728));
   ms00f80 north_input_NIB_storage_data_f_reg_1__3_ (.o(north_input_NIB_storage_data_f_1__3_),
	.ck(clk),
	.d(n12723));
   ms00f80 north_input_NIB_storage_data_f_reg_1__4_ (.o(north_input_NIB_storage_data_f_1__4_),
	.ck(clk),
	.d(n12718));
   ms00f80 north_input_NIB_storage_data_f_reg_1__5_ (.o(north_input_NIB_storage_data_f_1__5_),
	.ck(clk),
	.d(n12713));
   ms00f80 north_input_NIB_storage_data_f_reg_1__6_ (.o(north_input_NIB_storage_data_f_1__6_),
	.ck(clk),
	.d(n12708));
   ms00f80 north_input_NIB_storage_data_f_reg_1__7_ (.o(north_input_NIB_storage_data_f_1__7_),
	.ck(clk),
	.d(n12703));
   ms00f80 north_input_NIB_storage_data_f_reg_1__8_ (.o(north_input_NIB_storage_data_f_1__8_),
	.ck(clk),
	.d(n12698));
   ms00f80 north_input_NIB_storage_data_f_reg_1__9_ (.o(north_input_NIB_storage_data_f_1__9_),
	.ck(clk),
	.d(n12693));
   ms00f80 north_input_NIB_storage_data_f_reg_1__10_ (.o(north_input_NIB_storage_data_f_1__10_),
	.ck(clk),
	.d(n12688));
   ms00f80 north_input_NIB_storage_data_f_reg_1__11_ (.o(north_input_NIB_storage_data_f_1__11_),
	.ck(clk),
	.d(n12683));
   ms00f80 north_input_NIB_storage_data_f_reg_1__12_ (.o(north_input_NIB_storage_data_f_1__12_),
	.ck(clk),
	.d(n12678));
   ms00f80 north_input_NIB_storage_data_f_reg_1__13_ (.o(north_input_NIB_storage_data_f_1__13_),
	.ck(clk),
	.d(n12673));
   ms00f80 north_input_NIB_storage_data_f_reg_1__14_ (.o(north_input_NIB_storage_data_f_1__14_),
	.ck(clk),
	.d(n12668));
   ms00f80 north_input_NIB_storage_data_f_reg_1__15_ (.o(north_input_NIB_storage_data_f_1__15_),
	.ck(clk),
	.d(n12663));
   ms00f80 north_input_NIB_storage_data_f_reg_1__16_ (.o(north_input_NIB_storage_data_f_1__16_),
	.ck(clk),
	.d(n12658));
   ms00f80 north_input_NIB_storage_data_f_reg_1__17_ (.o(north_input_NIB_storage_data_f_1__17_),
	.ck(clk),
	.d(n12653));
   ms00f80 north_input_NIB_storage_data_f_reg_1__18_ (.o(north_input_NIB_storage_data_f_1__18_),
	.ck(clk),
	.d(n12648));
   ms00f80 north_input_NIB_storage_data_f_reg_1__19_ (.o(north_input_NIB_storage_data_f_1__19_),
	.ck(clk),
	.d(n12643));
   ms00f80 north_input_NIB_storage_data_f_reg_1__20_ (.o(north_input_NIB_storage_data_f_1__20_),
	.ck(clk),
	.d(n12638));
   ms00f80 north_input_NIB_storage_data_f_reg_1__21_ (.o(north_input_NIB_storage_data_f_1__21_),
	.ck(clk),
	.d(n12633));
   ms00f80 north_input_NIB_storage_data_f_reg_1__22_ (.o(north_input_NIB_storage_data_f_1__22_),
	.ck(clk),
	.d(n12628));
   ms00f80 north_input_NIB_storage_data_f_reg_1__23_ (.o(north_input_NIB_storage_data_f_1__23_),
	.ck(clk),
	.d(n12623));
   ms00f80 north_input_NIB_storage_data_f_reg_1__24_ (.o(north_input_NIB_storage_data_f_1__24_),
	.ck(clk),
	.d(n12618));
   ms00f80 north_input_NIB_storage_data_f_reg_1__25_ (.o(north_input_NIB_storage_data_f_1__25_),
	.ck(clk),
	.d(n12613));
   ms00f80 north_input_NIB_storage_data_f_reg_1__26_ (.o(north_input_NIB_storage_data_f_1__26_),
	.ck(clk),
	.d(n12608));
   ms00f80 north_input_NIB_storage_data_f_reg_1__27_ (.o(north_input_NIB_storage_data_f_1__27_),
	.ck(clk),
	.d(n12603));
   ms00f80 north_input_NIB_storage_data_f_reg_1__28_ (.o(north_input_NIB_storage_data_f_1__28_),
	.ck(clk),
	.d(n12598));
   ms00f80 north_input_NIB_storage_data_f_reg_1__29_ (.o(north_input_NIB_storage_data_f_1__29_),
	.ck(clk),
	.d(n12593));
   ms00f80 north_input_NIB_storage_data_f_reg_1__30_ (.o(north_input_NIB_storage_data_f_1__30_),
	.ck(clk),
	.d(n12588));
   ms00f80 north_input_NIB_storage_data_f_reg_1__31_ (.o(north_input_NIB_storage_data_f_1__31_),
	.ck(clk),
	.d(n12583));
   ms00f80 north_input_NIB_storage_data_f_reg_1__32_ (.o(north_input_NIB_storage_data_f_1__32_),
	.ck(clk),
	.d(n12578));
   ms00f80 north_input_NIB_storage_data_f_reg_1__33_ (.o(north_input_NIB_storage_data_f_1__33_),
	.ck(clk),
	.d(n12573));
   ms00f80 north_input_NIB_storage_data_f_reg_1__34_ (.o(north_input_NIB_storage_data_f_1__34_),
	.ck(clk),
	.d(n12568));
   ms00f80 north_input_NIB_storage_data_f_reg_1__35_ (.o(north_input_NIB_storage_data_f_1__35_),
	.ck(clk),
	.d(n12563));
   ms00f80 north_input_NIB_storage_data_f_reg_1__36_ (.o(north_input_NIB_storage_data_f_1__36_),
	.ck(clk),
	.d(n12558));
   ms00f80 north_input_NIB_storage_data_f_reg_1__37_ (.o(north_input_NIB_storage_data_f_1__37_),
	.ck(clk),
	.d(n12553));
   ms00f80 north_input_NIB_storage_data_f_reg_1__38_ (.o(north_input_NIB_storage_data_f_1__38_),
	.ck(clk),
	.d(n12548));
   ms00f80 north_input_NIB_storage_data_f_reg_1__39_ (.o(north_input_NIB_storage_data_f_1__39_),
	.ck(clk),
	.d(n12543));
   ms00f80 north_input_NIB_storage_data_f_reg_1__40_ (.o(north_input_NIB_storage_data_f_1__40_),
	.ck(clk),
	.d(n12538));
   ms00f80 north_input_NIB_storage_data_f_reg_1__41_ (.o(north_input_NIB_storage_data_f_1__41_),
	.ck(clk),
	.d(n12533));
   ms00f80 north_input_NIB_storage_data_f_reg_1__42_ (.o(north_input_NIB_storage_data_f_1__42_),
	.ck(clk),
	.d(n12528));
   ms00f80 north_input_NIB_storage_data_f_reg_1__43_ (.o(north_input_NIB_storage_data_f_1__43_),
	.ck(clk),
	.d(n12523));
   ms00f80 north_input_NIB_storage_data_f_reg_1__44_ (.o(north_input_NIB_storage_data_f_1__44_),
	.ck(clk),
	.d(n12518));
   ms00f80 north_input_NIB_storage_data_f_reg_1__45_ (.o(north_input_NIB_storage_data_f_1__45_),
	.ck(clk),
	.d(n12513));
   ms00f80 north_input_NIB_storage_data_f_reg_1__46_ (.o(north_input_NIB_storage_data_f_1__46_),
	.ck(clk),
	.d(n12508));
   ms00f80 north_input_NIB_storage_data_f_reg_1__47_ (.o(north_input_NIB_storage_data_f_1__47_),
	.ck(clk),
	.d(n12503));
   ms00f80 north_input_NIB_storage_data_f_reg_1__48_ (.o(north_input_NIB_storage_data_f_1__48_),
	.ck(clk),
	.d(n12498));
   ms00f80 north_input_NIB_storage_data_f_reg_1__49_ (.o(north_input_NIB_storage_data_f_1__49_),
	.ck(clk),
	.d(n12493));
   ms00f80 north_input_NIB_storage_data_f_reg_1__50_ (.o(north_input_NIB_storage_data_f_1__50_),
	.ck(clk),
	.d(n12488));
   ms00f80 north_input_NIB_storage_data_f_reg_1__51_ (.o(north_input_NIB_storage_data_f_1__51_),
	.ck(clk),
	.d(n12483));
   ms00f80 north_input_NIB_storage_data_f_reg_1__52_ (.o(north_input_NIB_storage_data_f_1__52_),
	.ck(clk),
	.d(n12478));
   ms00f80 north_input_NIB_storage_data_f_reg_1__53_ (.o(north_input_NIB_storage_data_f_1__53_),
	.ck(clk),
	.d(n12473));
   ms00f80 north_input_NIB_storage_data_f_reg_1__54_ (.o(north_input_NIB_storage_data_f_1__54_),
	.ck(clk),
	.d(n12468));
   ms00f80 north_input_NIB_storage_data_f_reg_1__55_ (.o(north_input_NIB_storage_data_f_1__55_),
	.ck(clk),
	.d(n12463));
   ms00f80 north_input_NIB_storage_data_f_reg_1__56_ (.o(north_input_NIB_storage_data_f_1__56_),
	.ck(clk),
	.d(n12458));
   ms00f80 north_input_NIB_storage_data_f_reg_1__57_ (.o(north_input_NIB_storage_data_f_1__57_),
	.ck(clk),
	.d(n12453));
   ms00f80 north_input_NIB_storage_data_f_reg_1__58_ (.o(north_input_NIB_storage_data_f_1__58_),
	.ck(clk),
	.d(n12448));
   ms00f80 north_input_NIB_storage_data_f_reg_1__59_ (.o(north_input_NIB_storage_data_f_1__59_),
	.ck(clk),
	.d(n12443));
   ms00f80 north_input_NIB_storage_data_f_reg_1__60_ (.o(north_input_NIB_storage_data_f_1__60_),
	.ck(clk),
	.d(n12438));
   ms00f80 north_input_NIB_storage_data_f_reg_1__61_ (.o(north_input_NIB_storage_data_f_1__61_),
	.ck(clk),
	.d(n12433));
   ms00f80 north_input_NIB_storage_data_f_reg_1__62_ (.o(north_input_NIB_storage_data_f_1__62_),
	.ck(clk),
	.d(n12428));
   ms00f80 north_input_NIB_storage_data_f_reg_1__63_ (.o(north_input_NIB_storage_data_f_1__63_),
	.ck(clk),
	.d(n12423));
   ms00f80 north_input_NIB_storage_data_f_reg_0__0_ (.o(north_input_NIB_storage_data_f_0__0_),
	.ck(clk),
	.d(n12418));
   ms00f80 north_input_NIB_storage_data_f_reg_0__1_ (.o(north_input_NIB_storage_data_f_0__1_),
	.ck(clk),
	.d(n12413));
   ms00f80 north_input_NIB_storage_data_f_reg_0__2_ (.o(north_input_NIB_storage_data_f_0__2_),
	.ck(clk),
	.d(n12408));
   ms00f80 north_input_NIB_storage_data_f_reg_0__3_ (.o(north_input_NIB_storage_data_f_0__3_),
	.ck(clk),
	.d(n12403));
   ms00f80 north_input_NIB_storage_data_f_reg_0__4_ (.o(north_input_NIB_storage_data_f_0__4_),
	.ck(clk),
	.d(n12398));
   ms00f80 north_input_NIB_storage_data_f_reg_0__5_ (.o(north_input_NIB_storage_data_f_0__5_),
	.ck(clk),
	.d(n12393));
   ms00f80 north_input_NIB_storage_data_f_reg_0__6_ (.o(north_input_NIB_storage_data_f_0__6_),
	.ck(clk),
	.d(n12388));
   ms00f80 north_input_NIB_storage_data_f_reg_0__7_ (.o(north_input_NIB_storage_data_f_0__7_),
	.ck(clk),
	.d(n12383));
   ms00f80 north_input_NIB_storage_data_f_reg_0__8_ (.o(north_input_NIB_storage_data_f_0__8_),
	.ck(clk),
	.d(n12378));
   ms00f80 north_input_NIB_storage_data_f_reg_0__9_ (.o(north_input_NIB_storage_data_f_0__9_),
	.ck(clk),
	.d(n12373));
   ms00f80 north_input_NIB_storage_data_f_reg_0__10_ (.o(north_input_NIB_storage_data_f_0__10_),
	.ck(clk),
	.d(n12368));
   ms00f80 north_input_NIB_storage_data_f_reg_0__11_ (.o(north_input_NIB_storage_data_f_0__11_),
	.ck(clk),
	.d(n12363));
   ms00f80 north_input_NIB_storage_data_f_reg_0__12_ (.o(north_input_NIB_storage_data_f_0__12_),
	.ck(clk),
	.d(n12358));
   ms00f80 north_input_NIB_storage_data_f_reg_0__13_ (.o(north_input_NIB_storage_data_f_0__13_),
	.ck(clk),
	.d(n12353));
   ms00f80 north_input_NIB_storage_data_f_reg_0__14_ (.o(north_input_NIB_storage_data_f_0__14_),
	.ck(clk),
	.d(n12348));
   ms00f80 north_input_NIB_storage_data_f_reg_0__15_ (.o(north_input_NIB_storage_data_f_0__15_),
	.ck(clk),
	.d(n12343));
   ms00f80 north_input_NIB_storage_data_f_reg_0__16_ (.o(north_input_NIB_storage_data_f_0__16_),
	.ck(clk),
	.d(n12338));
   ms00f80 north_input_NIB_storage_data_f_reg_0__17_ (.o(north_input_NIB_storage_data_f_0__17_),
	.ck(clk),
	.d(n12333));
   ms00f80 north_input_NIB_storage_data_f_reg_0__18_ (.o(north_input_NIB_storage_data_f_0__18_),
	.ck(clk),
	.d(n12328));
   ms00f80 north_input_NIB_storage_data_f_reg_0__19_ (.o(north_input_NIB_storage_data_f_0__19_),
	.ck(clk),
	.d(n12323));
   ms00f80 north_input_NIB_storage_data_f_reg_0__20_ (.o(north_input_NIB_storage_data_f_0__20_),
	.ck(clk),
	.d(n12318));
   ms00f80 north_input_NIB_storage_data_f_reg_0__21_ (.o(north_input_NIB_storage_data_f_0__21_),
	.ck(clk),
	.d(n12313));
   ms00f80 north_input_NIB_storage_data_f_reg_0__22_ (.o(north_input_NIB_storage_data_f_0__22_),
	.ck(clk),
	.d(n12308));
   ms00f80 north_input_NIB_storage_data_f_reg_0__23_ (.o(north_input_NIB_storage_data_f_0__23_),
	.ck(clk),
	.d(n12303));
   ms00f80 north_input_NIB_storage_data_f_reg_0__24_ (.o(north_input_NIB_storage_data_f_0__24_),
	.ck(clk),
	.d(n12298));
   ms00f80 north_input_NIB_storage_data_f_reg_0__25_ (.o(north_input_NIB_storage_data_f_0__25_),
	.ck(clk),
	.d(n12293));
   ms00f80 north_input_NIB_storage_data_f_reg_0__26_ (.o(north_input_NIB_storage_data_f_0__26_),
	.ck(clk),
	.d(n12288));
   ms00f80 north_input_NIB_storage_data_f_reg_0__27_ (.o(north_input_NIB_storage_data_f_0__27_),
	.ck(clk),
	.d(n12283));
   ms00f80 north_input_NIB_storage_data_f_reg_0__28_ (.o(north_input_NIB_storage_data_f_0__28_),
	.ck(clk),
	.d(n12278));
   ms00f80 north_input_NIB_storage_data_f_reg_0__29_ (.o(north_input_NIB_storage_data_f_0__29_),
	.ck(clk),
	.d(n12273));
   ms00f80 north_input_NIB_storage_data_f_reg_0__30_ (.o(north_input_NIB_storage_data_f_0__30_),
	.ck(clk),
	.d(n12268));
   ms00f80 north_input_NIB_storage_data_f_reg_0__31_ (.o(north_input_NIB_storage_data_f_0__31_),
	.ck(clk),
	.d(n12263));
   ms00f80 north_input_NIB_storage_data_f_reg_0__32_ (.o(north_input_NIB_storage_data_f_0__32_),
	.ck(clk),
	.d(n12258));
   ms00f80 north_input_NIB_storage_data_f_reg_0__33_ (.o(north_input_NIB_storage_data_f_0__33_),
	.ck(clk),
	.d(n12253));
   ms00f80 north_input_NIB_storage_data_f_reg_0__34_ (.o(north_input_NIB_storage_data_f_0__34_),
	.ck(clk),
	.d(n12248));
   ms00f80 north_input_NIB_storage_data_f_reg_0__35_ (.o(north_input_NIB_storage_data_f_0__35_),
	.ck(clk),
	.d(n12243));
   ms00f80 north_input_NIB_storage_data_f_reg_0__36_ (.o(north_input_NIB_storage_data_f_0__36_),
	.ck(clk),
	.d(n12238));
   ms00f80 north_input_NIB_storage_data_f_reg_0__37_ (.o(north_input_NIB_storage_data_f_0__37_),
	.ck(clk),
	.d(n12233));
   ms00f80 north_input_NIB_storage_data_f_reg_0__38_ (.o(north_input_NIB_storage_data_f_0__38_),
	.ck(clk),
	.d(n12228));
   ms00f80 north_input_NIB_storage_data_f_reg_0__39_ (.o(north_input_NIB_storage_data_f_0__39_),
	.ck(clk),
	.d(n12223));
   ms00f80 north_input_NIB_storage_data_f_reg_0__40_ (.o(north_input_NIB_storage_data_f_0__40_),
	.ck(clk),
	.d(n12218));
   ms00f80 north_input_NIB_storage_data_f_reg_0__41_ (.o(north_input_NIB_storage_data_f_0__41_),
	.ck(clk),
	.d(n12213));
   ms00f80 north_input_NIB_storage_data_f_reg_0__42_ (.o(north_input_NIB_storage_data_f_0__42_),
	.ck(clk),
	.d(n12208));
   ms00f80 north_input_NIB_storage_data_f_reg_0__43_ (.o(north_input_NIB_storage_data_f_0__43_),
	.ck(clk),
	.d(n12203));
   ms00f80 north_input_NIB_storage_data_f_reg_0__44_ (.o(north_input_NIB_storage_data_f_0__44_),
	.ck(clk),
	.d(n12198));
   ms00f80 north_input_NIB_storage_data_f_reg_0__45_ (.o(north_input_NIB_storage_data_f_0__45_),
	.ck(clk),
	.d(n12193));
   ms00f80 north_input_NIB_storage_data_f_reg_0__46_ (.o(north_input_NIB_storage_data_f_0__46_),
	.ck(clk),
	.d(n12188));
   ms00f80 north_input_NIB_storage_data_f_reg_0__47_ (.o(north_input_NIB_storage_data_f_0__47_),
	.ck(clk),
	.d(n12183));
   ms00f80 north_input_NIB_storage_data_f_reg_0__48_ (.o(north_input_NIB_storage_data_f_0__48_),
	.ck(clk),
	.d(n12178));
   ms00f80 north_input_NIB_storage_data_f_reg_0__49_ (.o(north_input_NIB_storage_data_f_0__49_),
	.ck(clk),
	.d(n12173));
   ms00f80 north_input_NIB_storage_data_f_reg_0__50_ (.o(north_input_NIB_storage_data_f_0__50_),
	.ck(clk),
	.d(n12168));
   ms00f80 north_input_NIB_storage_data_f_reg_0__51_ (.o(north_input_NIB_storage_data_f_0__51_),
	.ck(clk),
	.d(n12163));
   ms00f80 north_input_NIB_storage_data_f_reg_0__52_ (.o(north_input_NIB_storage_data_f_0__52_),
	.ck(clk),
	.d(n12158));
   ms00f80 north_input_NIB_storage_data_f_reg_0__53_ (.o(north_input_NIB_storage_data_f_0__53_),
	.ck(clk),
	.d(n12153));
   ms00f80 north_input_NIB_storage_data_f_reg_0__54_ (.o(north_input_NIB_storage_data_f_0__54_),
	.ck(clk),
	.d(n12148));
   ms00f80 north_input_NIB_storage_data_f_reg_0__55_ (.o(north_input_NIB_storage_data_f_0__55_),
	.ck(clk),
	.d(n12143));
   ms00f80 north_input_NIB_storage_data_f_reg_0__56_ (.o(north_input_NIB_storage_data_f_0__56_),
	.ck(clk),
	.d(n12138));
   ms00f80 north_input_NIB_storage_data_f_reg_0__57_ (.o(north_input_NIB_storage_data_f_0__57_),
	.ck(clk),
	.d(n12133));
   ms00f80 north_input_NIB_storage_data_f_reg_0__58_ (.o(north_input_NIB_storage_data_f_0__58_),
	.ck(clk),
	.d(n12128));
   ms00f80 north_input_NIB_storage_data_f_reg_0__59_ (.o(north_input_NIB_storage_data_f_0__59_),
	.ck(clk),
	.d(n12123));
   ms00f80 north_input_NIB_storage_data_f_reg_0__60_ (.o(north_input_NIB_storage_data_f_0__60_),
	.ck(clk),
	.d(n12118));
   ms00f80 north_input_NIB_storage_data_f_reg_0__61_ (.o(north_input_NIB_storage_data_f_0__61_),
	.ck(clk),
	.d(n12113));
   ms00f80 north_input_NIB_storage_data_f_reg_0__62_ (.o(north_input_NIB_storage_data_f_0__62_),
	.ck(clk),
	.d(n12108));
   ms00f80 north_input_NIB_storage_data_f_reg_0__63_ (.o(north_input_NIB_storage_data_f_0__63_),
	.ck(clk),
	.d(n12103));
   ms00f80 east_input_NIB_tail_ptr_f_reg_0_ (.o(east_input_NIB_tail_ptr_f_0_),
	.ck(clk),
	.d(n12098));
   ms00f80 east_input_NIB_tail_ptr_f_reg_1_ (.o(east_input_NIB_tail_ptr_f_1_),
	.ck(clk),
	.d(n12093));
   ms00f80 east_input_NIB_storage_data_f_reg_3__0_ (.o(east_input_NIB_storage_data_f_3__0_),
	.ck(clk),
	.d(n12088));
   ms00f80 east_input_NIB_storage_data_f_reg_3__1_ (.o(east_input_NIB_storage_data_f_3__1_),
	.ck(clk),
	.d(n12083));
   ms00f80 east_input_NIB_storage_data_f_reg_3__2_ (.o(east_input_NIB_storage_data_f_3__2_),
	.ck(clk),
	.d(n12078));
   ms00f80 east_input_NIB_storage_data_f_reg_3__3_ (.o(east_input_NIB_storage_data_f_3__3_),
	.ck(clk),
	.d(n12073));
   ms00f80 east_input_NIB_storage_data_f_reg_3__4_ (.o(east_input_NIB_storage_data_f_3__4_),
	.ck(clk),
	.d(n12068));
   ms00f80 east_input_NIB_storage_data_f_reg_3__5_ (.o(east_input_NIB_storage_data_f_3__5_),
	.ck(clk),
	.d(n12063));
   ms00f80 east_input_NIB_storage_data_f_reg_3__6_ (.o(east_input_NIB_storage_data_f_3__6_),
	.ck(clk),
	.d(n12058));
   ms00f80 east_input_NIB_storage_data_f_reg_3__7_ (.o(east_input_NIB_storage_data_f_3__7_),
	.ck(clk),
	.d(n12053));
   ms00f80 east_input_NIB_storage_data_f_reg_3__8_ (.o(east_input_NIB_storage_data_f_3__8_),
	.ck(clk),
	.d(n12048));
   ms00f80 east_input_NIB_storage_data_f_reg_3__9_ (.o(east_input_NIB_storage_data_f_3__9_),
	.ck(clk),
	.d(n12043));
   ms00f80 east_input_NIB_storage_data_f_reg_3__10_ (.o(east_input_NIB_storage_data_f_3__10_),
	.ck(clk),
	.d(n12038));
   ms00f80 east_input_NIB_storage_data_f_reg_3__11_ (.o(east_input_NIB_storage_data_f_3__11_),
	.ck(clk),
	.d(n12033));
   ms00f80 east_input_NIB_storage_data_f_reg_3__12_ (.o(east_input_NIB_storage_data_f_3__12_),
	.ck(clk),
	.d(n12028));
   ms00f80 east_input_NIB_storage_data_f_reg_3__13_ (.o(east_input_NIB_storage_data_f_3__13_),
	.ck(clk),
	.d(n12023));
   ms00f80 east_input_NIB_storage_data_f_reg_3__14_ (.o(east_input_NIB_storage_data_f_3__14_),
	.ck(clk),
	.d(n12018));
   ms00f80 east_input_NIB_storage_data_f_reg_3__15_ (.o(east_input_NIB_storage_data_f_3__15_),
	.ck(clk),
	.d(n12013));
   ms00f80 east_input_NIB_storage_data_f_reg_3__16_ (.o(east_input_NIB_storage_data_f_3__16_),
	.ck(clk),
	.d(n12008));
   ms00f80 east_input_NIB_storage_data_f_reg_3__17_ (.o(east_input_NIB_storage_data_f_3__17_),
	.ck(clk),
	.d(n12003));
   ms00f80 east_input_NIB_storage_data_f_reg_3__18_ (.o(east_input_NIB_storage_data_f_3__18_),
	.ck(clk),
	.d(n11998));
   ms00f80 east_input_NIB_storage_data_f_reg_3__19_ (.o(east_input_NIB_storage_data_f_3__19_),
	.ck(clk),
	.d(n11993));
   ms00f80 east_input_NIB_storage_data_f_reg_3__20_ (.o(east_input_NIB_storage_data_f_3__20_),
	.ck(clk),
	.d(n11988));
   ms00f80 east_input_NIB_storage_data_f_reg_3__21_ (.o(east_input_NIB_storage_data_f_3__21_),
	.ck(clk),
	.d(n11983));
   ms00f80 east_input_NIB_storage_data_f_reg_3__22_ (.o(east_input_NIB_storage_data_f_3__22_),
	.ck(clk),
	.d(n11978));
   ms00f80 east_input_NIB_storage_data_f_reg_3__23_ (.o(east_input_NIB_storage_data_f_3__23_),
	.ck(clk),
	.d(n11973));
   ms00f80 east_input_NIB_storage_data_f_reg_3__24_ (.o(east_input_NIB_storage_data_f_3__24_),
	.ck(clk),
	.d(n11968));
   ms00f80 east_input_NIB_storage_data_f_reg_3__25_ (.o(east_input_NIB_storage_data_f_3__25_),
	.ck(clk),
	.d(n11963));
   ms00f80 east_input_NIB_storage_data_f_reg_3__26_ (.o(east_input_NIB_storage_data_f_3__26_),
	.ck(clk),
	.d(n11958));
   ms00f80 east_input_NIB_storage_data_f_reg_3__27_ (.o(east_input_NIB_storage_data_f_3__27_),
	.ck(clk),
	.d(n11953));
   ms00f80 east_input_NIB_storage_data_f_reg_3__28_ (.o(east_input_NIB_storage_data_f_3__28_),
	.ck(clk),
	.d(n11948));
   ms00f80 east_input_NIB_storage_data_f_reg_3__29_ (.o(east_input_NIB_storage_data_f_3__29_),
	.ck(clk),
	.d(n11943));
   ms00f80 east_input_NIB_storage_data_f_reg_3__30_ (.o(east_input_NIB_storage_data_f_3__30_),
	.ck(clk),
	.d(n11938));
   ms00f80 east_input_NIB_storage_data_f_reg_3__31_ (.o(east_input_NIB_storage_data_f_3__31_),
	.ck(clk),
	.d(n11933));
   ms00f80 east_input_NIB_storage_data_f_reg_3__32_ (.o(east_input_NIB_storage_data_f_3__32_),
	.ck(clk),
	.d(n11928));
   ms00f80 east_input_NIB_storage_data_f_reg_3__33_ (.o(east_input_NIB_storage_data_f_3__33_),
	.ck(clk),
	.d(n11923));
   ms00f80 east_input_NIB_storage_data_f_reg_3__34_ (.o(east_input_NIB_storage_data_f_3__34_),
	.ck(clk),
	.d(n11918));
   ms00f80 east_input_NIB_storage_data_f_reg_3__35_ (.o(east_input_NIB_storage_data_f_3__35_),
	.ck(clk),
	.d(n11913));
   ms00f80 east_input_NIB_storage_data_f_reg_3__36_ (.o(east_input_NIB_storage_data_f_3__36_),
	.ck(clk),
	.d(n11908));
   ms00f80 east_input_NIB_storage_data_f_reg_3__37_ (.o(east_input_NIB_storage_data_f_3__37_),
	.ck(clk),
	.d(n11903));
   ms00f80 east_input_NIB_storage_data_f_reg_3__38_ (.o(east_input_NIB_storage_data_f_3__38_),
	.ck(clk),
	.d(n11898));
   ms00f80 east_input_NIB_storage_data_f_reg_3__39_ (.o(east_input_NIB_storage_data_f_3__39_),
	.ck(clk),
	.d(n11893));
   ms00f80 east_input_NIB_storage_data_f_reg_3__40_ (.o(east_input_NIB_storage_data_f_3__40_),
	.ck(clk),
	.d(n11888));
   ms00f80 east_input_NIB_storage_data_f_reg_3__41_ (.o(east_input_NIB_storage_data_f_3__41_),
	.ck(clk),
	.d(n11883));
   ms00f80 east_input_NIB_storage_data_f_reg_3__42_ (.o(east_input_NIB_storage_data_f_3__42_),
	.ck(clk),
	.d(n11878));
   ms00f80 east_input_NIB_storage_data_f_reg_3__43_ (.o(east_input_NIB_storage_data_f_3__43_),
	.ck(clk),
	.d(n11873));
   ms00f80 east_input_NIB_storage_data_f_reg_3__44_ (.o(east_input_NIB_storage_data_f_3__44_),
	.ck(clk),
	.d(n11868));
   ms00f80 east_input_NIB_storage_data_f_reg_3__45_ (.o(east_input_NIB_storage_data_f_3__45_),
	.ck(clk),
	.d(n11863));
   ms00f80 east_input_NIB_storage_data_f_reg_3__46_ (.o(east_input_NIB_storage_data_f_3__46_),
	.ck(clk),
	.d(n11858));
   ms00f80 east_input_NIB_storage_data_f_reg_3__47_ (.o(east_input_NIB_storage_data_f_3__47_),
	.ck(clk),
	.d(n11853));
   ms00f80 east_input_NIB_storage_data_f_reg_3__48_ (.o(east_input_NIB_storage_data_f_3__48_),
	.ck(clk),
	.d(n11848));
   ms00f80 east_input_NIB_storage_data_f_reg_3__49_ (.o(east_input_NIB_storage_data_f_3__49_),
	.ck(clk),
	.d(n11843));
   ms00f80 east_input_NIB_storage_data_f_reg_3__50_ (.o(east_input_NIB_storage_data_f_3__50_),
	.ck(clk),
	.d(n11838));
   ms00f80 east_input_NIB_storage_data_f_reg_3__51_ (.o(east_input_NIB_storage_data_f_3__51_),
	.ck(clk),
	.d(n11833));
   ms00f80 east_input_NIB_storage_data_f_reg_3__52_ (.o(east_input_NIB_storage_data_f_3__52_),
	.ck(clk),
	.d(n11828));
   ms00f80 east_input_NIB_storage_data_f_reg_3__53_ (.o(east_input_NIB_storage_data_f_3__53_),
	.ck(clk),
	.d(n11823));
   ms00f80 east_input_NIB_storage_data_f_reg_3__54_ (.o(east_input_NIB_storage_data_f_3__54_),
	.ck(clk),
	.d(n11818));
   ms00f80 east_input_NIB_storage_data_f_reg_3__55_ (.o(east_input_NIB_storage_data_f_3__55_),
	.ck(clk),
	.d(n11813));
   ms00f80 east_input_NIB_storage_data_f_reg_3__56_ (.o(east_input_NIB_storage_data_f_3__56_),
	.ck(clk),
	.d(n11808));
   ms00f80 east_input_NIB_storage_data_f_reg_3__57_ (.o(east_input_NIB_storage_data_f_3__57_),
	.ck(clk),
	.d(n11803));
   ms00f80 east_input_NIB_storage_data_f_reg_3__58_ (.o(east_input_NIB_storage_data_f_3__58_),
	.ck(clk),
	.d(n11798));
   ms00f80 east_input_NIB_storage_data_f_reg_3__59_ (.o(east_input_NIB_storage_data_f_3__59_),
	.ck(clk),
	.d(n11793));
   ms00f80 east_input_NIB_storage_data_f_reg_3__60_ (.o(east_input_NIB_storage_data_f_3__60_),
	.ck(clk),
	.d(n11788));
   ms00f80 east_input_NIB_storage_data_f_reg_3__61_ (.o(east_input_NIB_storage_data_f_3__61_),
	.ck(clk),
	.d(n11783));
   ms00f80 east_input_NIB_storage_data_f_reg_3__62_ (.o(east_input_NIB_storage_data_f_3__62_),
	.ck(clk),
	.d(n11778));
   ms00f80 east_input_NIB_storage_data_f_reg_3__63_ (.o(east_input_NIB_storage_data_f_3__63_),
	.ck(clk),
	.d(n11773));
   ms00f80 east_input_NIB_storage_data_f_reg_2__0_ (.o(east_input_NIB_storage_data_f_2__0_),
	.ck(clk),
	.d(n11768));
   ms00f80 east_input_NIB_storage_data_f_reg_2__1_ (.o(east_input_NIB_storage_data_f_2__1_),
	.ck(clk),
	.d(n11763));
   ms00f80 east_input_NIB_storage_data_f_reg_2__2_ (.o(east_input_NIB_storage_data_f_2__2_),
	.ck(clk),
	.d(n11758));
   ms00f80 east_input_NIB_storage_data_f_reg_2__3_ (.o(east_input_NIB_storage_data_f_2__3_),
	.ck(clk),
	.d(n11753));
   ms00f80 east_input_NIB_storage_data_f_reg_2__4_ (.o(east_input_NIB_storage_data_f_2__4_),
	.ck(clk),
	.d(n11748));
   ms00f80 east_input_NIB_storage_data_f_reg_2__5_ (.o(east_input_NIB_storage_data_f_2__5_),
	.ck(clk),
	.d(n11743));
   ms00f80 east_input_NIB_storage_data_f_reg_2__6_ (.o(east_input_NIB_storage_data_f_2__6_),
	.ck(clk),
	.d(n11738));
   ms00f80 east_input_NIB_storage_data_f_reg_2__7_ (.o(east_input_NIB_storage_data_f_2__7_),
	.ck(clk),
	.d(n11733));
   ms00f80 east_input_NIB_storage_data_f_reg_2__8_ (.o(east_input_NIB_storage_data_f_2__8_),
	.ck(clk),
	.d(n11728));
   ms00f80 east_input_NIB_storage_data_f_reg_2__9_ (.o(east_input_NIB_storage_data_f_2__9_),
	.ck(clk),
	.d(n11723));
   ms00f80 east_input_NIB_storage_data_f_reg_2__10_ (.o(east_input_NIB_storage_data_f_2__10_),
	.ck(clk),
	.d(n11718));
   ms00f80 east_input_NIB_storage_data_f_reg_2__11_ (.o(east_input_NIB_storage_data_f_2__11_),
	.ck(clk),
	.d(n11713));
   ms00f80 east_input_NIB_storage_data_f_reg_2__12_ (.o(east_input_NIB_storage_data_f_2__12_),
	.ck(clk),
	.d(n11708));
   ms00f80 east_input_NIB_storage_data_f_reg_2__13_ (.o(east_input_NIB_storage_data_f_2__13_),
	.ck(clk),
	.d(n11703));
   ms00f80 east_input_NIB_storage_data_f_reg_2__14_ (.o(east_input_NIB_storage_data_f_2__14_),
	.ck(clk),
	.d(n11698));
   ms00f80 east_input_NIB_storage_data_f_reg_2__15_ (.o(east_input_NIB_storage_data_f_2__15_),
	.ck(clk),
	.d(n11693));
   ms00f80 east_input_NIB_storage_data_f_reg_2__16_ (.o(east_input_NIB_storage_data_f_2__16_),
	.ck(clk),
	.d(n11688));
   ms00f80 east_input_NIB_storage_data_f_reg_2__17_ (.o(east_input_NIB_storage_data_f_2__17_),
	.ck(clk),
	.d(n11683));
   ms00f80 east_input_NIB_storage_data_f_reg_2__18_ (.o(east_input_NIB_storage_data_f_2__18_),
	.ck(clk),
	.d(n11678));
   ms00f80 east_input_NIB_storage_data_f_reg_2__19_ (.o(east_input_NIB_storage_data_f_2__19_),
	.ck(clk),
	.d(n11673));
   ms00f80 east_input_NIB_storage_data_f_reg_2__20_ (.o(east_input_NIB_storage_data_f_2__20_),
	.ck(clk),
	.d(n11668));
   ms00f80 east_input_NIB_storage_data_f_reg_2__21_ (.o(east_input_NIB_storage_data_f_2__21_),
	.ck(clk),
	.d(n11663));
   ms00f80 east_input_NIB_storage_data_f_reg_2__22_ (.o(east_input_NIB_storage_data_f_2__22_),
	.ck(clk),
	.d(n11658));
   ms00f80 east_input_NIB_storage_data_f_reg_2__23_ (.o(east_input_NIB_storage_data_f_2__23_),
	.ck(clk),
	.d(n11653));
   ms00f80 east_input_NIB_storage_data_f_reg_2__24_ (.o(east_input_NIB_storage_data_f_2__24_),
	.ck(clk),
	.d(n11648));
   ms00f80 east_input_NIB_storage_data_f_reg_2__25_ (.o(east_input_NIB_storage_data_f_2__25_),
	.ck(clk),
	.d(n11643));
   ms00f80 east_input_NIB_storage_data_f_reg_2__26_ (.o(east_input_NIB_storage_data_f_2__26_),
	.ck(clk),
	.d(n11638));
   ms00f80 east_input_NIB_storage_data_f_reg_2__27_ (.o(east_input_NIB_storage_data_f_2__27_),
	.ck(clk),
	.d(n11633));
   ms00f80 east_input_NIB_storage_data_f_reg_2__28_ (.o(east_input_NIB_storage_data_f_2__28_),
	.ck(clk),
	.d(n11628));
   ms00f80 east_input_NIB_storage_data_f_reg_2__29_ (.o(east_input_NIB_storage_data_f_2__29_),
	.ck(clk),
	.d(n11623));
   ms00f80 east_input_NIB_storage_data_f_reg_2__30_ (.o(east_input_NIB_storage_data_f_2__30_),
	.ck(clk),
	.d(n11618));
   ms00f80 east_input_NIB_storage_data_f_reg_2__31_ (.o(east_input_NIB_storage_data_f_2__31_),
	.ck(clk),
	.d(n11613));
   ms00f80 east_input_NIB_storage_data_f_reg_2__32_ (.o(east_input_NIB_storage_data_f_2__32_),
	.ck(clk),
	.d(n11608));
   ms00f80 east_input_NIB_storage_data_f_reg_2__33_ (.o(east_input_NIB_storage_data_f_2__33_),
	.ck(clk),
	.d(n11603));
   ms00f80 east_input_NIB_storage_data_f_reg_2__34_ (.o(east_input_NIB_storage_data_f_2__34_),
	.ck(clk),
	.d(n11598));
   ms00f80 east_input_NIB_storage_data_f_reg_2__35_ (.o(east_input_NIB_storage_data_f_2__35_),
	.ck(clk),
	.d(n11593));
   ms00f80 east_input_NIB_storage_data_f_reg_2__36_ (.o(east_input_NIB_storage_data_f_2__36_),
	.ck(clk),
	.d(n11588));
   ms00f80 east_input_NIB_storage_data_f_reg_2__37_ (.o(east_input_NIB_storage_data_f_2__37_),
	.ck(clk),
	.d(n11583));
   ms00f80 east_input_NIB_storage_data_f_reg_2__38_ (.o(east_input_NIB_storage_data_f_2__38_),
	.ck(clk),
	.d(n11578));
   ms00f80 east_input_NIB_storage_data_f_reg_2__39_ (.o(east_input_NIB_storage_data_f_2__39_),
	.ck(clk),
	.d(n11573));
   ms00f80 east_input_NIB_storage_data_f_reg_2__40_ (.o(east_input_NIB_storage_data_f_2__40_),
	.ck(clk),
	.d(n11568));
   ms00f80 east_input_NIB_storage_data_f_reg_2__41_ (.o(east_input_NIB_storage_data_f_2__41_),
	.ck(clk),
	.d(n11563));
   ms00f80 east_input_NIB_storage_data_f_reg_2__42_ (.o(east_input_NIB_storage_data_f_2__42_),
	.ck(clk),
	.d(n11558));
   ms00f80 east_input_NIB_storage_data_f_reg_2__43_ (.o(east_input_NIB_storage_data_f_2__43_),
	.ck(clk),
	.d(n11553));
   ms00f80 east_input_NIB_storage_data_f_reg_2__44_ (.o(east_input_NIB_storage_data_f_2__44_),
	.ck(clk),
	.d(n11548));
   ms00f80 east_input_NIB_storage_data_f_reg_2__45_ (.o(east_input_NIB_storage_data_f_2__45_),
	.ck(clk),
	.d(n11543));
   ms00f80 east_input_NIB_storage_data_f_reg_2__46_ (.o(east_input_NIB_storage_data_f_2__46_),
	.ck(clk),
	.d(n11538));
   ms00f80 east_input_NIB_storage_data_f_reg_2__47_ (.o(east_input_NIB_storage_data_f_2__47_),
	.ck(clk),
	.d(n11533));
   ms00f80 east_input_NIB_storage_data_f_reg_2__48_ (.o(east_input_NIB_storage_data_f_2__48_),
	.ck(clk),
	.d(n11528));
   ms00f80 east_input_NIB_storage_data_f_reg_2__49_ (.o(east_input_NIB_storage_data_f_2__49_),
	.ck(clk),
	.d(n11523));
   ms00f80 east_input_NIB_storage_data_f_reg_2__50_ (.o(east_input_NIB_storage_data_f_2__50_),
	.ck(clk),
	.d(n11518));
   ms00f80 east_input_NIB_storage_data_f_reg_2__51_ (.o(east_input_NIB_storage_data_f_2__51_),
	.ck(clk),
	.d(n11513));
   ms00f80 east_input_NIB_storage_data_f_reg_2__52_ (.o(east_input_NIB_storage_data_f_2__52_),
	.ck(clk),
	.d(n11508));
   ms00f80 east_input_NIB_storage_data_f_reg_2__53_ (.o(east_input_NIB_storage_data_f_2__53_),
	.ck(clk),
	.d(n11503));
   ms00f80 east_input_NIB_storage_data_f_reg_2__54_ (.o(east_input_NIB_storage_data_f_2__54_),
	.ck(clk),
	.d(n11498));
   ms00f80 east_input_NIB_storage_data_f_reg_2__55_ (.o(east_input_NIB_storage_data_f_2__55_),
	.ck(clk),
	.d(n11493));
   ms00f80 east_input_NIB_storage_data_f_reg_2__56_ (.o(east_input_NIB_storage_data_f_2__56_),
	.ck(clk),
	.d(n11488));
   ms00f80 east_input_NIB_storage_data_f_reg_2__57_ (.o(east_input_NIB_storage_data_f_2__57_),
	.ck(clk),
	.d(n11483));
   ms00f80 east_input_NIB_storage_data_f_reg_2__58_ (.o(east_input_NIB_storage_data_f_2__58_),
	.ck(clk),
	.d(n11478));
   ms00f80 east_input_NIB_storage_data_f_reg_2__59_ (.o(east_input_NIB_storage_data_f_2__59_),
	.ck(clk),
	.d(n11473));
   ms00f80 east_input_NIB_storage_data_f_reg_2__60_ (.o(east_input_NIB_storage_data_f_2__60_),
	.ck(clk),
	.d(n11468));
   ms00f80 east_input_NIB_storage_data_f_reg_2__61_ (.o(east_input_NIB_storage_data_f_2__61_),
	.ck(clk),
	.d(n11463));
   ms00f80 east_input_NIB_storage_data_f_reg_2__62_ (.o(east_input_NIB_storage_data_f_2__62_),
	.ck(clk),
	.d(n11458));
   ms00f80 east_input_NIB_storage_data_f_reg_2__63_ (.o(east_input_NIB_storage_data_f_2__63_),
	.ck(clk),
	.d(n11453));
   ms00f80 east_input_NIB_storage_data_f_reg_1__0_ (.o(east_input_NIB_storage_data_f_1__0_),
	.ck(clk),
	.d(n11448));
   ms00f80 east_input_NIB_storage_data_f_reg_1__1_ (.o(east_input_NIB_storage_data_f_1__1_),
	.ck(clk),
	.d(n11443));
   ms00f80 east_input_NIB_storage_data_f_reg_1__2_ (.o(east_input_NIB_storage_data_f_1__2_),
	.ck(clk),
	.d(n11438));
   ms00f80 east_input_NIB_storage_data_f_reg_1__3_ (.o(east_input_NIB_storage_data_f_1__3_),
	.ck(clk),
	.d(n11433));
   ms00f80 east_input_NIB_storage_data_f_reg_1__4_ (.o(east_input_NIB_storage_data_f_1__4_),
	.ck(clk),
	.d(n11428));
   ms00f80 east_input_NIB_storage_data_f_reg_1__5_ (.o(east_input_NIB_storage_data_f_1__5_),
	.ck(clk),
	.d(n11423));
   ms00f80 east_input_NIB_storage_data_f_reg_1__6_ (.o(east_input_NIB_storage_data_f_1__6_),
	.ck(clk),
	.d(n11418));
   ms00f80 east_input_NIB_storage_data_f_reg_1__7_ (.o(east_input_NIB_storage_data_f_1__7_),
	.ck(clk),
	.d(n11413));
   ms00f80 east_input_NIB_storage_data_f_reg_1__8_ (.o(east_input_NIB_storage_data_f_1__8_),
	.ck(clk),
	.d(n11408));
   ms00f80 east_input_NIB_storage_data_f_reg_1__9_ (.o(east_input_NIB_storage_data_f_1__9_),
	.ck(clk),
	.d(n11403));
   ms00f80 east_input_NIB_storage_data_f_reg_1__10_ (.o(east_input_NIB_storage_data_f_1__10_),
	.ck(clk),
	.d(n11398));
   ms00f80 east_input_NIB_storage_data_f_reg_1__11_ (.o(east_input_NIB_storage_data_f_1__11_),
	.ck(clk),
	.d(n11393));
   ms00f80 east_input_NIB_storage_data_f_reg_1__12_ (.o(east_input_NIB_storage_data_f_1__12_),
	.ck(clk),
	.d(n11388));
   ms00f80 east_input_NIB_storage_data_f_reg_1__13_ (.o(east_input_NIB_storage_data_f_1__13_),
	.ck(clk),
	.d(n11383));
   ms00f80 east_input_NIB_storage_data_f_reg_1__14_ (.o(east_input_NIB_storage_data_f_1__14_),
	.ck(clk),
	.d(n11378));
   ms00f80 east_input_NIB_storage_data_f_reg_1__15_ (.o(east_input_NIB_storage_data_f_1__15_),
	.ck(clk),
	.d(n11373));
   ms00f80 east_input_NIB_storage_data_f_reg_1__16_ (.o(east_input_NIB_storage_data_f_1__16_),
	.ck(clk),
	.d(n11368));
   ms00f80 east_input_NIB_storage_data_f_reg_1__17_ (.o(east_input_NIB_storage_data_f_1__17_),
	.ck(clk),
	.d(n11363));
   ms00f80 east_input_NIB_storage_data_f_reg_1__18_ (.o(east_input_NIB_storage_data_f_1__18_),
	.ck(clk),
	.d(n11358));
   ms00f80 east_input_NIB_storage_data_f_reg_1__19_ (.o(east_input_NIB_storage_data_f_1__19_),
	.ck(clk),
	.d(n11353));
   ms00f80 east_input_NIB_storage_data_f_reg_1__20_ (.o(east_input_NIB_storage_data_f_1__20_),
	.ck(clk),
	.d(n11348));
   ms00f80 east_input_NIB_storage_data_f_reg_1__21_ (.o(east_input_NIB_storage_data_f_1__21_),
	.ck(clk),
	.d(n11343));
   ms00f80 east_input_NIB_storage_data_f_reg_1__22_ (.o(east_input_NIB_storage_data_f_1__22_),
	.ck(clk),
	.d(n11338));
   ms00f80 east_input_NIB_storage_data_f_reg_1__23_ (.o(east_input_NIB_storage_data_f_1__23_),
	.ck(clk),
	.d(n11333));
   ms00f80 east_input_NIB_storage_data_f_reg_1__24_ (.o(east_input_NIB_storage_data_f_1__24_),
	.ck(clk),
	.d(n11328));
   ms00f80 east_input_NIB_storage_data_f_reg_1__25_ (.o(east_input_NIB_storage_data_f_1__25_),
	.ck(clk),
	.d(n11323));
   ms00f80 east_input_NIB_storage_data_f_reg_1__26_ (.o(east_input_NIB_storage_data_f_1__26_),
	.ck(clk),
	.d(n11318));
   ms00f80 east_input_NIB_storage_data_f_reg_1__27_ (.o(east_input_NIB_storage_data_f_1__27_),
	.ck(clk),
	.d(n11313));
   ms00f80 east_input_NIB_storage_data_f_reg_1__28_ (.o(east_input_NIB_storage_data_f_1__28_),
	.ck(clk),
	.d(n11308));
   ms00f80 east_input_NIB_storage_data_f_reg_1__29_ (.o(east_input_NIB_storage_data_f_1__29_),
	.ck(clk),
	.d(n11303));
   ms00f80 east_input_NIB_storage_data_f_reg_1__30_ (.o(east_input_NIB_storage_data_f_1__30_),
	.ck(clk),
	.d(n11298));
   ms00f80 east_input_NIB_storage_data_f_reg_1__31_ (.o(east_input_NIB_storage_data_f_1__31_),
	.ck(clk),
	.d(n11293));
   ms00f80 east_input_NIB_storage_data_f_reg_1__32_ (.o(east_input_NIB_storage_data_f_1__32_),
	.ck(clk),
	.d(n11288));
   ms00f80 east_input_NIB_storage_data_f_reg_1__33_ (.o(east_input_NIB_storage_data_f_1__33_),
	.ck(clk),
	.d(n11283));
   ms00f80 east_input_NIB_storage_data_f_reg_1__34_ (.o(east_input_NIB_storage_data_f_1__34_),
	.ck(clk),
	.d(n11278));
   ms00f80 east_input_NIB_storage_data_f_reg_1__35_ (.o(east_input_NIB_storage_data_f_1__35_),
	.ck(clk),
	.d(n11273));
   ms00f80 east_input_NIB_storage_data_f_reg_1__36_ (.o(east_input_NIB_storage_data_f_1__36_),
	.ck(clk),
	.d(n11268));
   ms00f80 east_input_NIB_storage_data_f_reg_1__37_ (.o(east_input_NIB_storage_data_f_1__37_),
	.ck(clk),
	.d(n11263));
   ms00f80 east_input_NIB_storage_data_f_reg_1__38_ (.o(east_input_NIB_storage_data_f_1__38_),
	.ck(clk),
	.d(n11258));
   ms00f80 east_input_NIB_storage_data_f_reg_1__39_ (.o(east_input_NIB_storage_data_f_1__39_),
	.ck(clk),
	.d(n11253));
   ms00f80 east_input_NIB_storage_data_f_reg_1__40_ (.o(east_input_NIB_storage_data_f_1__40_),
	.ck(clk),
	.d(n11248));
   ms00f80 east_input_NIB_storage_data_f_reg_1__41_ (.o(east_input_NIB_storage_data_f_1__41_),
	.ck(clk),
	.d(n11243));
   ms00f80 east_input_NIB_storage_data_f_reg_1__42_ (.o(east_input_NIB_storage_data_f_1__42_),
	.ck(clk),
	.d(n11238));
   ms00f80 east_input_NIB_storage_data_f_reg_1__43_ (.o(east_input_NIB_storage_data_f_1__43_),
	.ck(clk),
	.d(n11233));
   ms00f80 east_input_NIB_storage_data_f_reg_1__44_ (.o(east_input_NIB_storage_data_f_1__44_),
	.ck(clk),
	.d(n11228));
   ms00f80 east_input_NIB_storage_data_f_reg_1__45_ (.o(east_input_NIB_storage_data_f_1__45_),
	.ck(clk),
	.d(n11223));
   ms00f80 east_input_NIB_storage_data_f_reg_1__46_ (.o(east_input_NIB_storage_data_f_1__46_),
	.ck(clk),
	.d(n11218));
   ms00f80 east_input_NIB_storage_data_f_reg_1__47_ (.o(east_input_NIB_storage_data_f_1__47_),
	.ck(clk),
	.d(n11213));
   ms00f80 east_input_NIB_storage_data_f_reg_1__48_ (.o(east_input_NIB_storage_data_f_1__48_),
	.ck(clk),
	.d(n11208));
   ms00f80 east_input_NIB_storage_data_f_reg_1__49_ (.o(east_input_NIB_storage_data_f_1__49_),
	.ck(clk),
	.d(n11203));
   ms00f80 east_input_NIB_storage_data_f_reg_1__50_ (.o(east_input_NIB_storage_data_f_1__50_),
	.ck(clk),
	.d(n11198));
   ms00f80 east_input_NIB_storage_data_f_reg_1__51_ (.o(east_input_NIB_storage_data_f_1__51_),
	.ck(clk),
	.d(n11193));
   ms00f80 east_input_NIB_storage_data_f_reg_1__52_ (.o(east_input_NIB_storage_data_f_1__52_),
	.ck(clk),
	.d(n11188));
   ms00f80 east_input_NIB_storage_data_f_reg_1__53_ (.o(east_input_NIB_storage_data_f_1__53_),
	.ck(clk),
	.d(n11183));
   ms00f80 east_input_NIB_storage_data_f_reg_1__54_ (.o(east_input_NIB_storage_data_f_1__54_),
	.ck(clk),
	.d(n11178));
   ms00f80 east_input_NIB_storage_data_f_reg_1__55_ (.o(east_input_NIB_storage_data_f_1__55_),
	.ck(clk),
	.d(n11173));
   ms00f80 east_input_NIB_storage_data_f_reg_1__56_ (.o(east_input_NIB_storage_data_f_1__56_),
	.ck(clk),
	.d(n11168));
   ms00f80 east_input_NIB_storage_data_f_reg_1__57_ (.o(east_input_NIB_storage_data_f_1__57_),
	.ck(clk),
	.d(n11163));
   ms00f80 east_input_NIB_storage_data_f_reg_1__58_ (.o(east_input_NIB_storage_data_f_1__58_),
	.ck(clk),
	.d(n11158));
   ms00f80 east_input_NIB_storage_data_f_reg_1__59_ (.o(east_input_NIB_storage_data_f_1__59_),
	.ck(clk),
	.d(n11153));
   ms00f80 east_input_NIB_storage_data_f_reg_1__60_ (.o(east_input_NIB_storage_data_f_1__60_),
	.ck(clk),
	.d(n11148));
   ms00f80 east_input_NIB_storage_data_f_reg_1__61_ (.o(east_input_NIB_storage_data_f_1__61_),
	.ck(clk),
	.d(n11143));
   ms00f80 east_input_NIB_storage_data_f_reg_1__62_ (.o(east_input_NIB_storage_data_f_1__62_),
	.ck(clk),
	.d(n11138));
   ms00f80 east_input_NIB_storage_data_f_reg_1__63_ (.o(east_input_NIB_storage_data_f_1__63_),
	.ck(clk),
	.d(n11133));
   ms00f80 east_input_NIB_storage_data_f_reg_0__0_ (.o(east_input_NIB_storage_data_f_0__0_),
	.ck(clk),
	.d(n11128));
   ms00f80 east_input_NIB_storage_data_f_reg_0__1_ (.o(east_input_NIB_storage_data_f_0__1_),
	.ck(clk),
	.d(n11123));
   ms00f80 east_input_NIB_storage_data_f_reg_0__2_ (.o(east_input_NIB_storage_data_f_0__2_),
	.ck(clk),
	.d(n11118));
   ms00f80 east_input_NIB_storage_data_f_reg_0__3_ (.o(east_input_NIB_storage_data_f_0__3_),
	.ck(clk),
	.d(n11113));
   ms00f80 east_input_NIB_storage_data_f_reg_0__4_ (.o(east_input_NIB_storage_data_f_0__4_),
	.ck(clk),
	.d(n11108));
   ms00f80 east_input_NIB_storage_data_f_reg_0__5_ (.o(east_input_NIB_storage_data_f_0__5_),
	.ck(clk),
	.d(n11103));
   ms00f80 east_input_NIB_storage_data_f_reg_0__6_ (.o(east_input_NIB_storage_data_f_0__6_),
	.ck(clk),
	.d(n11098));
   ms00f80 east_input_NIB_storage_data_f_reg_0__7_ (.o(east_input_NIB_storage_data_f_0__7_),
	.ck(clk),
	.d(n11093));
   ms00f80 east_input_NIB_storage_data_f_reg_0__8_ (.o(east_input_NIB_storage_data_f_0__8_),
	.ck(clk),
	.d(n11088));
   ms00f80 east_input_NIB_storage_data_f_reg_0__9_ (.o(east_input_NIB_storage_data_f_0__9_),
	.ck(clk),
	.d(n11083));
   ms00f80 east_input_NIB_storage_data_f_reg_0__10_ (.o(east_input_NIB_storage_data_f_0__10_),
	.ck(clk),
	.d(n11078));
   ms00f80 east_input_NIB_storage_data_f_reg_0__11_ (.o(east_input_NIB_storage_data_f_0__11_),
	.ck(clk),
	.d(n11073));
   ms00f80 east_input_NIB_storage_data_f_reg_0__12_ (.o(east_input_NIB_storage_data_f_0__12_),
	.ck(clk),
	.d(n11068));
   ms00f80 east_input_NIB_storage_data_f_reg_0__13_ (.o(east_input_NIB_storage_data_f_0__13_),
	.ck(clk),
	.d(n11063));
   ms00f80 east_input_NIB_storage_data_f_reg_0__14_ (.o(east_input_NIB_storage_data_f_0__14_),
	.ck(clk),
	.d(n11058));
   ms00f80 east_input_NIB_storage_data_f_reg_0__15_ (.o(east_input_NIB_storage_data_f_0__15_),
	.ck(clk),
	.d(n11053));
   ms00f80 east_input_NIB_storage_data_f_reg_0__16_ (.o(east_input_NIB_storage_data_f_0__16_),
	.ck(clk),
	.d(n11048));
   ms00f80 east_input_NIB_storage_data_f_reg_0__17_ (.o(east_input_NIB_storage_data_f_0__17_),
	.ck(clk),
	.d(n11043));
   ms00f80 east_input_NIB_storage_data_f_reg_0__18_ (.o(east_input_NIB_storage_data_f_0__18_),
	.ck(clk),
	.d(n11038));
   ms00f80 east_input_NIB_storage_data_f_reg_0__19_ (.o(east_input_NIB_storage_data_f_0__19_),
	.ck(clk),
	.d(n11033));
   ms00f80 east_input_NIB_storage_data_f_reg_0__20_ (.o(east_input_NIB_storage_data_f_0__20_),
	.ck(clk),
	.d(n11028));
   ms00f80 east_input_NIB_storage_data_f_reg_0__21_ (.o(east_input_NIB_storage_data_f_0__21_),
	.ck(clk),
	.d(n11023));
   ms00f80 east_input_NIB_storage_data_f_reg_0__22_ (.o(east_input_NIB_storage_data_f_0__22_),
	.ck(clk),
	.d(n11018));
   ms00f80 east_input_NIB_storage_data_f_reg_0__23_ (.o(east_input_NIB_storage_data_f_0__23_),
	.ck(clk),
	.d(n11013));
   ms00f80 east_input_NIB_storage_data_f_reg_0__24_ (.o(east_input_NIB_storage_data_f_0__24_),
	.ck(clk),
	.d(n11008));
   ms00f80 east_input_NIB_storage_data_f_reg_0__25_ (.o(east_input_NIB_storage_data_f_0__25_),
	.ck(clk),
	.d(n11003));
   ms00f80 east_input_NIB_storage_data_f_reg_0__26_ (.o(east_input_NIB_storage_data_f_0__26_),
	.ck(clk),
	.d(n10998));
   ms00f80 east_input_NIB_storage_data_f_reg_0__27_ (.o(east_input_NIB_storage_data_f_0__27_),
	.ck(clk),
	.d(n10993));
   ms00f80 east_input_NIB_storage_data_f_reg_0__28_ (.o(east_input_NIB_storage_data_f_0__28_),
	.ck(clk),
	.d(n10988));
   ms00f80 east_input_NIB_storage_data_f_reg_0__29_ (.o(east_input_NIB_storage_data_f_0__29_),
	.ck(clk),
	.d(n10983));
   ms00f80 east_input_NIB_storage_data_f_reg_0__30_ (.o(east_input_NIB_storage_data_f_0__30_),
	.ck(clk),
	.d(n10978));
   ms00f80 east_input_NIB_storage_data_f_reg_0__31_ (.o(east_input_NIB_storage_data_f_0__31_),
	.ck(clk),
	.d(n10973));
   ms00f80 east_input_NIB_storage_data_f_reg_0__32_ (.o(east_input_NIB_storage_data_f_0__32_),
	.ck(clk),
	.d(n10968));
   ms00f80 east_input_NIB_storage_data_f_reg_0__33_ (.o(east_input_NIB_storage_data_f_0__33_),
	.ck(clk),
	.d(n10963));
   ms00f80 east_input_NIB_storage_data_f_reg_0__34_ (.o(east_input_NIB_storage_data_f_0__34_),
	.ck(clk),
	.d(n10958));
   ms00f80 east_input_NIB_storage_data_f_reg_0__35_ (.o(east_input_NIB_storage_data_f_0__35_),
	.ck(clk),
	.d(n10953));
   ms00f80 east_input_NIB_storage_data_f_reg_0__36_ (.o(east_input_NIB_storage_data_f_0__36_),
	.ck(clk),
	.d(n10948));
   ms00f80 east_input_NIB_storage_data_f_reg_0__37_ (.o(east_input_NIB_storage_data_f_0__37_),
	.ck(clk),
	.d(n10943));
   ms00f80 east_input_NIB_storage_data_f_reg_0__38_ (.o(east_input_NIB_storage_data_f_0__38_),
	.ck(clk),
	.d(n10938));
   ms00f80 east_input_NIB_storage_data_f_reg_0__39_ (.o(east_input_NIB_storage_data_f_0__39_),
	.ck(clk),
	.d(n10933));
   ms00f80 east_input_NIB_storage_data_f_reg_0__40_ (.o(east_input_NIB_storage_data_f_0__40_),
	.ck(clk),
	.d(n10928));
   ms00f80 east_input_NIB_storage_data_f_reg_0__41_ (.o(east_input_NIB_storage_data_f_0__41_),
	.ck(clk),
	.d(n10923));
   ms00f80 east_input_NIB_storage_data_f_reg_0__42_ (.o(east_input_NIB_storage_data_f_0__42_),
	.ck(clk),
	.d(n10918));
   ms00f80 east_input_NIB_storage_data_f_reg_0__43_ (.o(east_input_NIB_storage_data_f_0__43_),
	.ck(clk),
	.d(n10913));
   ms00f80 east_input_NIB_storage_data_f_reg_0__44_ (.o(east_input_NIB_storage_data_f_0__44_),
	.ck(clk),
	.d(n10908));
   ms00f80 east_input_NIB_storage_data_f_reg_0__45_ (.o(east_input_NIB_storage_data_f_0__45_),
	.ck(clk),
	.d(n10903));
   ms00f80 east_input_NIB_storage_data_f_reg_0__46_ (.o(east_input_NIB_storage_data_f_0__46_),
	.ck(clk),
	.d(n10898));
   ms00f80 east_input_NIB_storage_data_f_reg_0__47_ (.o(east_input_NIB_storage_data_f_0__47_),
	.ck(clk),
	.d(n10893));
   ms00f80 east_input_NIB_storage_data_f_reg_0__48_ (.o(east_input_NIB_storage_data_f_0__48_),
	.ck(clk),
	.d(n10888));
   ms00f80 east_input_NIB_storage_data_f_reg_0__49_ (.o(east_input_NIB_storage_data_f_0__49_),
	.ck(clk),
	.d(n10883));
   ms00f80 east_input_NIB_storage_data_f_reg_0__50_ (.o(east_input_NIB_storage_data_f_0__50_),
	.ck(clk),
	.d(n10878));
   ms00f80 east_input_NIB_storage_data_f_reg_0__51_ (.o(east_input_NIB_storage_data_f_0__51_),
	.ck(clk),
	.d(n10873));
   ms00f80 east_input_NIB_storage_data_f_reg_0__52_ (.o(east_input_NIB_storage_data_f_0__52_),
	.ck(clk),
	.d(n10868));
   ms00f80 east_input_NIB_storage_data_f_reg_0__53_ (.o(east_input_NIB_storage_data_f_0__53_),
	.ck(clk),
	.d(n10863));
   ms00f80 east_input_NIB_storage_data_f_reg_0__54_ (.o(east_input_NIB_storage_data_f_0__54_),
	.ck(clk),
	.d(n10858));
   ms00f80 east_input_NIB_storage_data_f_reg_0__55_ (.o(east_input_NIB_storage_data_f_0__55_),
	.ck(clk),
	.d(n10853));
   ms00f80 east_input_NIB_storage_data_f_reg_0__56_ (.o(east_input_NIB_storage_data_f_0__56_),
	.ck(clk),
	.d(n10848));
   ms00f80 east_input_NIB_storage_data_f_reg_0__57_ (.o(east_input_NIB_storage_data_f_0__57_),
	.ck(clk),
	.d(n10843));
   ms00f80 east_input_NIB_storage_data_f_reg_0__58_ (.o(east_input_NIB_storage_data_f_0__58_),
	.ck(clk),
	.d(n10838));
   ms00f80 east_input_NIB_storage_data_f_reg_0__59_ (.o(east_input_NIB_storage_data_f_0__59_),
	.ck(clk),
	.d(n10833));
   ms00f80 east_input_NIB_storage_data_f_reg_0__60_ (.o(east_input_NIB_storage_data_f_0__60_),
	.ck(clk),
	.d(n10828));
   ms00f80 east_input_NIB_storage_data_f_reg_0__61_ (.o(east_input_NIB_storage_data_f_0__61_),
	.ck(clk),
	.d(n10823));
   ms00f80 east_input_NIB_storage_data_f_reg_0__62_ (.o(east_input_NIB_storage_data_f_0__62_),
	.ck(clk),
	.d(n10818));
   ms00f80 east_input_NIB_storage_data_f_reg_0__63_ (.o(east_input_NIB_storage_data_f_0__63_),
	.ck(clk),
	.d(n10813));
   ms00f80 south_input_NIB_tail_ptr_f_reg_0_ (.o(south_input_NIB_tail_ptr_f_0_),
	.ck(clk),
	.d(n10808));
   ms00f80 south_input_NIB_tail_ptr_f_reg_1_ (.o(south_input_NIB_tail_ptr_f_1_),
	.ck(clk),
	.d(n10803));
   ms00f80 south_input_NIB_storage_data_f_reg_3__0_ (.o(south_input_NIB_storage_data_f_3__0_),
	.ck(clk),
	.d(n10798));
   ms00f80 south_input_NIB_storage_data_f_reg_3__1_ (.o(south_input_NIB_storage_data_f_3__1_),
	.ck(clk),
	.d(n10793));
   ms00f80 south_input_NIB_storage_data_f_reg_3__2_ (.o(south_input_NIB_storage_data_f_3__2_),
	.ck(clk),
	.d(n10788));
   ms00f80 south_input_NIB_storage_data_f_reg_3__3_ (.o(south_input_NIB_storage_data_f_3__3_),
	.ck(clk),
	.d(n10783));
   ms00f80 south_input_NIB_storage_data_f_reg_3__4_ (.o(south_input_NIB_storage_data_f_3__4_),
	.ck(clk),
	.d(n10778));
   ms00f80 south_input_NIB_storage_data_f_reg_3__5_ (.o(south_input_NIB_storage_data_f_3__5_),
	.ck(clk),
	.d(n10773));
   ms00f80 south_input_NIB_storage_data_f_reg_3__6_ (.o(south_input_NIB_storage_data_f_3__6_),
	.ck(clk),
	.d(n10768));
   ms00f80 south_input_NIB_storage_data_f_reg_3__7_ (.o(south_input_NIB_storage_data_f_3__7_),
	.ck(clk),
	.d(n10763));
   ms00f80 south_input_NIB_storage_data_f_reg_3__8_ (.o(south_input_NIB_storage_data_f_3__8_),
	.ck(clk),
	.d(n10758));
   ms00f80 south_input_NIB_storage_data_f_reg_3__9_ (.o(south_input_NIB_storage_data_f_3__9_),
	.ck(clk),
	.d(n10753));
   ms00f80 south_input_NIB_storage_data_f_reg_3__10_ (.o(south_input_NIB_storage_data_f_3__10_),
	.ck(clk),
	.d(n10748));
   ms00f80 south_input_NIB_storage_data_f_reg_3__11_ (.o(south_input_NIB_storage_data_f_3__11_),
	.ck(clk),
	.d(n10743));
   ms00f80 south_input_NIB_storage_data_f_reg_3__12_ (.o(south_input_NIB_storage_data_f_3__12_),
	.ck(clk),
	.d(n10738));
   ms00f80 south_input_NIB_storage_data_f_reg_3__13_ (.o(south_input_NIB_storage_data_f_3__13_),
	.ck(clk),
	.d(n10733));
   ms00f80 south_input_NIB_storage_data_f_reg_3__14_ (.o(south_input_NIB_storage_data_f_3__14_),
	.ck(clk),
	.d(n10728));
   ms00f80 south_input_NIB_storage_data_f_reg_3__15_ (.o(south_input_NIB_storage_data_f_3__15_),
	.ck(clk),
	.d(n10723));
   ms00f80 south_input_NIB_storage_data_f_reg_3__16_ (.o(south_input_NIB_storage_data_f_3__16_),
	.ck(clk),
	.d(n10718));
   ms00f80 south_input_NIB_storage_data_f_reg_3__17_ (.o(south_input_NIB_storage_data_f_3__17_),
	.ck(clk),
	.d(n10713));
   ms00f80 south_input_NIB_storage_data_f_reg_3__18_ (.o(south_input_NIB_storage_data_f_3__18_),
	.ck(clk),
	.d(n10708));
   ms00f80 south_input_NIB_storage_data_f_reg_3__19_ (.o(south_input_NIB_storage_data_f_3__19_),
	.ck(clk),
	.d(n10703));
   ms00f80 south_input_NIB_storage_data_f_reg_3__20_ (.o(south_input_NIB_storage_data_f_3__20_),
	.ck(clk),
	.d(n10698));
   ms00f80 south_input_NIB_storage_data_f_reg_3__21_ (.o(south_input_NIB_storage_data_f_3__21_),
	.ck(clk),
	.d(n10693));
   ms00f80 south_input_NIB_storage_data_f_reg_3__22_ (.o(south_input_NIB_storage_data_f_3__22_),
	.ck(clk),
	.d(n10688));
   ms00f80 south_input_NIB_storage_data_f_reg_3__23_ (.o(south_input_NIB_storage_data_f_3__23_),
	.ck(clk),
	.d(n10683));
   ms00f80 south_input_NIB_storage_data_f_reg_3__24_ (.o(south_input_NIB_storage_data_f_3__24_),
	.ck(clk),
	.d(n10678));
   ms00f80 south_input_NIB_storage_data_f_reg_3__25_ (.o(south_input_NIB_storage_data_f_3__25_),
	.ck(clk),
	.d(n10673));
   ms00f80 south_input_NIB_storage_data_f_reg_3__26_ (.o(south_input_NIB_storage_data_f_3__26_),
	.ck(clk),
	.d(n10668));
   ms00f80 south_input_NIB_storage_data_f_reg_3__27_ (.o(south_input_NIB_storage_data_f_3__27_),
	.ck(clk),
	.d(n10663));
   ms00f80 south_input_NIB_storage_data_f_reg_3__28_ (.o(south_input_NIB_storage_data_f_3__28_),
	.ck(clk),
	.d(n10658));
   ms00f80 south_input_NIB_storage_data_f_reg_3__29_ (.o(south_input_NIB_storage_data_f_3__29_),
	.ck(clk),
	.d(n10653));
   ms00f80 south_input_NIB_storage_data_f_reg_3__30_ (.o(south_input_NIB_storage_data_f_3__30_),
	.ck(clk),
	.d(n10648));
   ms00f80 south_input_NIB_storage_data_f_reg_3__31_ (.o(south_input_NIB_storage_data_f_3__31_),
	.ck(clk),
	.d(n10643));
   ms00f80 south_input_NIB_storage_data_f_reg_3__32_ (.o(south_input_NIB_storage_data_f_3__32_),
	.ck(clk),
	.d(n10638));
   ms00f80 south_input_NIB_storage_data_f_reg_3__33_ (.o(south_input_NIB_storage_data_f_3__33_),
	.ck(clk),
	.d(n10633));
   ms00f80 south_input_NIB_storage_data_f_reg_3__34_ (.o(south_input_NIB_storage_data_f_3__34_),
	.ck(clk),
	.d(n10628));
   ms00f80 south_input_NIB_storage_data_f_reg_3__35_ (.o(south_input_NIB_storage_data_f_3__35_),
	.ck(clk),
	.d(n10623));
   ms00f80 south_input_NIB_storage_data_f_reg_3__36_ (.o(south_input_NIB_storage_data_f_3__36_),
	.ck(clk),
	.d(n10618));
   ms00f80 south_input_NIB_storage_data_f_reg_3__37_ (.o(south_input_NIB_storage_data_f_3__37_),
	.ck(clk),
	.d(n10613));
   ms00f80 south_input_NIB_storage_data_f_reg_3__38_ (.o(south_input_NIB_storage_data_f_3__38_),
	.ck(clk),
	.d(n10608));
   ms00f80 south_input_NIB_storage_data_f_reg_3__39_ (.o(south_input_NIB_storage_data_f_3__39_),
	.ck(clk),
	.d(n10603));
   ms00f80 south_input_NIB_storage_data_f_reg_3__40_ (.o(south_input_NIB_storage_data_f_3__40_),
	.ck(clk),
	.d(n10598));
   ms00f80 south_input_NIB_storage_data_f_reg_3__41_ (.o(south_input_NIB_storage_data_f_3__41_),
	.ck(clk),
	.d(n10593));
   ms00f80 south_input_NIB_storage_data_f_reg_3__42_ (.o(south_input_NIB_storage_data_f_3__42_),
	.ck(clk),
	.d(n10588));
   ms00f80 south_input_NIB_storage_data_f_reg_3__43_ (.o(south_input_NIB_storage_data_f_3__43_),
	.ck(clk),
	.d(n10583));
   ms00f80 south_input_NIB_storage_data_f_reg_3__44_ (.o(south_input_NIB_storage_data_f_3__44_),
	.ck(clk),
	.d(n10578));
   ms00f80 south_input_NIB_storage_data_f_reg_3__45_ (.o(south_input_NIB_storage_data_f_3__45_),
	.ck(clk),
	.d(n10573));
   ms00f80 south_input_NIB_storage_data_f_reg_3__46_ (.o(south_input_NIB_storage_data_f_3__46_),
	.ck(clk),
	.d(n10568));
   ms00f80 south_input_NIB_storage_data_f_reg_3__47_ (.o(south_input_NIB_storage_data_f_3__47_),
	.ck(clk),
	.d(n10563));
   ms00f80 south_input_NIB_storage_data_f_reg_3__48_ (.o(south_input_NIB_storage_data_f_3__48_),
	.ck(clk),
	.d(n10558));
   ms00f80 south_input_NIB_storage_data_f_reg_3__49_ (.o(south_input_NIB_storage_data_f_3__49_),
	.ck(clk),
	.d(n10553));
   ms00f80 south_input_NIB_storage_data_f_reg_3__50_ (.o(south_input_NIB_storage_data_f_3__50_),
	.ck(clk),
	.d(n10548));
   ms00f80 south_input_NIB_storage_data_f_reg_3__51_ (.o(south_input_NIB_storage_data_f_3__51_),
	.ck(clk),
	.d(n10543));
   ms00f80 south_input_NIB_storage_data_f_reg_3__52_ (.o(south_input_NIB_storage_data_f_3__52_),
	.ck(clk),
	.d(n10538));
   ms00f80 south_input_NIB_storage_data_f_reg_3__53_ (.o(south_input_NIB_storage_data_f_3__53_),
	.ck(clk),
	.d(n10533));
   ms00f80 south_input_NIB_storage_data_f_reg_3__54_ (.o(south_input_NIB_storage_data_f_3__54_),
	.ck(clk),
	.d(n10528));
   ms00f80 south_input_NIB_storage_data_f_reg_3__55_ (.o(south_input_NIB_storage_data_f_3__55_),
	.ck(clk),
	.d(n10523));
   ms00f80 south_input_NIB_storage_data_f_reg_3__56_ (.o(south_input_NIB_storage_data_f_3__56_),
	.ck(clk),
	.d(n10518));
   ms00f80 south_input_NIB_storage_data_f_reg_3__57_ (.o(south_input_NIB_storage_data_f_3__57_),
	.ck(clk),
	.d(n10513));
   ms00f80 south_input_NIB_storage_data_f_reg_3__58_ (.o(south_input_NIB_storage_data_f_3__58_),
	.ck(clk),
	.d(n10508));
   ms00f80 south_input_NIB_storage_data_f_reg_3__59_ (.o(south_input_NIB_storage_data_f_3__59_),
	.ck(clk),
	.d(n10503));
   ms00f80 south_input_NIB_storage_data_f_reg_3__60_ (.o(south_input_NIB_storage_data_f_3__60_),
	.ck(clk),
	.d(n10498));
   ms00f80 south_input_NIB_storage_data_f_reg_3__61_ (.o(south_input_NIB_storage_data_f_3__61_),
	.ck(clk),
	.d(n10493));
   ms00f80 south_input_NIB_storage_data_f_reg_3__62_ (.o(south_input_NIB_storage_data_f_3__62_),
	.ck(clk),
	.d(n10488));
   ms00f80 south_input_NIB_storage_data_f_reg_3__63_ (.o(south_input_NIB_storage_data_f_3__63_),
	.ck(clk),
	.d(n10483));
   ms00f80 south_input_NIB_storage_data_f_reg_2__0_ (.o(south_input_NIB_storage_data_f_2__0_),
	.ck(clk),
	.d(n10478));
   ms00f80 south_input_NIB_storage_data_f_reg_2__1_ (.o(south_input_NIB_storage_data_f_2__1_),
	.ck(clk),
	.d(n10473));
   ms00f80 south_input_NIB_storage_data_f_reg_2__2_ (.o(south_input_NIB_storage_data_f_2__2_),
	.ck(clk),
	.d(n10468));
   ms00f80 south_input_NIB_storage_data_f_reg_2__3_ (.o(south_input_NIB_storage_data_f_2__3_),
	.ck(clk),
	.d(n10463));
   ms00f80 south_input_NIB_storage_data_f_reg_2__4_ (.o(south_input_NIB_storage_data_f_2__4_),
	.ck(clk),
	.d(n10458));
   ms00f80 south_input_NIB_storage_data_f_reg_2__5_ (.o(south_input_NIB_storage_data_f_2__5_),
	.ck(clk),
	.d(n10453));
   ms00f80 south_input_NIB_storage_data_f_reg_2__6_ (.o(south_input_NIB_storage_data_f_2__6_),
	.ck(clk),
	.d(n10448));
   ms00f80 south_input_NIB_storage_data_f_reg_2__7_ (.o(south_input_NIB_storage_data_f_2__7_),
	.ck(clk),
	.d(n10443));
   ms00f80 south_input_NIB_storage_data_f_reg_2__8_ (.o(south_input_NIB_storage_data_f_2__8_),
	.ck(clk),
	.d(n10438));
   ms00f80 south_input_NIB_storage_data_f_reg_2__9_ (.o(south_input_NIB_storage_data_f_2__9_),
	.ck(clk),
	.d(n10433));
   ms00f80 south_input_NIB_storage_data_f_reg_2__10_ (.o(south_input_NIB_storage_data_f_2__10_),
	.ck(clk),
	.d(n10428));
   ms00f80 south_input_NIB_storage_data_f_reg_2__11_ (.o(south_input_NIB_storage_data_f_2__11_),
	.ck(clk),
	.d(n10423));
   ms00f80 south_input_NIB_storage_data_f_reg_2__12_ (.o(south_input_NIB_storage_data_f_2__12_),
	.ck(clk),
	.d(n10418));
   ms00f80 south_input_NIB_storage_data_f_reg_2__13_ (.o(south_input_NIB_storage_data_f_2__13_),
	.ck(clk),
	.d(n10413));
   ms00f80 south_input_NIB_storage_data_f_reg_2__14_ (.o(south_input_NIB_storage_data_f_2__14_),
	.ck(clk),
	.d(n10408));
   ms00f80 south_input_NIB_storage_data_f_reg_2__15_ (.o(south_input_NIB_storage_data_f_2__15_),
	.ck(clk),
	.d(n10403));
   ms00f80 south_input_NIB_storage_data_f_reg_2__16_ (.o(south_input_NIB_storage_data_f_2__16_),
	.ck(clk),
	.d(n10398));
   ms00f80 south_input_NIB_storage_data_f_reg_2__17_ (.o(south_input_NIB_storage_data_f_2__17_),
	.ck(clk),
	.d(n10393));
   ms00f80 south_input_NIB_storage_data_f_reg_2__18_ (.o(south_input_NIB_storage_data_f_2__18_),
	.ck(clk),
	.d(n10388));
   ms00f80 south_input_NIB_storage_data_f_reg_2__19_ (.o(south_input_NIB_storage_data_f_2__19_),
	.ck(clk),
	.d(n10383));
   ms00f80 south_input_NIB_storage_data_f_reg_2__20_ (.o(south_input_NIB_storage_data_f_2__20_),
	.ck(clk),
	.d(n10378));
   ms00f80 south_input_NIB_storage_data_f_reg_2__21_ (.o(south_input_NIB_storage_data_f_2__21_),
	.ck(clk),
	.d(n10373));
   ms00f80 south_input_NIB_storage_data_f_reg_2__22_ (.o(south_input_NIB_storage_data_f_2__22_),
	.ck(clk),
	.d(n10368));
   ms00f80 south_input_NIB_storage_data_f_reg_2__23_ (.o(south_input_NIB_storage_data_f_2__23_),
	.ck(clk),
	.d(n10363));
   ms00f80 south_input_NIB_storage_data_f_reg_2__24_ (.o(south_input_NIB_storage_data_f_2__24_),
	.ck(clk),
	.d(n10358));
   ms00f80 south_input_NIB_storage_data_f_reg_2__25_ (.o(south_input_NIB_storage_data_f_2__25_),
	.ck(clk),
	.d(n10353));
   ms00f80 south_input_NIB_storage_data_f_reg_2__26_ (.o(south_input_NIB_storage_data_f_2__26_),
	.ck(clk),
	.d(n10348));
   ms00f80 south_input_NIB_storage_data_f_reg_2__27_ (.o(south_input_NIB_storage_data_f_2__27_),
	.ck(clk),
	.d(n10343));
   ms00f80 south_input_NIB_storage_data_f_reg_2__28_ (.o(south_input_NIB_storage_data_f_2__28_),
	.ck(clk),
	.d(n10338));
   ms00f80 south_input_NIB_storage_data_f_reg_2__29_ (.o(south_input_NIB_storage_data_f_2__29_),
	.ck(clk),
	.d(n10333));
   ms00f80 south_input_NIB_storage_data_f_reg_2__30_ (.o(south_input_NIB_storage_data_f_2__30_),
	.ck(clk),
	.d(n10328));
   ms00f80 south_input_NIB_storage_data_f_reg_2__31_ (.o(south_input_NIB_storage_data_f_2__31_),
	.ck(clk),
	.d(n10323));
   ms00f80 south_input_NIB_storage_data_f_reg_2__32_ (.o(south_input_NIB_storage_data_f_2__32_),
	.ck(clk),
	.d(n10318));
   ms00f80 south_input_NIB_storage_data_f_reg_2__33_ (.o(south_input_NIB_storage_data_f_2__33_),
	.ck(clk),
	.d(n10313));
   ms00f80 south_input_NIB_storage_data_f_reg_2__34_ (.o(south_input_NIB_storage_data_f_2__34_),
	.ck(clk),
	.d(n10308));
   ms00f80 south_input_NIB_storage_data_f_reg_2__35_ (.o(south_input_NIB_storage_data_f_2__35_),
	.ck(clk),
	.d(n10303));
   ms00f80 south_input_NIB_storage_data_f_reg_2__36_ (.o(south_input_NIB_storage_data_f_2__36_),
	.ck(clk),
	.d(n10298));
   ms00f80 south_input_NIB_storage_data_f_reg_2__37_ (.o(south_input_NIB_storage_data_f_2__37_),
	.ck(clk),
	.d(n10293));
   ms00f80 south_input_NIB_storage_data_f_reg_2__38_ (.o(south_input_NIB_storage_data_f_2__38_),
	.ck(clk),
	.d(n10288));
   ms00f80 south_input_NIB_storage_data_f_reg_2__39_ (.o(south_input_NIB_storage_data_f_2__39_),
	.ck(clk),
	.d(n10283));
   ms00f80 south_input_NIB_storage_data_f_reg_2__40_ (.o(south_input_NIB_storage_data_f_2__40_),
	.ck(clk),
	.d(n10278));
   ms00f80 south_input_NIB_storage_data_f_reg_2__41_ (.o(south_input_NIB_storage_data_f_2__41_),
	.ck(clk),
	.d(n10273));
   ms00f80 south_input_NIB_storage_data_f_reg_2__42_ (.o(south_input_NIB_storage_data_f_2__42_),
	.ck(clk),
	.d(n10268));
   ms00f80 south_input_NIB_storage_data_f_reg_2__43_ (.o(south_input_NIB_storage_data_f_2__43_),
	.ck(clk),
	.d(n10263));
   ms00f80 south_input_NIB_storage_data_f_reg_2__44_ (.o(south_input_NIB_storage_data_f_2__44_),
	.ck(clk),
	.d(n10258));
   ms00f80 south_input_NIB_storage_data_f_reg_2__45_ (.o(south_input_NIB_storage_data_f_2__45_),
	.ck(clk),
	.d(n10253));
   ms00f80 south_input_NIB_storage_data_f_reg_2__46_ (.o(south_input_NIB_storage_data_f_2__46_),
	.ck(clk),
	.d(n10248));
   ms00f80 south_input_NIB_storage_data_f_reg_2__47_ (.o(south_input_NIB_storage_data_f_2__47_),
	.ck(clk),
	.d(n10243));
   ms00f80 south_input_NIB_storage_data_f_reg_2__48_ (.o(south_input_NIB_storage_data_f_2__48_),
	.ck(clk),
	.d(n10238));
   ms00f80 south_input_NIB_storage_data_f_reg_2__49_ (.o(south_input_NIB_storage_data_f_2__49_),
	.ck(clk),
	.d(n10233));
   ms00f80 south_input_NIB_storage_data_f_reg_2__50_ (.o(south_input_NIB_storage_data_f_2__50_),
	.ck(clk),
	.d(n10228));
   ms00f80 south_input_NIB_storage_data_f_reg_2__51_ (.o(south_input_NIB_storage_data_f_2__51_),
	.ck(clk),
	.d(n10223));
   ms00f80 south_input_NIB_storage_data_f_reg_2__52_ (.o(south_input_NIB_storage_data_f_2__52_),
	.ck(clk),
	.d(n10218));
   ms00f80 south_input_NIB_storage_data_f_reg_2__53_ (.o(south_input_NIB_storage_data_f_2__53_),
	.ck(clk),
	.d(n10213));
   ms00f80 south_input_NIB_storage_data_f_reg_2__54_ (.o(south_input_NIB_storage_data_f_2__54_),
	.ck(clk),
	.d(n10208));
   ms00f80 south_input_NIB_storage_data_f_reg_2__55_ (.o(south_input_NIB_storage_data_f_2__55_),
	.ck(clk),
	.d(n10203));
   ms00f80 south_input_NIB_storage_data_f_reg_2__56_ (.o(south_input_NIB_storage_data_f_2__56_),
	.ck(clk),
	.d(n10198));
   ms00f80 south_input_NIB_storage_data_f_reg_2__57_ (.o(south_input_NIB_storage_data_f_2__57_),
	.ck(clk),
	.d(n10193));
   ms00f80 south_input_NIB_storage_data_f_reg_2__58_ (.o(south_input_NIB_storage_data_f_2__58_),
	.ck(clk),
	.d(n10188));
   ms00f80 south_input_NIB_storage_data_f_reg_2__59_ (.o(south_input_NIB_storage_data_f_2__59_),
	.ck(clk),
	.d(n10183));
   ms00f80 south_input_NIB_storage_data_f_reg_2__60_ (.o(south_input_NIB_storage_data_f_2__60_),
	.ck(clk),
	.d(n10178));
   ms00f80 south_input_NIB_storage_data_f_reg_2__61_ (.o(south_input_NIB_storage_data_f_2__61_),
	.ck(clk),
	.d(n10173));
   ms00f80 south_input_NIB_storage_data_f_reg_2__62_ (.o(south_input_NIB_storage_data_f_2__62_),
	.ck(clk),
	.d(n10168));
   ms00f80 south_input_NIB_storage_data_f_reg_2__63_ (.o(south_input_NIB_storage_data_f_2__63_),
	.ck(clk),
	.d(n10163));
   ms00f80 south_input_NIB_storage_data_f_reg_1__0_ (.o(south_input_NIB_storage_data_f_1__0_),
	.ck(clk),
	.d(n10158));
   ms00f80 south_input_NIB_storage_data_f_reg_1__1_ (.o(south_input_NIB_storage_data_f_1__1_),
	.ck(clk),
	.d(n10153));
   ms00f80 south_input_NIB_storage_data_f_reg_1__2_ (.o(south_input_NIB_storage_data_f_1__2_),
	.ck(clk),
	.d(n10148));
   ms00f80 south_input_NIB_storage_data_f_reg_1__3_ (.o(south_input_NIB_storage_data_f_1__3_),
	.ck(clk),
	.d(n10143));
   ms00f80 south_input_NIB_storage_data_f_reg_1__4_ (.o(south_input_NIB_storage_data_f_1__4_),
	.ck(clk),
	.d(n10138));
   ms00f80 south_input_NIB_storage_data_f_reg_1__5_ (.o(south_input_NIB_storage_data_f_1__5_),
	.ck(clk),
	.d(n10133));
   ms00f80 south_input_NIB_storage_data_f_reg_1__6_ (.o(south_input_NIB_storage_data_f_1__6_),
	.ck(clk),
	.d(n10128));
   ms00f80 south_input_NIB_storage_data_f_reg_1__7_ (.o(south_input_NIB_storage_data_f_1__7_),
	.ck(clk),
	.d(n10123));
   ms00f80 south_input_NIB_storage_data_f_reg_1__8_ (.o(south_input_NIB_storage_data_f_1__8_),
	.ck(clk),
	.d(n10118));
   ms00f80 south_input_NIB_storage_data_f_reg_1__9_ (.o(south_input_NIB_storage_data_f_1__9_),
	.ck(clk),
	.d(n10113));
   ms00f80 south_input_NIB_storage_data_f_reg_1__10_ (.o(south_input_NIB_storage_data_f_1__10_),
	.ck(clk),
	.d(n10108));
   ms00f80 south_input_NIB_storage_data_f_reg_1__11_ (.o(south_input_NIB_storage_data_f_1__11_),
	.ck(clk),
	.d(n10103));
   ms00f80 south_input_NIB_storage_data_f_reg_1__12_ (.o(south_input_NIB_storage_data_f_1__12_),
	.ck(clk),
	.d(n10098));
   ms00f80 south_input_NIB_storage_data_f_reg_1__13_ (.o(south_input_NIB_storage_data_f_1__13_),
	.ck(clk),
	.d(n10093));
   ms00f80 south_input_NIB_storage_data_f_reg_1__14_ (.o(south_input_NIB_storage_data_f_1__14_),
	.ck(clk),
	.d(n10088));
   ms00f80 south_input_NIB_storage_data_f_reg_1__15_ (.o(south_input_NIB_storage_data_f_1__15_),
	.ck(clk),
	.d(n10083));
   ms00f80 south_input_NIB_storage_data_f_reg_1__16_ (.o(south_input_NIB_storage_data_f_1__16_),
	.ck(clk),
	.d(n10078));
   ms00f80 south_input_NIB_storage_data_f_reg_1__17_ (.o(south_input_NIB_storage_data_f_1__17_),
	.ck(clk),
	.d(n10073));
   ms00f80 south_input_NIB_storage_data_f_reg_1__18_ (.o(south_input_NIB_storage_data_f_1__18_),
	.ck(clk),
	.d(n10068));
   ms00f80 south_input_NIB_storage_data_f_reg_1__19_ (.o(south_input_NIB_storage_data_f_1__19_),
	.ck(clk),
	.d(n10063));
   ms00f80 south_input_NIB_storage_data_f_reg_1__20_ (.o(south_input_NIB_storage_data_f_1__20_),
	.ck(clk),
	.d(n10058));
   ms00f80 south_input_NIB_storage_data_f_reg_1__21_ (.o(south_input_NIB_storage_data_f_1__21_),
	.ck(clk),
	.d(n10053));
   ms00f80 south_input_NIB_storage_data_f_reg_1__22_ (.o(south_input_NIB_storage_data_f_1__22_),
	.ck(clk),
	.d(n10048));
   ms00f80 south_input_NIB_storage_data_f_reg_1__23_ (.o(south_input_NIB_storage_data_f_1__23_),
	.ck(clk),
	.d(n10043));
   ms00f80 south_input_NIB_storage_data_f_reg_1__24_ (.o(south_input_NIB_storage_data_f_1__24_),
	.ck(clk),
	.d(n10038));
   ms00f80 south_input_NIB_storage_data_f_reg_1__25_ (.o(south_input_NIB_storage_data_f_1__25_),
	.ck(clk),
	.d(n10033));
   ms00f80 south_input_NIB_storage_data_f_reg_1__26_ (.o(south_input_NIB_storage_data_f_1__26_),
	.ck(clk),
	.d(n10028));
   ms00f80 south_input_NIB_storage_data_f_reg_1__27_ (.o(south_input_NIB_storage_data_f_1__27_),
	.ck(clk),
	.d(n10023));
   ms00f80 south_input_NIB_storage_data_f_reg_1__28_ (.o(south_input_NIB_storage_data_f_1__28_),
	.ck(clk),
	.d(n10018));
   ms00f80 south_input_NIB_storage_data_f_reg_1__29_ (.o(south_input_NIB_storage_data_f_1__29_),
	.ck(clk),
	.d(n10013));
   ms00f80 south_input_NIB_storage_data_f_reg_1__30_ (.o(south_input_NIB_storage_data_f_1__30_),
	.ck(clk),
	.d(n10008));
   ms00f80 south_input_NIB_storage_data_f_reg_1__31_ (.o(south_input_NIB_storage_data_f_1__31_),
	.ck(clk),
	.d(n10003));
   ms00f80 south_input_NIB_storage_data_f_reg_1__32_ (.o(south_input_NIB_storage_data_f_1__32_),
	.ck(clk),
	.d(n9998));
   ms00f80 south_input_NIB_storage_data_f_reg_1__33_ (.o(south_input_NIB_storage_data_f_1__33_),
	.ck(clk),
	.d(n9993));
   ms00f80 south_input_NIB_storage_data_f_reg_1__34_ (.o(south_input_NIB_storage_data_f_1__34_),
	.ck(clk),
	.d(n9988));
   ms00f80 south_input_NIB_storage_data_f_reg_1__35_ (.o(south_input_NIB_storage_data_f_1__35_),
	.ck(clk),
	.d(n9983));
   ms00f80 south_input_NIB_storage_data_f_reg_1__36_ (.o(south_input_NIB_storage_data_f_1__36_),
	.ck(clk),
	.d(n9978));
   ms00f80 south_input_NIB_storage_data_f_reg_1__37_ (.o(south_input_NIB_storage_data_f_1__37_),
	.ck(clk),
	.d(n9973));
   ms00f80 south_input_NIB_storage_data_f_reg_1__38_ (.o(south_input_NIB_storage_data_f_1__38_),
	.ck(clk),
	.d(n9968));
   ms00f80 south_input_NIB_storage_data_f_reg_1__39_ (.o(south_input_NIB_storage_data_f_1__39_),
	.ck(clk),
	.d(n9963));
   ms00f80 south_input_NIB_storage_data_f_reg_1__40_ (.o(south_input_NIB_storage_data_f_1__40_),
	.ck(clk),
	.d(n9958));
   ms00f80 south_input_NIB_storage_data_f_reg_1__41_ (.o(south_input_NIB_storage_data_f_1__41_),
	.ck(clk),
	.d(n9953));
   ms00f80 south_input_NIB_storage_data_f_reg_1__42_ (.o(south_input_NIB_storage_data_f_1__42_),
	.ck(clk),
	.d(n9948));
   ms00f80 south_input_NIB_storage_data_f_reg_1__43_ (.o(south_input_NIB_storage_data_f_1__43_),
	.ck(clk),
	.d(n9943));
   ms00f80 south_input_NIB_storage_data_f_reg_1__44_ (.o(south_input_NIB_storage_data_f_1__44_),
	.ck(clk),
	.d(n9938));
   ms00f80 south_input_NIB_storage_data_f_reg_1__45_ (.o(south_input_NIB_storage_data_f_1__45_),
	.ck(clk),
	.d(n9933));
   ms00f80 south_input_NIB_storage_data_f_reg_1__46_ (.o(south_input_NIB_storage_data_f_1__46_),
	.ck(clk),
	.d(n9928));
   ms00f80 south_input_NIB_storage_data_f_reg_1__47_ (.o(south_input_NIB_storage_data_f_1__47_),
	.ck(clk),
	.d(n9923));
   ms00f80 south_input_NIB_storage_data_f_reg_1__48_ (.o(south_input_NIB_storage_data_f_1__48_),
	.ck(clk),
	.d(n9918));
   ms00f80 south_input_NIB_storage_data_f_reg_1__49_ (.o(south_input_NIB_storage_data_f_1__49_),
	.ck(clk),
	.d(n9913));
   ms00f80 south_input_NIB_storage_data_f_reg_1__50_ (.o(south_input_NIB_storage_data_f_1__50_),
	.ck(clk),
	.d(n9908));
   ms00f80 south_input_NIB_storage_data_f_reg_1__51_ (.o(south_input_NIB_storage_data_f_1__51_),
	.ck(clk),
	.d(n9903));
   ms00f80 south_input_NIB_storage_data_f_reg_1__52_ (.o(south_input_NIB_storage_data_f_1__52_),
	.ck(clk),
	.d(n9898));
   ms00f80 south_input_NIB_storage_data_f_reg_1__53_ (.o(south_input_NIB_storage_data_f_1__53_),
	.ck(clk),
	.d(n9893));
   ms00f80 south_input_NIB_storage_data_f_reg_1__54_ (.o(south_input_NIB_storage_data_f_1__54_),
	.ck(clk),
	.d(n9888));
   ms00f80 south_input_NIB_storage_data_f_reg_1__55_ (.o(south_input_NIB_storage_data_f_1__55_),
	.ck(clk),
	.d(n9883));
   ms00f80 south_input_NIB_storage_data_f_reg_1__56_ (.o(south_input_NIB_storage_data_f_1__56_),
	.ck(clk),
	.d(n9878));
   ms00f80 south_input_NIB_storage_data_f_reg_1__57_ (.o(south_input_NIB_storage_data_f_1__57_),
	.ck(clk),
	.d(n9873));
   ms00f80 south_input_NIB_storage_data_f_reg_1__58_ (.o(south_input_NIB_storage_data_f_1__58_),
	.ck(clk),
	.d(n9868));
   ms00f80 south_input_NIB_storage_data_f_reg_1__59_ (.o(south_input_NIB_storage_data_f_1__59_),
	.ck(clk),
	.d(n9863));
   ms00f80 south_input_NIB_storage_data_f_reg_1__60_ (.o(south_input_NIB_storage_data_f_1__60_),
	.ck(clk),
	.d(n9858));
   ms00f80 south_input_NIB_storage_data_f_reg_1__61_ (.o(south_input_NIB_storage_data_f_1__61_),
	.ck(clk),
	.d(n9853));
   ms00f80 south_input_NIB_storage_data_f_reg_1__62_ (.o(south_input_NIB_storage_data_f_1__62_),
	.ck(clk),
	.d(n9848));
   ms00f80 south_input_NIB_storage_data_f_reg_1__63_ (.o(south_input_NIB_storage_data_f_1__63_),
	.ck(clk),
	.d(n9843));
   ms00f80 south_input_NIB_storage_data_f_reg_0__0_ (.o(south_input_NIB_storage_data_f_0__0_),
	.ck(clk),
	.d(n9838));
   ms00f80 south_input_NIB_storage_data_f_reg_0__1_ (.o(south_input_NIB_storage_data_f_0__1_),
	.ck(clk),
	.d(n9833));
   ms00f80 south_input_NIB_storage_data_f_reg_0__2_ (.o(south_input_NIB_storage_data_f_0__2_),
	.ck(clk),
	.d(n9828));
   ms00f80 south_input_NIB_storage_data_f_reg_0__3_ (.o(south_input_NIB_storage_data_f_0__3_),
	.ck(clk),
	.d(n9823));
   ms00f80 south_input_NIB_storage_data_f_reg_0__4_ (.o(south_input_NIB_storage_data_f_0__4_),
	.ck(clk),
	.d(n9818));
   ms00f80 south_input_NIB_storage_data_f_reg_0__5_ (.o(south_input_NIB_storage_data_f_0__5_),
	.ck(clk),
	.d(n9813));
   ms00f80 south_input_NIB_storage_data_f_reg_0__6_ (.o(south_input_NIB_storage_data_f_0__6_),
	.ck(clk),
	.d(n9808));
   ms00f80 south_input_NIB_storage_data_f_reg_0__7_ (.o(south_input_NIB_storage_data_f_0__7_),
	.ck(clk),
	.d(n9803));
   ms00f80 south_input_NIB_storage_data_f_reg_0__8_ (.o(south_input_NIB_storage_data_f_0__8_),
	.ck(clk),
	.d(n9798));
   ms00f80 south_input_NIB_storage_data_f_reg_0__9_ (.o(south_input_NIB_storage_data_f_0__9_),
	.ck(clk),
	.d(n9793));
   ms00f80 south_input_NIB_storage_data_f_reg_0__10_ (.o(south_input_NIB_storage_data_f_0__10_),
	.ck(clk),
	.d(n9788));
   ms00f80 south_input_NIB_storage_data_f_reg_0__11_ (.o(south_input_NIB_storage_data_f_0__11_),
	.ck(clk),
	.d(n9783));
   ms00f80 south_input_NIB_storage_data_f_reg_0__12_ (.o(south_input_NIB_storage_data_f_0__12_),
	.ck(clk),
	.d(n9778));
   ms00f80 south_input_NIB_storage_data_f_reg_0__13_ (.o(south_input_NIB_storage_data_f_0__13_),
	.ck(clk),
	.d(n9773));
   ms00f80 south_input_NIB_storage_data_f_reg_0__14_ (.o(south_input_NIB_storage_data_f_0__14_),
	.ck(clk),
	.d(n9768));
   ms00f80 south_input_NIB_storage_data_f_reg_0__15_ (.o(south_input_NIB_storage_data_f_0__15_),
	.ck(clk),
	.d(n9763));
   ms00f80 south_input_NIB_storage_data_f_reg_0__16_ (.o(south_input_NIB_storage_data_f_0__16_),
	.ck(clk),
	.d(n9758));
   ms00f80 south_input_NIB_storage_data_f_reg_0__17_ (.o(south_input_NIB_storage_data_f_0__17_),
	.ck(clk),
	.d(n9753));
   ms00f80 south_input_NIB_storage_data_f_reg_0__18_ (.o(south_input_NIB_storage_data_f_0__18_),
	.ck(clk),
	.d(n9748));
   ms00f80 south_input_NIB_storage_data_f_reg_0__19_ (.o(south_input_NIB_storage_data_f_0__19_),
	.ck(clk),
	.d(n9743));
   ms00f80 south_input_NIB_storage_data_f_reg_0__20_ (.o(south_input_NIB_storage_data_f_0__20_),
	.ck(clk),
	.d(n9738));
   ms00f80 south_input_NIB_storage_data_f_reg_0__21_ (.o(south_input_NIB_storage_data_f_0__21_),
	.ck(clk),
	.d(n9733));
   ms00f80 south_input_NIB_storage_data_f_reg_0__22_ (.o(south_input_NIB_storage_data_f_0__22_),
	.ck(clk),
	.d(n9728));
   ms00f80 south_input_NIB_storage_data_f_reg_0__23_ (.o(south_input_NIB_storage_data_f_0__23_),
	.ck(clk),
	.d(n9723));
   ms00f80 south_input_NIB_storage_data_f_reg_0__24_ (.o(south_input_NIB_storage_data_f_0__24_),
	.ck(clk),
	.d(n9718));
   ms00f80 south_input_NIB_storage_data_f_reg_0__25_ (.o(south_input_NIB_storage_data_f_0__25_),
	.ck(clk),
	.d(n9713));
   ms00f80 south_input_NIB_storage_data_f_reg_0__26_ (.o(south_input_NIB_storage_data_f_0__26_),
	.ck(clk),
	.d(n9708));
   ms00f80 south_input_NIB_storage_data_f_reg_0__27_ (.o(south_input_NIB_storage_data_f_0__27_),
	.ck(clk),
	.d(n9703));
   ms00f80 south_input_NIB_storage_data_f_reg_0__28_ (.o(south_input_NIB_storage_data_f_0__28_),
	.ck(clk),
	.d(n9698));
   ms00f80 south_input_NIB_storage_data_f_reg_0__29_ (.o(south_input_NIB_storage_data_f_0__29_),
	.ck(clk),
	.d(n9693));
   ms00f80 south_input_NIB_storage_data_f_reg_0__30_ (.o(south_input_NIB_storage_data_f_0__30_),
	.ck(clk),
	.d(n9688));
   ms00f80 south_input_NIB_storage_data_f_reg_0__31_ (.o(south_input_NIB_storage_data_f_0__31_),
	.ck(clk),
	.d(n9683));
   ms00f80 south_input_NIB_storage_data_f_reg_0__32_ (.o(south_input_NIB_storage_data_f_0__32_),
	.ck(clk),
	.d(n9678));
   ms00f80 south_input_NIB_storage_data_f_reg_0__33_ (.o(south_input_NIB_storage_data_f_0__33_),
	.ck(clk),
	.d(n9673));
   ms00f80 south_input_NIB_storage_data_f_reg_0__34_ (.o(south_input_NIB_storage_data_f_0__34_),
	.ck(clk),
	.d(n9668));
   ms00f80 south_input_NIB_storage_data_f_reg_0__35_ (.o(south_input_NIB_storage_data_f_0__35_),
	.ck(clk),
	.d(n9663));
   ms00f80 south_input_NIB_storage_data_f_reg_0__36_ (.o(south_input_NIB_storage_data_f_0__36_),
	.ck(clk),
	.d(n9658));
   ms00f80 south_input_NIB_storage_data_f_reg_0__37_ (.o(south_input_NIB_storage_data_f_0__37_),
	.ck(clk),
	.d(n9653));
   ms00f80 south_input_NIB_storage_data_f_reg_0__38_ (.o(south_input_NIB_storage_data_f_0__38_),
	.ck(clk),
	.d(n9648));
   ms00f80 south_input_NIB_storage_data_f_reg_0__39_ (.o(south_input_NIB_storage_data_f_0__39_),
	.ck(clk),
	.d(n9643));
   ms00f80 south_input_NIB_storage_data_f_reg_0__40_ (.o(south_input_NIB_storage_data_f_0__40_),
	.ck(clk),
	.d(n9638));
   ms00f80 south_input_NIB_storage_data_f_reg_0__41_ (.o(south_input_NIB_storage_data_f_0__41_),
	.ck(clk),
	.d(n9633));
   ms00f80 south_input_NIB_storage_data_f_reg_0__42_ (.o(south_input_NIB_storage_data_f_0__42_),
	.ck(clk),
	.d(n9628));
   ms00f80 south_input_NIB_storage_data_f_reg_0__43_ (.o(south_input_NIB_storage_data_f_0__43_),
	.ck(clk),
	.d(n9623));
   ms00f80 south_input_NIB_storage_data_f_reg_0__44_ (.o(south_input_NIB_storage_data_f_0__44_),
	.ck(clk),
	.d(n9618));
   ms00f80 south_input_NIB_storage_data_f_reg_0__45_ (.o(south_input_NIB_storage_data_f_0__45_),
	.ck(clk),
	.d(n9613));
   ms00f80 south_input_NIB_storage_data_f_reg_0__46_ (.o(south_input_NIB_storage_data_f_0__46_),
	.ck(clk),
	.d(n9608));
   ms00f80 south_input_NIB_storage_data_f_reg_0__47_ (.o(south_input_NIB_storage_data_f_0__47_),
	.ck(clk),
	.d(n9603));
   ms00f80 south_input_NIB_storage_data_f_reg_0__48_ (.o(south_input_NIB_storage_data_f_0__48_),
	.ck(clk),
	.d(n9598));
   ms00f80 south_input_NIB_storage_data_f_reg_0__49_ (.o(south_input_NIB_storage_data_f_0__49_),
	.ck(clk),
	.d(n9593));
   ms00f80 south_input_NIB_storage_data_f_reg_0__50_ (.o(south_input_NIB_storage_data_f_0__50_),
	.ck(clk),
	.d(n9588));
   ms00f80 south_input_NIB_storage_data_f_reg_0__51_ (.o(south_input_NIB_storage_data_f_0__51_),
	.ck(clk),
	.d(n9583));
   ms00f80 south_input_NIB_storage_data_f_reg_0__52_ (.o(south_input_NIB_storage_data_f_0__52_),
	.ck(clk),
	.d(n9578));
   ms00f80 south_input_NIB_storage_data_f_reg_0__53_ (.o(south_input_NIB_storage_data_f_0__53_),
	.ck(clk),
	.d(n9573));
   ms00f80 south_input_NIB_storage_data_f_reg_0__54_ (.o(south_input_NIB_storage_data_f_0__54_),
	.ck(clk),
	.d(n9568));
   ms00f80 south_input_NIB_storage_data_f_reg_0__55_ (.o(south_input_NIB_storage_data_f_0__55_),
	.ck(clk),
	.d(n9563));
   ms00f80 south_input_NIB_storage_data_f_reg_0__56_ (.o(south_input_NIB_storage_data_f_0__56_),
	.ck(clk),
	.d(n9558));
   ms00f80 south_input_NIB_storage_data_f_reg_0__57_ (.o(south_input_NIB_storage_data_f_0__57_),
	.ck(clk),
	.d(n9553));
   ms00f80 south_input_NIB_storage_data_f_reg_0__58_ (.o(south_input_NIB_storage_data_f_0__58_),
	.ck(clk),
	.d(n9548));
   ms00f80 south_input_NIB_storage_data_f_reg_0__59_ (.o(south_input_NIB_storage_data_f_0__59_),
	.ck(clk),
	.d(n9543));
   ms00f80 south_input_NIB_storage_data_f_reg_0__60_ (.o(south_input_NIB_storage_data_f_0__60_),
	.ck(clk),
	.d(n9538));
   ms00f80 south_input_NIB_storage_data_f_reg_0__61_ (.o(south_input_NIB_storage_data_f_0__61_),
	.ck(clk),
	.d(n9533));
   ms00f80 south_input_NIB_storage_data_f_reg_0__62_ (.o(south_input_NIB_storage_data_f_0__62_),
	.ck(clk),
	.d(n9528));
   ms00f80 south_input_NIB_storage_data_f_reg_0__63_ (.o(south_input_NIB_storage_data_f_0__63_),
	.ck(clk),
	.d(n9523));
   ms00f80 west_input_NIB_tail_ptr_f_reg_0_ (.o(west_input_NIB_tail_ptr_f_0_),
	.ck(clk),
	.d(n9518));
   ms00f80 west_input_NIB_tail_ptr_f_reg_1_ (.o(west_input_NIB_tail_ptr_f_1_),
	.ck(clk),
	.d(n9513));
   ms00f80 west_input_NIB_storage_data_f_reg_3__0_ (.o(west_input_NIB_storage_data_f_3__0_),
	.ck(clk),
	.d(n9508));
   ms00f80 west_input_NIB_storage_data_f_reg_3__1_ (.o(west_input_NIB_storage_data_f_3__1_),
	.ck(clk),
	.d(n9503));
   ms00f80 west_input_NIB_storage_data_f_reg_3__2_ (.o(west_input_NIB_storage_data_f_3__2_),
	.ck(clk),
	.d(n9498));
   ms00f80 west_input_NIB_storage_data_f_reg_3__3_ (.o(west_input_NIB_storage_data_f_3__3_),
	.ck(clk),
	.d(n9493));
   ms00f80 west_input_NIB_storage_data_f_reg_3__4_ (.o(west_input_NIB_storage_data_f_3__4_),
	.ck(clk),
	.d(n9488));
   ms00f80 west_input_NIB_storage_data_f_reg_3__5_ (.o(west_input_NIB_storage_data_f_3__5_),
	.ck(clk),
	.d(n9483));
   ms00f80 west_input_NIB_storage_data_f_reg_3__6_ (.o(west_input_NIB_storage_data_f_3__6_),
	.ck(clk),
	.d(n9478));
   ms00f80 west_input_NIB_storage_data_f_reg_3__7_ (.o(west_input_NIB_storage_data_f_3__7_),
	.ck(clk),
	.d(n9473));
   ms00f80 west_input_NIB_storage_data_f_reg_3__8_ (.o(west_input_NIB_storage_data_f_3__8_),
	.ck(clk),
	.d(n9468));
   ms00f80 west_input_NIB_storage_data_f_reg_3__9_ (.o(west_input_NIB_storage_data_f_3__9_),
	.ck(clk),
	.d(n9463));
   ms00f80 west_input_NIB_storage_data_f_reg_3__10_ (.o(west_input_NIB_storage_data_f_3__10_),
	.ck(clk),
	.d(n9458));
   ms00f80 west_input_NIB_storage_data_f_reg_3__11_ (.o(west_input_NIB_storage_data_f_3__11_),
	.ck(clk),
	.d(n9453));
   ms00f80 west_input_NIB_storage_data_f_reg_3__12_ (.o(west_input_NIB_storage_data_f_3__12_),
	.ck(clk),
	.d(n9448));
   ms00f80 west_input_NIB_storage_data_f_reg_3__13_ (.o(west_input_NIB_storage_data_f_3__13_),
	.ck(clk),
	.d(n9443));
   ms00f80 west_input_NIB_storage_data_f_reg_3__14_ (.o(west_input_NIB_storage_data_f_3__14_),
	.ck(clk),
	.d(n9438));
   ms00f80 west_input_NIB_storage_data_f_reg_3__15_ (.o(west_input_NIB_storage_data_f_3__15_),
	.ck(clk),
	.d(n9433));
   ms00f80 west_input_NIB_storage_data_f_reg_3__16_ (.o(west_input_NIB_storage_data_f_3__16_),
	.ck(clk),
	.d(n9428));
   ms00f80 west_input_NIB_storage_data_f_reg_3__17_ (.o(west_input_NIB_storage_data_f_3__17_),
	.ck(clk),
	.d(n9423));
   ms00f80 west_input_NIB_storage_data_f_reg_3__18_ (.o(west_input_NIB_storage_data_f_3__18_),
	.ck(clk),
	.d(n9418));
   ms00f80 west_input_NIB_storage_data_f_reg_3__19_ (.o(west_input_NIB_storage_data_f_3__19_),
	.ck(clk),
	.d(n9413));
   ms00f80 west_input_NIB_storage_data_f_reg_3__20_ (.o(west_input_NIB_storage_data_f_3__20_),
	.ck(clk),
	.d(n9408));
   ms00f80 west_input_NIB_storage_data_f_reg_3__21_ (.o(west_input_NIB_storage_data_f_3__21_),
	.ck(clk),
	.d(n9403));
   ms00f80 west_input_NIB_storage_data_f_reg_3__22_ (.o(west_input_NIB_storage_data_f_3__22_),
	.ck(clk),
	.d(n9398));
   ms00f80 west_input_NIB_storage_data_f_reg_3__23_ (.o(west_input_NIB_storage_data_f_3__23_),
	.ck(clk),
	.d(n9393));
   ms00f80 west_input_NIB_storage_data_f_reg_3__24_ (.o(west_input_NIB_storage_data_f_3__24_),
	.ck(clk),
	.d(n9388));
   ms00f80 west_input_NIB_storage_data_f_reg_3__25_ (.o(west_input_NIB_storage_data_f_3__25_),
	.ck(clk),
	.d(n9383));
   ms00f80 west_input_NIB_storage_data_f_reg_3__26_ (.o(west_input_NIB_storage_data_f_3__26_),
	.ck(clk),
	.d(n9378));
   ms00f80 west_input_NIB_storage_data_f_reg_3__27_ (.o(west_input_NIB_storage_data_f_3__27_),
	.ck(clk),
	.d(n9373));
   ms00f80 west_input_NIB_storage_data_f_reg_3__28_ (.o(west_input_NIB_storage_data_f_3__28_),
	.ck(clk),
	.d(n9368));
   ms00f80 west_input_NIB_storage_data_f_reg_3__29_ (.o(west_input_NIB_storage_data_f_3__29_),
	.ck(clk),
	.d(n9363));
   ms00f80 west_input_NIB_storage_data_f_reg_3__30_ (.o(west_input_NIB_storage_data_f_3__30_),
	.ck(clk),
	.d(n9358));
   ms00f80 west_input_NIB_storage_data_f_reg_3__31_ (.o(west_input_NIB_storage_data_f_3__31_),
	.ck(clk),
	.d(n9353));
   ms00f80 west_input_NIB_storage_data_f_reg_3__32_ (.o(west_input_NIB_storage_data_f_3__32_),
	.ck(clk),
	.d(n9348));
   ms00f80 west_input_NIB_storage_data_f_reg_3__33_ (.o(west_input_NIB_storage_data_f_3__33_),
	.ck(clk),
	.d(n9343));
   ms00f80 west_input_NIB_storage_data_f_reg_3__34_ (.o(west_input_NIB_storage_data_f_3__34_),
	.ck(clk),
	.d(n9338));
   ms00f80 west_input_NIB_storage_data_f_reg_3__35_ (.o(west_input_NIB_storage_data_f_3__35_),
	.ck(clk),
	.d(n9333));
   ms00f80 west_input_NIB_storage_data_f_reg_3__36_ (.o(west_input_NIB_storage_data_f_3__36_),
	.ck(clk),
	.d(n9328));
   ms00f80 west_input_NIB_storage_data_f_reg_3__37_ (.o(west_input_NIB_storage_data_f_3__37_),
	.ck(clk),
	.d(n9323));
   ms00f80 west_input_NIB_storage_data_f_reg_3__38_ (.o(west_input_NIB_storage_data_f_3__38_),
	.ck(clk),
	.d(n9318));
   ms00f80 west_input_NIB_storage_data_f_reg_3__39_ (.o(west_input_NIB_storage_data_f_3__39_),
	.ck(clk),
	.d(n9313));
   ms00f80 west_input_NIB_storage_data_f_reg_3__40_ (.o(west_input_NIB_storage_data_f_3__40_),
	.ck(clk),
	.d(n9308));
   ms00f80 west_input_NIB_storage_data_f_reg_3__41_ (.o(west_input_NIB_storage_data_f_3__41_),
	.ck(clk),
	.d(n9303));
   ms00f80 west_input_NIB_storage_data_f_reg_3__42_ (.o(west_input_NIB_storage_data_f_3__42_),
	.ck(clk),
	.d(n9298));
   ms00f80 west_input_NIB_storage_data_f_reg_3__43_ (.o(west_input_NIB_storage_data_f_3__43_),
	.ck(clk),
	.d(n9293));
   ms00f80 west_input_NIB_storage_data_f_reg_3__44_ (.o(west_input_NIB_storage_data_f_3__44_),
	.ck(clk),
	.d(n9288));
   ms00f80 west_input_NIB_storage_data_f_reg_3__45_ (.o(west_input_NIB_storage_data_f_3__45_),
	.ck(clk),
	.d(n9283));
   ms00f80 west_input_NIB_storage_data_f_reg_3__46_ (.o(west_input_NIB_storage_data_f_3__46_),
	.ck(clk),
	.d(n9278));
   ms00f80 west_input_NIB_storage_data_f_reg_3__47_ (.o(west_input_NIB_storage_data_f_3__47_),
	.ck(clk),
	.d(n9273));
   ms00f80 west_input_NIB_storage_data_f_reg_3__48_ (.o(west_input_NIB_storage_data_f_3__48_),
	.ck(clk),
	.d(n9268));
   ms00f80 west_input_NIB_storage_data_f_reg_3__49_ (.o(west_input_NIB_storage_data_f_3__49_),
	.ck(clk),
	.d(n9263));
   ms00f80 west_input_NIB_storage_data_f_reg_3__50_ (.o(west_input_NIB_storage_data_f_3__50_),
	.ck(clk),
	.d(n9258));
   ms00f80 west_input_NIB_storage_data_f_reg_3__51_ (.o(west_input_NIB_storage_data_f_3__51_),
	.ck(clk),
	.d(n9253));
   ms00f80 west_input_NIB_storage_data_f_reg_3__52_ (.o(west_input_NIB_storage_data_f_3__52_),
	.ck(clk),
	.d(n9248));
   ms00f80 west_input_NIB_storage_data_f_reg_3__53_ (.o(west_input_NIB_storage_data_f_3__53_),
	.ck(clk),
	.d(n9243));
   ms00f80 west_input_NIB_storage_data_f_reg_3__54_ (.o(west_input_NIB_storage_data_f_3__54_),
	.ck(clk),
	.d(n9238));
   ms00f80 west_input_NIB_storage_data_f_reg_3__55_ (.o(west_input_NIB_storage_data_f_3__55_),
	.ck(clk),
	.d(n9233));
   ms00f80 west_input_NIB_storage_data_f_reg_3__56_ (.o(west_input_NIB_storage_data_f_3__56_),
	.ck(clk),
	.d(n9228));
   ms00f80 west_input_NIB_storage_data_f_reg_3__57_ (.o(west_input_NIB_storage_data_f_3__57_),
	.ck(clk),
	.d(n9223));
   ms00f80 west_input_NIB_storage_data_f_reg_3__58_ (.o(west_input_NIB_storage_data_f_3__58_),
	.ck(clk),
	.d(n9218));
   ms00f80 west_input_NIB_storage_data_f_reg_3__59_ (.o(west_input_NIB_storage_data_f_3__59_),
	.ck(clk),
	.d(n9213));
   ms00f80 west_input_NIB_storage_data_f_reg_3__60_ (.o(west_input_NIB_storage_data_f_3__60_),
	.ck(clk),
	.d(n9208));
   ms00f80 west_input_NIB_storage_data_f_reg_3__61_ (.o(west_input_NIB_storage_data_f_3__61_),
	.ck(clk),
	.d(n9203));
   ms00f80 west_input_NIB_storage_data_f_reg_3__62_ (.o(west_input_NIB_storage_data_f_3__62_),
	.ck(clk),
	.d(n9198));
   ms00f80 west_input_NIB_storage_data_f_reg_3__63_ (.o(west_input_NIB_storage_data_f_3__63_),
	.ck(clk),
	.d(n9193));
   ms00f80 west_input_NIB_storage_data_f_reg_2__0_ (.o(west_input_NIB_storage_data_f_2__0_),
	.ck(clk),
	.d(n9188));
   ms00f80 west_input_NIB_storage_data_f_reg_2__1_ (.o(west_input_NIB_storage_data_f_2__1_),
	.ck(clk),
	.d(n9183));
   ms00f80 west_input_NIB_storage_data_f_reg_2__2_ (.o(west_input_NIB_storage_data_f_2__2_),
	.ck(clk),
	.d(n9178));
   ms00f80 west_input_NIB_storage_data_f_reg_2__3_ (.o(west_input_NIB_storage_data_f_2__3_),
	.ck(clk),
	.d(n9173));
   ms00f80 west_input_NIB_storage_data_f_reg_2__4_ (.o(west_input_NIB_storage_data_f_2__4_),
	.ck(clk),
	.d(n9168));
   ms00f80 west_input_NIB_storage_data_f_reg_2__5_ (.o(west_input_NIB_storage_data_f_2__5_),
	.ck(clk),
	.d(n9163));
   ms00f80 west_input_NIB_storage_data_f_reg_2__6_ (.o(west_input_NIB_storage_data_f_2__6_),
	.ck(clk),
	.d(n9158));
   ms00f80 west_input_NIB_storage_data_f_reg_2__7_ (.o(west_input_NIB_storage_data_f_2__7_),
	.ck(clk),
	.d(n9153));
   ms00f80 west_input_NIB_storage_data_f_reg_2__8_ (.o(west_input_NIB_storage_data_f_2__8_),
	.ck(clk),
	.d(n9148));
   ms00f80 west_input_NIB_storage_data_f_reg_2__9_ (.o(west_input_NIB_storage_data_f_2__9_),
	.ck(clk),
	.d(n9143));
   ms00f80 west_input_NIB_storage_data_f_reg_2__10_ (.o(west_input_NIB_storage_data_f_2__10_),
	.ck(clk),
	.d(n9138));
   ms00f80 west_input_NIB_storage_data_f_reg_2__11_ (.o(west_input_NIB_storage_data_f_2__11_),
	.ck(clk),
	.d(n9133));
   ms00f80 west_input_NIB_storage_data_f_reg_2__12_ (.o(west_input_NIB_storage_data_f_2__12_),
	.ck(clk),
	.d(n9128));
   ms00f80 west_input_NIB_storage_data_f_reg_2__13_ (.o(west_input_NIB_storage_data_f_2__13_),
	.ck(clk),
	.d(n9123));
   ms00f80 west_input_NIB_storage_data_f_reg_2__14_ (.o(west_input_NIB_storage_data_f_2__14_),
	.ck(clk),
	.d(n9118));
   ms00f80 west_input_NIB_storage_data_f_reg_2__15_ (.o(west_input_NIB_storage_data_f_2__15_),
	.ck(clk),
	.d(n9113));
   ms00f80 west_input_NIB_storage_data_f_reg_2__16_ (.o(west_input_NIB_storage_data_f_2__16_),
	.ck(clk),
	.d(n9108));
   ms00f80 west_input_NIB_storage_data_f_reg_2__17_ (.o(west_input_NIB_storage_data_f_2__17_),
	.ck(clk),
	.d(n9103));
   ms00f80 west_input_NIB_storage_data_f_reg_2__18_ (.o(west_input_NIB_storage_data_f_2__18_),
	.ck(clk),
	.d(n9098));
   ms00f80 west_input_NIB_storage_data_f_reg_2__19_ (.o(west_input_NIB_storage_data_f_2__19_),
	.ck(clk),
	.d(n9093));
   ms00f80 west_input_NIB_storage_data_f_reg_2__20_ (.o(west_input_NIB_storage_data_f_2__20_),
	.ck(clk),
	.d(n9088));
   ms00f80 west_input_NIB_storage_data_f_reg_2__21_ (.o(west_input_NIB_storage_data_f_2__21_),
	.ck(clk),
	.d(n9083));
   ms00f80 west_input_NIB_storage_data_f_reg_2__22_ (.o(west_input_NIB_storage_data_f_2__22_),
	.ck(clk),
	.d(n9078));
   ms00f80 west_input_NIB_storage_data_f_reg_2__23_ (.o(west_input_NIB_storage_data_f_2__23_),
	.ck(clk),
	.d(n9073));
   ms00f80 west_input_NIB_storage_data_f_reg_2__24_ (.o(west_input_NIB_storage_data_f_2__24_),
	.ck(clk),
	.d(n9068));
   ms00f80 west_input_NIB_storage_data_f_reg_2__25_ (.o(west_input_NIB_storage_data_f_2__25_),
	.ck(clk),
	.d(n9063));
   ms00f80 west_input_NIB_storage_data_f_reg_2__26_ (.o(west_input_NIB_storage_data_f_2__26_),
	.ck(clk),
	.d(n9058));
   ms00f80 west_input_NIB_storage_data_f_reg_2__27_ (.o(west_input_NIB_storage_data_f_2__27_),
	.ck(clk),
	.d(n9053));
   ms00f80 west_input_NIB_storage_data_f_reg_2__28_ (.o(west_input_NIB_storage_data_f_2__28_),
	.ck(clk),
	.d(n9048));
   ms00f80 west_input_NIB_storage_data_f_reg_2__29_ (.o(west_input_NIB_storage_data_f_2__29_),
	.ck(clk),
	.d(n9043));
   ms00f80 west_input_NIB_storage_data_f_reg_2__30_ (.o(west_input_NIB_storage_data_f_2__30_),
	.ck(clk),
	.d(n9038));
   ms00f80 west_input_NIB_storage_data_f_reg_2__31_ (.o(west_input_NIB_storage_data_f_2__31_),
	.ck(clk),
	.d(n9033));
   ms00f80 west_input_NIB_storage_data_f_reg_2__32_ (.o(west_input_NIB_storage_data_f_2__32_),
	.ck(clk),
	.d(n9028));
   ms00f80 west_input_NIB_storage_data_f_reg_2__33_ (.o(west_input_NIB_storage_data_f_2__33_),
	.ck(clk),
	.d(n9023));
   ms00f80 west_input_NIB_storage_data_f_reg_2__34_ (.o(west_input_NIB_storage_data_f_2__34_),
	.ck(clk),
	.d(n9018));
   ms00f80 west_input_NIB_storage_data_f_reg_2__35_ (.o(west_input_NIB_storage_data_f_2__35_),
	.ck(clk),
	.d(n9013));
   ms00f80 west_input_NIB_storage_data_f_reg_2__36_ (.o(west_input_NIB_storage_data_f_2__36_),
	.ck(clk),
	.d(n9008));
   ms00f80 west_input_NIB_storage_data_f_reg_2__37_ (.o(west_input_NIB_storage_data_f_2__37_),
	.ck(clk),
	.d(n9003));
   ms00f80 west_input_NIB_storage_data_f_reg_2__38_ (.o(west_input_NIB_storage_data_f_2__38_),
	.ck(clk),
	.d(n8998));
   ms00f80 west_input_NIB_storage_data_f_reg_2__39_ (.o(west_input_NIB_storage_data_f_2__39_),
	.ck(clk),
	.d(n8993));
   ms00f80 west_input_NIB_storage_data_f_reg_2__40_ (.o(west_input_NIB_storage_data_f_2__40_),
	.ck(clk),
	.d(n8988));
   ms00f80 west_input_NIB_storage_data_f_reg_2__41_ (.o(west_input_NIB_storage_data_f_2__41_),
	.ck(clk),
	.d(n8983));
   ms00f80 west_input_NIB_storage_data_f_reg_2__42_ (.o(west_input_NIB_storage_data_f_2__42_),
	.ck(clk),
	.d(n8978));
   ms00f80 west_input_NIB_storage_data_f_reg_2__43_ (.o(west_input_NIB_storage_data_f_2__43_),
	.ck(clk),
	.d(n8973));
   ms00f80 west_input_NIB_storage_data_f_reg_2__44_ (.o(west_input_NIB_storage_data_f_2__44_),
	.ck(clk),
	.d(n8968));
   ms00f80 west_input_NIB_storage_data_f_reg_2__45_ (.o(west_input_NIB_storage_data_f_2__45_),
	.ck(clk),
	.d(n8963));
   ms00f80 west_input_NIB_storage_data_f_reg_2__46_ (.o(west_input_NIB_storage_data_f_2__46_),
	.ck(clk),
	.d(n8958));
   ms00f80 west_input_NIB_storage_data_f_reg_2__47_ (.o(west_input_NIB_storage_data_f_2__47_),
	.ck(clk),
	.d(n8953));
   ms00f80 west_input_NIB_storage_data_f_reg_2__48_ (.o(west_input_NIB_storage_data_f_2__48_),
	.ck(clk),
	.d(n8948));
   ms00f80 west_input_NIB_storage_data_f_reg_2__49_ (.o(west_input_NIB_storage_data_f_2__49_),
	.ck(clk),
	.d(n8943));
   ms00f80 west_input_NIB_storage_data_f_reg_2__50_ (.o(west_input_NIB_storage_data_f_2__50_),
	.ck(clk),
	.d(n8938));
   ms00f80 west_input_NIB_storage_data_f_reg_2__51_ (.o(west_input_NIB_storage_data_f_2__51_),
	.ck(clk),
	.d(n8933));
   ms00f80 west_input_NIB_storage_data_f_reg_2__52_ (.o(west_input_NIB_storage_data_f_2__52_),
	.ck(clk),
	.d(n8928));
   ms00f80 west_input_NIB_storage_data_f_reg_2__53_ (.o(west_input_NIB_storage_data_f_2__53_),
	.ck(clk),
	.d(n8923));
   ms00f80 west_input_NIB_storage_data_f_reg_2__54_ (.o(west_input_NIB_storage_data_f_2__54_),
	.ck(clk),
	.d(n8918));
   ms00f80 west_input_NIB_storage_data_f_reg_2__55_ (.o(west_input_NIB_storage_data_f_2__55_),
	.ck(clk),
	.d(n8913));
   ms00f80 west_input_NIB_storage_data_f_reg_2__56_ (.o(west_input_NIB_storage_data_f_2__56_),
	.ck(clk),
	.d(n8908));
   ms00f80 west_input_NIB_storage_data_f_reg_2__57_ (.o(west_input_NIB_storage_data_f_2__57_),
	.ck(clk),
	.d(n8903));
   ms00f80 west_input_NIB_storage_data_f_reg_2__58_ (.o(west_input_NIB_storage_data_f_2__58_),
	.ck(clk),
	.d(n8898));
   ms00f80 west_input_NIB_storage_data_f_reg_2__59_ (.o(west_input_NIB_storage_data_f_2__59_),
	.ck(clk),
	.d(n8893));
   ms00f80 west_input_NIB_storage_data_f_reg_2__60_ (.o(west_input_NIB_storage_data_f_2__60_),
	.ck(clk),
	.d(n8888));
   ms00f80 west_input_NIB_storage_data_f_reg_2__61_ (.o(west_input_NIB_storage_data_f_2__61_),
	.ck(clk),
	.d(n8883));
   ms00f80 west_input_NIB_storage_data_f_reg_2__62_ (.o(west_input_NIB_storage_data_f_2__62_),
	.ck(clk),
	.d(n8878));
   ms00f80 west_input_NIB_storage_data_f_reg_2__63_ (.o(west_input_NIB_storage_data_f_2__63_),
	.ck(clk),
	.d(n8873));
   ms00f80 west_input_NIB_storage_data_f_reg_1__0_ (.o(west_input_NIB_storage_data_f_1__0_),
	.ck(clk),
	.d(n8868));
   ms00f80 west_input_NIB_storage_data_f_reg_1__1_ (.o(west_input_NIB_storage_data_f_1__1_),
	.ck(clk),
	.d(n8863));
   ms00f80 west_input_NIB_storage_data_f_reg_1__2_ (.o(west_input_NIB_storage_data_f_1__2_),
	.ck(clk),
	.d(n8858));
   ms00f80 west_input_NIB_storage_data_f_reg_1__3_ (.o(west_input_NIB_storage_data_f_1__3_),
	.ck(clk),
	.d(n8853));
   ms00f80 west_input_NIB_storage_data_f_reg_1__4_ (.o(west_input_NIB_storage_data_f_1__4_),
	.ck(clk),
	.d(n8848));
   ms00f80 west_input_NIB_storage_data_f_reg_1__5_ (.o(west_input_NIB_storage_data_f_1__5_),
	.ck(clk),
	.d(n8843));
   ms00f80 west_input_NIB_storage_data_f_reg_1__6_ (.o(west_input_NIB_storage_data_f_1__6_),
	.ck(clk),
	.d(n8838));
   ms00f80 west_input_NIB_storage_data_f_reg_1__7_ (.o(west_input_NIB_storage_data_f_1__7_),
	.ck(clk),
	.d(n8833));
   ms00f80 west_input_NIB_storage_data_f_reg_1__8_ (.o(west_input_NIB_storage_data_f_1__8_),
	.ck(clk),
	.d(n8828));
   ms00f80 west_input_NIB_storage_data_f_reg_1__9_ (.o(west_input_NIB_storage_data_f_1__9_),
	.ck(clk),
	.d(n8823));
   ms00f80 west_input_NIB_storage_data_f_reg_1__10_ (.o(west_input_NIB_storage_data_f_1__10_),
	.ck(clk),
	.d(n8818));
   ms00f80 west_input_NIB_storage_data_f_reg_1__11_ (.o(west_input_NIB_storage_data_f_1__11_),
	.ck(clk),
	.d(n8813));
   ms00f80 west_input_NIB_storage_data_f_reg_1__12_ (.o(west_input_NIB_storage_data_f_1__12_),
	.ck(clk),
	.d(n8808));
   ms00f80 west_input_NIB_storage_data_f_reg_1__13_ (.o(west_input_NIB_storage_data_f_1__13_),
	.ck(clk),
	.d(n8803));
   ms00f80 west_input_NIB_storage_data_f_reg_1__14_ (.o(west_input_NIB_storage_data_f_1__14_),
	.ck(clk),
	.d(n8798));
   ms00f80 west_input_NIB_storage_data_f_reg_1__15_ (.o(west_input_NIB_storage_data_f_1__15_),
	.ck(clk),
	.d(n8793));
   ms00f80 west_input_NIB_storage_data_f_reg_1__16_ (.o(west_input_NIB_storage_data_f_1__16_),
	.ck(clk),
	.d(n8788));
   ms00f80 west_input_NIB_storage_data_f_reg_1__17_ (.o(west_input_NIB_storage_data_f_1__17_),
	.ck(clk),
	.d(n8783));
   ms00f80 west_input_NIB_storage_data_f_reg_1__18_ (.o(west_input_NIB_storage_data_f_1__18_),
	.ck(clk),
	.d(n8778));
   ms00f80 west_input_NIB_storage_data_f_reg_1__19_ (.o(west_input_NIB_storage_data_f_1__19_),
	.ck(clk),
	.d(n8773));
   ms00f80 west_input_NIB_storage_data_f_reg_1__20_ (.o(west_input_NIB_storage_data_f_1__20_),
	.ck(clk),
	.d(n8768));
   ms00f80 west_input_NIB_storage_data_f_reg_1__21_ (.o(west_input_NIB_storage_data_f_1__21_),
	.ck(clk),
	.d(n8763));
   ms00f80 west_input_NIB_storage_data_f_reg_1__22_ (.o(west_input_NIB_storage_data_f_1__22_),
	.ck(clk),
	.d(n8758));
   ms00f80 west_input_NIB_storage_data_f_reg_1__23_ (.o(west_input_NIB_storage_data_f_1__23_),
	.ck(clk),
	.d(n8753));
   ms00f80 west_input_NIB_storage_data_f_reg_1__24_ (.o(west_input_NIB_storage_data_f_1__24_),
	.ck(clk),
	.d(n8748));
   ms00f80 west_input_NIB_storage_data_f_reg_1__25_ (.o(west_input_NIB_storage_data_f_1__25_),
	.ck(clk),
	.d(n8743));
   ms00f80 west_input_NIB_storage_data_f_reg_1__26_ (.o(west_input_NIB_storage_data_f_1__26_),
	.ck(clk),
	.d(n8738));
   ms00f80 west_input_NIB_storage_data_f_reg_1__27_ (.o(west_input_NIB_storage_data_f_1__27_),
	.ck(clk),
	.d(n8733));
   ms00f80 west_input_NIB_storage_data_f_reg_1__28_ (.o(west_input_NIB_storage_data_f_1__28_),
	.ck(clk),
	.d(n8728));
   ms00f80 west_input_NIB_storage_data_f_reg_1__29_ (.o(west_input_NIB_storage_data_f_1__29_),
	.ck(clk),
	.d(n8723));
   ms00f80 west_input_NIB_storage_data_f_reg_1__30_ (.o(west_input_NIB_storage_data_f_1__30_),
	.ck(clk),
	.d(n8718));
   ms00f80 west_input_NIB_storage_data_f_reg_1__31_ (.o(west_input_NIB_storage_data_f_1__31_),
	.ck(clk),
	.d(n8713));
   ms00f80 west_input_NIB_storage_data_f_reg_1__32_ (.o(west_input_NIB_storage_data_f_1__32_),
	.ck(clk),
	.d(n8708));
   ms00f80 west_input_NIB_storage_data_f_reg_1__33_ (.o(west_input_NIB_storage_data_f_1__33_),
	.ck(clk),
	.d(n8703));
   ms00f80 west_input_NIB_storage_data_f_reg_1__34_ (.o(west_input_NIB_storage_data_f_1__34_),
	.ck(clk),
	.d(n8698));
   ms00f80 west_input_NIB_storage_data_f_reg_1__35_ (.o(west_input_NIB_storage_data_f_1__35_),
	.ck(clk),
	.d(n8693));
   ms00f80 west_input_NIB_storage_data_f_reg_1__36_ (.o(west_input_NIB_storage_data_f_1__36_),
	.ck(clk),
	.d(n8688));
   ms00f80 west_input_NIB_storage_data_f_reg_1__37_ (.o(west_input_NIB_storage_data_f_1__37_),
	.ck(clk),
	.d(n8683));
   ms00f80 west_input_NIB_storage_data_f_reg_1__38_ (.o(west_input_NIB_storage_data_f_1__38_),
	.ck(clk),
	.d(n8678));
   ms00f80 west_input_NIB_storage_data_f_reg_1__39_ (.o(west_input_NIB_storage_data_f_1__39_),
	.ck(clk),
	.d(n8673));
   ms00f80 west_input_NIB_storage_data_f_reg_1__40_ (.o(west_input_NIB_storage_data_f_1__40_),
	.ck(clk),
	.d(n8668));
   ms00f80 west_input_NIB_storage_data_f_reg_1__41_ (.o(west_input_NIB_storage_data_f_1__41_),
	.ck(clk),
	.d(n8663));
   ms00f80 west_input_NIB_storage_data_f_reg_1__42_ (.o(west_input_NIB_storage_data_f_1__42_),
	.ck(clk),
	.d(n8658));
   ms00f80 west_input_NIB_storage_data_f_reg_1__43_ (.o(west_input_NIB_storage_data_f_1__43_),
	.ck(clk),
	.d(n8653));
   ms00f80 west_input_NIB_storage_data_f_reg_1__44_ (.o(west_input_NIB_storage_data_f_1__44_),
	.ck(clk),
	.d(n8648));
   ms00f80 west_input_NIB_storage_data_f_reg_1__45_ (.o(west_input_NIB_storage_data_f_1__45_),
	.ck(clk),
	.d(n8643));
   ms00f80 west_input_NIB_storage_data_f_reg_1__46_ (.o(west_input_NIB_storage_data_f_1__46_),
	.ck(clk),
	.d(n8638));
   ms00f80 west_input_NIB_storage_data_f_reg_1__47_ (.o(west_input_NIB_storage_data_f_1__47_),
	.ck(clk),
	.d(n8633));
   ms00f80 west_input_NIB_storage_data_f_reg_1__48_ (.o(west_input_NIB_storage_data_f_1__48_),
	.ck(clk),
	.d(n8628));
   ms00f80 west_input_NIB_storage_data_f_reg_1__49_ (.o(west_input_NIB_storage_data_f_1__49_),
	.ck(clk),
	.d(n8623));
   ms00f80 west_input_NIB_storage_data_f_reg_1__50_ (.o(west_input_NIB_storage_data_f_1__50_),
	.ck(clk),
	.d(n8618));
   ms00f80 west_input_NIB_storage_data_f_reg_1__51_ (.o(west_input_NIB_storage_data_f_1__51_),
	.ck(clk),
	.d(n8613));
   ms00f80 west_input_NIB_storage_data_f_reg_1__52_ (.o(west_input_NIB_storage_data_f_1__52_),
	.ck(clk),
	.d(n8608));
   ms00f80 west_input_NIB_storage_data_f_reg_1__53_ (.o(west_input_NIB_storage_data_f_1__53_),
	.ck(clk),
	.d(n8603));
   ms00f80 west_input_NIB_storage_data_f_reg_1__54_ (.o(west_input_NIB_storage_data_f_1__54_),
	.ck(clk),
	.d(n8598));
   ms00f80 west_input_NIB_storage_data_f_reg_1__55_ (.o(west_input_NIB_storage_data_f_1__55_),
	.ck(clk),
	.d(n8593));
   ms00f80 west_input_NIB_storage_data_f_reg_1__56_ (.o(west_input_NIB_storage_data_f_1__56_),
	.ck(clk),
	.d(n8588));
   ms00f80 west_input_NIB_storage_data_f_reg_1__57_ (.o(west_input_NIB_storage_data_f_1__57_),
	.ck(clk),
	.d(n8583));
   ms00f80 west_input_NIB_storage_data_f_reg_1__58_ (.o(west_input_NIB_storage_data_f_1__58_),
	.ck(clk),
	.d(n8578));
   ms00f80 west_input_NIB_storage_data_f_reg_1__59_ (.o(west_input_NIB_storage_data_f_1__59_),
	.ck(clk),
	.d(n8573));
   ms00f80 west_input_NIB_storage_data_f_reg_1__60_ (.o(west_input_NIB_storage_data_f_1__60_),
	.ck(clk),
	.d(n8568));
   ms00f80 west_input_NIB_storage_data_f_reg_1__61_ (.o(west_input_NIB_storage_data_f_1__61_),
	.ck(clk),
	.d(n8563));
   ms00f80 west_input_NIB_storage_data_f_reg_1__62_ (.o(west_input_NIB_storage_data_f_1__62_),
	.ck(clk),
	.d(n8558));
   ms00f80 west_input_NIB_storage_data_f_reg_1__63_ (.o(west_input_NIB_storage_data_f_1__63_),
	.ck(clk),
	.d(n8553));
   ms00f80 west_input_NIB_storage_data_f_reg_0__0_ (.o(west_input_NIB_storage_data_f_0__0_),
	.ck(clk),
	.d(n8548));
   ms00f80 west_input_NIB_storage_data_f_reg_0__1_ (.o(west_input_NIB_storage_data_f_0__1_),
	.ck(clk),
	.d(n8543));
   ms00f80 west_input_NIB_storage_data_f_reg_0__2_ (.o(west_input_NIB_storage_data_f_0__2_),
	.ck(clk),
	.d(n8538));
   ms00f80 west_input_NIB_storage_data_f_reg_0__3_ (.o(west_input_NIB_storage_data_f_0__3_),
	.ck(clk),
	.d(n8533));
   ms00f80 west_input_NIB_storage_data_f_reg_0__4_ (.o(west_input_NIB_storage_data_f_0__4_),
	.ck(clk),
	.d(n8528));
   ms00f80 west_input_NIB_storage_data_f_reg_0__5_ (.o(west_input_NIB_storage_data_f_0__5_),
	.ck(clk),
	.d(n8523));
   ms00f80 west_input_NIB_storage_data_f_reg_0__6_ (.o(west_input_NIB_storage_data_f_0__6_),
	.ck(clk),
	.d(n8518));
   ms00f80 west_input_NIB_storage_data_f_reg_0__7_ (.o(west_input_NIB_storage_data_f_0__7_),
	.ck(clk),
	.d(n8513));
   ms00f80 west_input_NIB_storage_data_f_reg_0__8_ (.o(west_input_NIB_storage_data_f_0__8_),
	.ck(clk),
	.d(n8508));
   ms00f80 west_input_NIB_storage_data_f_reg_0__9_ (.o(west_input_NIB_storage_data_f_0__9_),
	.ck(clk),
	.d(n8503));
   ms00f80 west_input_NIB_storage_data_f_reg_0__10_ (.o(west_input_NIB_storage_data_f_0__10_),
	.ck(clk),
	.d(n8498));
   ms00f80 west_input_NIB_storage_data_f_reg_0__11_ (.o(west_input_NIB_storage_data_f_0__11_),
	.ck(clk),
	.d(n8493));
   ms00f80 west_input_NIB_storage_data_f_reg_0__12_ (.o(west_input_NIB_storage_data_f_0__12_),
	.ck(clk),
	.d(n8488));
   ms00f80 west_input_NIB_storage_data_f_reg_0__13_ (.o(west_input_NIB_storage_data_f_0__13_),
	.ck(clk),
	.d(n8483));
   ms00f80 west_input_NIB_storage_data_f_reg_0__14_ (.o(west_input_NIB_storage_data_f_0__14_),
	.ck(clk),
	.d(n8478));
   ms00f80 west_input_NIB_storage_data_f_reg_0__15_ (.o(west_input_NIB_storage_data_f_0__15_),
	.ck(clk),
	.d(n8473));
   ms00f80 west_input_NIB_storage_data_f_reg_0__16_ (.o(west_input_NIB_storage_data_f_0__16_),
	.ck(clk),
	.d(n8468));
   ms00f80 west_input_NIB_storage_data_f_reg_0__17_ (.o(west_input_NIB_storage_data_f_0__17_),
	.ck(clk),
	.d(n8463));
   ms00f80 west_input_NIB_storage_data_f_reg_0__18_ (.o(west_input_NIB_storage_data_f_0__18_),
	.ck(clk),
	.d(n8458));
   ms00f80 west_input_NIB_storage_data_f_reg_0__19_ (.o(west_input_NIB_storage_data_f_0__19_),
	.ck(clk),
	.d(n8453));
   ms00f80 west_input_NIB_storage_data_f_reg_0__20_ (.o(west_input_NIB_storage_data_f_0__20_),
	.ck(clk),
	.d(n8448));
   ms00f80 west_input_NIB_storage_data_f_reg_0__21_ (.o(west_input_NIB_storage_data_f_0__21_),
	.ck(clk),
	.d(n8443));
   ms00f80 west_input_NIB_storage_data_f_reg_0__22_ (.o(west_input_NIB_storage_data_f_0__22_),
	.ck(clk),
	.d(n8438));
   ms00f80 west_input_NIB_storage_data_f_reg_0__23_ (.o(west_input_NIB_storage_data_f_0__23_),
	.ck(clk),
	.d(n8433));
   ms00f80 west_input_NIB_storage_data_f_reg_0__24_ (.o(west_input_NIB_storage_data_f_0__24_),
	.ck(clk),
	.d(n8428));
   ms00f80 west_input_NIB_storage_data_f_reg_0__25_ (.o(west_input_NIB_storage_data_f_0__25_),
	.ck(clk),
	.d(n8423));
   ms00f80 west_input_NIB_storage_data_f_reg_0__26_ (.o(west_input_NIB_storage_data_f_0__26_),
	.ck(clk),
	.d(n8418));
   ms00f80 west_input_NIB_storage_data_f_reg_0__27_ (.o(west_input_NIB_storage_data_f_0__27_),
	.ck(clk),
	.d(n8413));
   ms00f80 west_input_NIB_storage_data_f_reg_0__28_ (.o(west_input_NIB_storage_data_f_0__28_),
	.ck(clk),
	.d(n8408));
   ms00f80 west_input_NIB_storage_data_f_reg_0__29_ (.o(west_input_NIB_storage_data_f_0__29_),
	.ck(clk),
	.d(n8403));
   ms00f80 west_input_NIB_storage_data_f_reg_0__30_ (.o(west_input_NIB_storage_data_f_0__30_),
	.ck(clk),
	.d(n8398));
   ms00f80 west_input_NIB_storage_data_f_reg_0__31_ (.o(west_input_NIB_storage_data_f_0__31_),
	.ck(clk),
	.d(n8393));
   ms00f80 west_input_NIB_storage_data_f_reg_0__32_ (.o(west_input_NIB_storage_data_f_0__32_),
	.ck(clk),
	.d(n8388));
   ms00f80 west_input_NIB_storage_data_f_reg_0__33_ (.o(west_input_NIB_storage_data_f_0__33_),
	.ck(clk),
	.d(n8383));
   ms00f80 west_input_NIB_storage_data_f_reg_0__34_ (.o(west_input_NIB_storage_data_f_0__34_),
	.ck(clk),
	.d(n8378));
   ms00f80 west_input_NIB_storage_data_f_reg_0__35_ (.o(west_input_NIB_storage_data_f_0__35_),
	.ck(clk),
	.d(n8373));
   ms00f80 west_input_NIB_storage_data_f_reg_0__36_ (.o(west_input_NIB_storage_data_f_0__36_),
	.ck(clk),
	.d(n8368));
   ms00f80 west_input_NIB_storage_data_f_reg_0__37_ (.o(west_input_NIB_storage_data_f_0__37_),
	.ck(clk),
	.d(n8363));
   ms00f80 west_input_NIB_storage_data_f_reg_0__38_ (.o(west_input_NIB_storage_data_f_0__38_),
	.ck(clk),
	.d(n8358));
   ms00f80 west_input_NIB_storage_data_f_reg_0__39_ (.o(west_input_NIB_storage_data_f_0__39_),
	.ck(clk),
	.d(n8353));
   ms00f80 west_input_NIB_storage_data_f_reg_0__40_ (.o(west_input_NIB_storage_data_f_0__40_),
	.ck(clk),
	.d(n8348));
   ms00f80 west_input_NIB_storage_data_f_reg_0__41_ (.o(west_input_NIB_storage_data_f_0__41_),
	.ck(clk),
	.d(n8343));
   ms00f80 west_input_NIB_storage_data_f_reg_0__42_ (.o(west_input_NIB_storage_data_f_0__42_),
	.ck(clk),
	.d(n8338));
   ms00f80 west_input_NIB_storage_data_f_reg_0__43_ (.o(west_input_NIB_storage_data_f_0__43_),
	.ck(clk),
	.d(n8333));
   ms00f80 west_input_NIB_storage_data_f_reg_0__44_ (.o(west_input_NIB_storage_data_f_0__44_),
	.ck(clk),
	.d(n8328));
   ms00f80 west_input_NIB_storage_data_f_reg_0__45_ (.o(west_input_NIB_storage_data_f_0__45_),
	.ck(clk),
	.d(n8323));
   ms00f80 west_input_NIB_storage_data_f_reg_0__46_ (.o(west_input_NIB_storage_data_f_0__46_),
	.ck(clk),
	.d(n8318));
   ms00f80 west_input_NIB_storage_data_f_reg_0__47_ (.o(west_input_NIB_storage_data_f_0__47_),
	.ck(clk),
	.d(n8313));
   ms00f80 west_input_NIB_storage_data_f_reg_0__48_ (.o(west_input_NIB_storage_data_f_0__48_),
	.ck(clk),
	.d(n8308));
   ms00f80 west_input_NIB_storage_data_f_reg_0__49_ (.o(west_input_NIB_storage_data_f_0__49_),
	.ck(clk),
	.d(n8303));
   ms00f80 west_input_NIB_storage_data_f_reg_0__50_ (.o(west_input_NIB_storage_data_f_0__50_),
	.ck(clk),
	.d(n8298));
   ms00f80 west_input_NIB_storage_data_f_reg_0__51_ (.o(west_input_NIB_storage_data_f_0__51_),
	.ck(clk),
	.d(n8293));
   ms00f80 west_input_NIB_storage_data_f_reg_0__52_ (.o(west_input_NIB_storage_data_f_0__52_),
	.ck(clk),
	.d(n8288));
   ms00f80 west_input_NIB_storage_data_f_reg_0__53_ (.o(west_input_NIB_storage_data_f_0__53_),
	.ck(clk),
	.d(n8283));
   ms00f80 west_input_NIB_storage_data_f_reg_0__54_ (.o(west_input_NIB_storage_data_f_0__54_),
	.ck(clk),
	.d(n8278));
   ms00f80 west_input_NIB_storage_data_f_reg_0__55_ (.o(west_input_NIB_storage_data_f_0__55_),
	.ck(clk),
	.d(n8273));
   ms00f80 west_input_NIB_storage_data_f_reg_0__56_ (.o(west_input_NIB_storage_data_f_0__56_),
	.ck(clk),
	.d(n8268));
   ms00f80 west_input_NIB_storage_data_f_reg_0__57_ (.o(west_input_NIB_storage_data_f_0__57_),
	.ck(clk),
	.d(n8263));
   ms00f80 west_input_NIB_storage_data_f_reg_0__58_ (.o(west_input_NIB_storage_data_f_0__58_),
	.ck(clk),
	.d(n8258));
   ms00f80 west_input_NIB_storage_data_f_reg_0__59_ (.o(west_input_NIB_storage_data_f_0__59_),
	.ck(clk),
	.d(n8253));
   ms00f80 west_input_NIB_storage_data_f_reg_0__60_ (.o(west_input_NIB_storage_data_f_0__60_),
	.ck(clk),
	.d(n8248));
   ms00f80 west_input_NIB_storage_data_f_reg_0__61_ (.o(west_input_NIB_storage_data_f_0__61_),
	.ck(clk),
	.d(n8243));
   ms00f80 west_input_NIB_storage_data_f_reg_0__62_ (.o(west_input_NIB_storage_data_f_0__62_),
	.ck(clk),
	.d(n8238));
   ms00f80 west_input_NIB_storage_data_f_reg_0__63_ (.o(west_input_NIB_storage_data_f_0__63_),
	.ck(clk),
	.d(n8233));
   ms00f80 proc_input_NIB_tail_ptr_f_reg_0_ (.o(proc_input_NIB_tail_ptr_f_0_),
	.ck(clk),
	.d(n8228));
   ms00f80 proc_input_NIB_tail_ptr_f_reg_1_ (.o(proc_input_NIB_tail_ptr_f_1_),
	.ck(clk),
	.d(n8223));
   ms00f80 proc_input_NIB_tail_ptr_f_reg_2_ (.o(proc_input_NIB_tail_ptr_f_2_),
	.ck(clk),
	.d(n8218));
   ms00f80 proc_input_NIB_tail_ptr_f_reg_3_ (.o(proc_input_NIB_tail_ptr_f_3_),
	.ck(clk),
	.d(n8213));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__0_ (.o(proc_input_NIB_storage_data_f_15__0_),
	.ck(clk),
	.d(n8208));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__1_ (.o(proc_input_NIB_storage_data_f_15__1_),
	.ck(clk),
	.d(n8203));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__2_ (.o(proc_input_NIB_storage_data_f_15__2_),
	.ck(clk),
	.d(n8198));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__3_ (.o(proc_input_NIB_storage_data_f_15__3_),
	.ck(clk),
	.d(n8193));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__4_ (.o(proc_input_NIB_storage_data_f_15__4_),
	.ck(clk),
	.d(n8188));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__5_ (.o(proc_input_NIB_storage_data_f_15__5_),
	.ck(clk),
	.d(n8183));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__6_ (.o(proc_input_NIB_storage_data_f_15__6_),
	.ck(clk),
	.d(n8178));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__7_ (.o(proc_input_NIB_storage_data_f_15__7_),
	.ck(clk),
	.d(n8173));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__8_ (.o(proc_input_NIB_storage_data_f_15__8_),
	.ck(clk),
	.d(n8168));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__9_ (.o(proc_input_NIB_storage_data_f_15__9_),
	.ck(clk),
	.d(n8163));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__10_ (.o(proc_input_NIB_storage_data_f_15__10_),
	.ck(clk),
	.d(n8158));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__11_ (.o(proc_input_NIB_storage_data_f_15__11_),
	.ck(clk),
	.d(n8153));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__12_ (.o(proc_input_NIB_storage_data_f_15__12_),
	.ck(clk),
	.d(n8148));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__13_ (.o(proc_input_NIB_storage_data_f_15__13_),
	.ck(clk),
	.d(n8143));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__14_ (.o(proc_input_NIB_storage_data_f_15__14_),
	.ck(clk),
	.d(n8138));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__15_ (.o(proc_input_NIB_storage_data_f_15__15_),
	.ck(clk),
	.d(n8133));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__16_ (.o(proc_input_NIB_storage_data_f_15__16_),
	.ck(clk),
	.d(n8128));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__17_ (.o(proc_input_NIB_storage_data_f_15__17_),
	.ck(clk),
	.d(n8123));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__18_ (.o(proc_input_NIB_storage_data_f_15__18_),
	.ck(clk),
	.d(n8118));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__19_ (.o(proc_input_NIB_storage_data_f_15__19_),
	.ck(clk),
	.d(n8113));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__20_ (.o(proc_input_NIB_storage_data_f_15__20_),
	.ck(clk),
	.d(n8108));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__21_ (.o(proc_input_NIB_storage_data_f_15__21_),
	.ck(clk),
	.d(n8103));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__22_ (.o(proc_input_NIB_storage_data_f_15__22_),
	.ck(clk),
	.d(n8098));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__23_ (.o(proc_input_NIB_storage_data_f_15__23_),
	.ck(clk),
	.d(n8093));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__24_ (.o(proc_input_NIB_storage_data_f_15__24_),
	.ck(clk),
	.d(n8088));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__25_ (.o(proc_input_NIB_storage_data_f_15__25_),
	.ck(clk),
	.d(n8083));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__26_ (.o(proc_input_NIB_storage_data_f_15__26_),
	.ck(clk),
	.d(n8078));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__27_ (.o(proc_input_NIB_storage_data_f_15__27_),
	.ck(clk),
	.d(n8073));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__28_ (.o(proc_input_NIB_storage_data_f_15__28_),
	.ck(clk),
	.d(n8068));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__29_ (.o(proc_input_NIB_storage_data_f_15__29_),
	.ck(clk),
	.d(n8063));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__30_ (.o(proc_input_NIB_storage_data_f_15__30_),
	.ck(clk),
	.d(n8058));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__31_ (.o(proc_input_NIB_storage_data_f_15__31_),
	.ck(clk),
	.d(n8053));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__32_ (.o(proc_input_NIB_storage_data_f_15__32_),
	.ck(clk),
	.d(n8048));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__33_ (.o(proc_input_NIB_storage_data_f_15__33_),
	.ck(clk),
	.d(n8043));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__34_ (.o(proc_input_NIB_storage_data_f_15__34_),
	.ck(clk),
	.d(n8038));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__35_ (.o(proc_input_NIB_storage_data_f_15__35_),
	.ck(clk),
	.d(n8033));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__36_ (.o(proc_input_NIB_storage_data_f_15__36_),
	.ck(clk),
	.d(n8028));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__37_ (.o(proc_input_NIB_storage_data_f_15__37_),
	.ck(clk),
	.d(n8023));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__38_ (.o(proc_input_NIB_storage_data_f_15__38_),
	.ck(clk),
	.d(n8018));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__39_ (.o(proc_input_NIB_storage_data_f_15__39_),
	.ck(clk),
	.d(n8013));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__40_ (.o(proc_input_NIB_storage_data_f_15__40_),
	.ck(clk),
	.d(n8008));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__41_ (.o(proc_input_NIB_storage_data_f_15__41_),
	.ck(clk),
	.d(n8003));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__42_ (.o(proc_input_NIB_storage_data_f_15__42_),
	.ck(clk),
	.d(n7998));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__43_ (.o(proc_input_NIB_storage_data_f_15__43_),
	.ck(clk),
	.d(n7993));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__44_ (.o(proc_input_NIB_storage_data_f_15__44_),
	.ck(clk),
	.d(n7988));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__45_ (.o(proc_input_NIB_storage_data_f_15__45_),
	.ck(clk),
	.d(n7983));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__46_ (.o(proc_input_NIB_storage_data_f_15__46_),
	.ck(clk),
	.d(n7978));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__47_ (.o(proc_input_NIB_storage_data_f_15__47_),
	.ck(clk),
	.d(n7973));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__48_ (.o(proc_input_NIB_storage_data_f_15__48_),
	.ck(clk),
	.d(n7968));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__49_ (.o(proc_input_NIB_storage_data_f_15__49_),
	.ck(clk),
	.d(n7963));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__50_ (.o(proc_input_NIB_storage_data_f_15__50_),
	.ck(clk),
	.d(n7958));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__51_ (.o(proc_input_NIB_storage_data_f_15__51_),
	.ck(clk),
	.d(n7953));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__52_ (.o(proc_input_NIB_storage_data_f_15__52_),
	.ck(clk),
	.d(n7948));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__53_ (.o(proc_input_NIB_storage_data_f_15__53_),
	.ck(clk),
	.d(n7943));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__54_ (.o(proc_input_NIB_storage_data_f_15__54_),
	.ck(clk),
	.d(n7938));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__55_ (.o(proc_input_NIB_storage_data_f_15__55_),
	.ck(clk),
	.d(n7933));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__56_ (.o(proc_input_NIB_storage_data_f_15__56_),
	.ck(clk),
	.d(n7928));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__57_ (.o(proc_input_NIB_storage_data_f_15__57_),
	.ck(clk),
	.d(n7923));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__58_ (.o(proc_input_NIB_storage_data_f_15__58_),
	.ck(clk),
	.d(n7918));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__59_ (.o(proc_input_NIB_storage_data_f_15__59_),
	.ck(clk),
	.d(n7913));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__60_ (.o(proc_input_NIB_storage_data_f_15__60_),
	.ck(clk),
	.d(n7908));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__61_ (.o(proc_input_NIB_storage_data_f_15__61_),
	.ck(clk),
	.d(n7903));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__62_ (.o(proc_input_NIB_storage_data_f_15__62_),
	.ck(clk),
	.d(n7898));
   ms00f80 proc_input_NIB_storage_data_f_reg_15__63_ (.o(proc_input_NIB_storage_data_f_15__63_),
	.ck(clk),
	.d(n7893));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__0_ (.o(proc_input_NIB_storage_data_f_14__0_),
	.ck(clk),
	.d(n7888));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__1_ (.o(proc_input_NIB_storage_data_f_14__1_),
	.ck(clk),
	.d(n7883));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__2_ (.o(proc_input_NIB_storage_data_f_14__2_),
	.ck(clk),
	.d(n7878));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__3_ (.o(proc_input_NIB_storage_data_f_14__3_),
	.ck(clk),
	.d(n7873));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__4_ (.o(proc_input_NIB_storage_data_f_14__4_),
	.ck(clk),
	.d(n7868));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__5_ (.o(proc_input_NIB_storage_data_f_14__5_),
	.ck(clk),
	.d(n7863));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__6_ (.o(proc_input_NIB_storage_data_f_14__6_),
	.ck(clk),
	.d(n7858));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__7_ (.o(proc_input_NIB_storage_data_f_14__7_),
	.ck(clk),
	.d(n7853));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__8_ (.o(proc_input_NIB_storage_data_f_14__8_),
	.ck(clk),
	.d(n7848));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__9_ (.o(proc_input_NIB_storage_data_f_14__9_),
	.ck(clk),
	.d(n7843));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__10_ (.o(proc_input_NIB_storage_data_f_14__10_),
	.ck(clk),
	.d(n7838));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__11_ (.o(proc_input_NIB_storage_data_f_14__11_),
	.ck(clk),
	.d(n7833));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__12_ (.o(proc_input_NIB_storage_data_f_14__12_),
	.ck(clk),
	.d(n7828));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__13_ (.o(proc_input_NIB_storage_data_f_14__13_),
	.ck(clk),
	.d(n7823));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__14_ (.o(proc_input_NIB_storage_data_f_14__14_),
	.ck(clk),
	.d(n7818));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__15_ (.o(proc_input_NIB_storage_data_f_14__15_),
	.ck(clk),
	.d(n7813));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__16_ (.o(proc_input_NIB_storage_data_f_14__16_),
	.ck(clk),
	.d(n7808));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__17_ (.o(proc_input_NIB_storage_data_f_14__17_),
	.ck(clk),
	.d(n7803));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__18_ (.o(proc_input_NIB_storage_data_f_14__18_),
	.ck(clk),
	.d(n7798));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__19_ (.o(proc_input_NIB_storage_data_f_14__19_),
	.ck(clk),
	.d(n7793));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__20_ (.o(proc_input_NIB_storage_data_f_14__20_),
	.ck(clk),
	.d(n7788));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__21_ (.o(proc_input_NIB_storage_data_f_14__21_),
	.ck(clk),
	.d(n7783));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__22_ (.o(proc_input_NIB_storage_data_f_14__22_),
	.ck(clk),
	.d(n7778));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__23_ (.o(proc_input_NIB_storage_data_f_14__23_),
	.ck(clk),
	.d(n7773));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__24_ (.o(proc_input_NIB_storage_data_f_14__24_),
	.ck(clk),
	.d(n7768));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__25_ (.o(proc_input_NIB_storage_data_f_14__25_),
	.ck(clk),
	.d(n7763));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__26_ (.o(proc_input_NIB_storage_data_f_14__26_),
	.ck(clk),
	.d(n7758));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__27_ (.o(proc_input_NIB_storage_data_f_14__27_),
	.ck(clk),
	.d(n7753));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__28_ (.o(proc_input_NIB_storage_data_f_14__28_),
	.ck(clk),
	.d(n7748));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__29_ (.o(proc_input_NIB_storage_data_f_14__29_),
	.ck(clk),
	.d(n7743));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__30_ (.o(proc_input_NIB_storage_data_f_14__30_),
	.ck(clk),
	.d(n7738));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__31_ (.o(proc_input_NIB_storage_data_f_14__31_),
	.ck(clk),
	.d(n7733));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__32_ (.o(proc_input_NIB_storage_data_f_14__32_),
	.ck(clk),
	.d(n7728));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__33_ (.o(proc_input_NIB_storage_data_f_14__33_),
	.ck(clk),
	.d(n7723));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__34_ (.o(proc_input_NIB_storage_data_f_14__34_),
	.ck(clk),
	.d(n7718));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__35_ (.o(proc_input_NIB_storage_data_f_14__35_),
	.ck(clk),
	.d(n7713));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__36_ (.o(proc_input_NIB_storage_data_f_14__36_),
	.ck(clk),
	.d(n7708));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__37_ (.o(proc_input_NIB_storage_data_f_14__37_),
	.ck(clk),
	.d(n7703));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__38_ (.o(proc_input_NIB_storage_data_f_14__38_),
	.ck(clk),
	.d(n7698));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__39_ (.o(proc_input_NIB_storage_data_f_14__39_),
	.ck(clk),
	.d(n7693));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__40_ (.o(proc_input_NIB_storage_data_f_14__40_),
	.ck(clk),
	.d(n7688));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__41_ (.o(proc_input_NIB_storage_data_f_14__41_),
	.ck(clk),
	.d(n7683));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__42_ (.o(proc_input_NIB_storage_data_f_14__42_),
	.ck(clk),
	.d(n7678));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__43_ (.o(proc_input_NIB_storage_data_f_14__43_),
	.ck(clk),
	.d(n7673));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__44_ (.o(proc_input_NIB_storage_data_f_14__44_),
	.ck(clk),
	.d(n7668));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__45_ (.o(proc_input_NIB_storage_data_f_14__45_),
	.ck(clk),
	.d(n7663));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__46_ (.o(proc_input_NIB_storage_data_f_14__46_),
	.ck(clk),
	.d(n7658));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__47_ (.o(proc_input_NIB_storage_data_f_14__47_),
	.ck(clk),
	.d(n7653));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__48_ (.o(proc_input_NIB_storage_data_f_14__48_),
	.ck(clk),
	.d(n7648));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__49_ (.o(proc_input_NIB_storage_data_f_14__49_),
	.ck(clk),
	.d(n7643));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__50_ (.o(proc_input_NIB_storage_data_f_14__50_),
	.ck(clk),
	.d(n7638));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__51_ (.o(proc_input_NIB_storage_data_f_14__51_),
	.ck(clk),
	.d(n7633));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__52_ (.o(proc_input_NIB_storage_data_f_14__52_),
	.ck(clk),
	.d(n7628));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__53_ (.o(proc_input_NIB_storage_data_f_14__53_),
	.ck(clk),
	.d(n7623));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__54_ (.o(proc_input_NIB_storage_data_f_14__54_),
	.ck(clk),
	.d(n7618));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__55_ (.o(proc_input_NIB_storage_data_f_14__55_),
	.ck(clk),
	.d(n7613));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__56_ (.o(proc_input_NIB_storage_data_f_14__56_),
	.ck(clk),
	.d(n7608));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__57_ (.o(proc_input_NIB_storage_data_f_14__57_),
	.ck(clk),
	.d(n7603));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__58_ (.o(proc_input_NIB_storage_data_f_14__58_),
	.ck(clk),
	.d(n7598));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__59_ (.o(proc_input_NIB_storage_data_f_14__59_),
	.ck(clk),
	.d(n7593));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__60_ (.o(proc_input_NIB_storage_data_f_14__60_),
	.ck(clk),
	.d(n7588));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__61_ (.o(proc_input_NIB_storage_data_f_14__61_),
	.ck(clk),
	.d(n7583));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__62_ (.o(proc_input_NIB_storage_data_f_14__62_),
	.ck(clk),
	.d(n7578));
   ms00f80 proc_input_NIB_storage_data_f_reg_14__63_ (.o(proc_input_NIB_storage_data_f_14__63_),
	.ck(clk),
	.d(n7573));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__0_ (.o(proc_input_NIB_storage_data_f_13__0_),
	.ck(clk),
	.d(n7568));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__1_ (.o(proc_input_NIB_storage_data_f_13__1_),
	.ck(clk),
	.d(n7563));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__2_ (.o(proc_input_NIB_storage_data_f_13__2_),
	.ck(clk),
	.d(n7558));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__3_ (.o(proc_input_NIB_storage_data_f_13__3_),
	.ck(clk),
	.d(n7553));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__4_ (.o(proc_input_NIB_storage_data_f_13__4_),
	.ck(clk),
	.d(n7548));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__5_ (.o(proc_input_NIB_storage_data_f_13__5_),
	.ck(clk),
	.d(n7543));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__6_ (.o(proc_input_NIB_storage_data_f_13__6_),
	.ck(clk),
	.d(n7538));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__7_ (.o(proc_input_NIB_storage_data_f_13__7_),
	.ck(clk),
	.d(n7533));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__8_ (.o(proc_input_NIB_storage_data_f_13__8_),
	.ck(clk),
	.d(n7528));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__9_ (.o(proc_input_NIB_storage_data_f_13__9_),
	.ck(clk),
	.d(n7523));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__10_ (.o(proc_input_NIB_storage_data_f_13__10_),
	.ck(clk),
	.d(n7518));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__11_ (.o(proc_input_NIB_storage_data_f_13__11_),
	.ck(clk),
	.d(n7513));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__12_ (.o(proc_input_NIB_storage_data_f_13__12_),
	.ck(clk),
	.d(n7508));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__13_ (.o(proc_input_NIB_storage_data_f_13__13_),
	.ck(clk),
	.d(n7503));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__14_ (.o(proc_input_NIB_storage_data_f_13__14_),
	.ck(clk),
	.d(n7498));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__15_ (.o(proc_input_NIB_storage_data_f_13__15_),
	.ck(clk),
	.d(n7493));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__16_ (.o(proc_input_NIB_storage_data_f_13__16_),
	.ck(clk),
	.d(n7488));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__17_ (.o(proc_input_NIB_storage_data_f_13__17_),
	.ck(clk),
	.d(n7483));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__18_ (.o(proc_input_NIB_storage_data_f_13__18_),
	.ck(clk),
	.d(n7478));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__19_ (.o(proc_input_NIB_storage_data_f_13__19_),
	.ck(clk),
	.d(n7473));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__20_ (.o(proc_input_NIB_storage_data_f_13__20_),
	.ck(clk),
	.d(n7468));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__21_ (.o(proc_input_NIB_storage_data_f_13__21_),
	.ck(clk),
	.d(n7463));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__22_ (.o(proc_input_NIB_storage_data_f_13__22_),
	.ck(clk),
	.d(n7458));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__23_ (.o(proc_input_NIB_storage_data_f_13__23_),
	.ck(clk),
	.d(n7453));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__24_ (.o(proc_input_NIB_storage_data_f_13__24_),
	.ck(clk),
	.d(n7448));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__25_ (.o(proc_input_NIB_storage_data_f_13__25_),
	.ck(clk),
	.d(n7443));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__26_ (.o(proc_input_NIB_storage_data_f_13__26_),
	.ck(clk),
	.d(n7438));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__27_ (.o(proc_input_NIB_storage_data_f_13__27_),
	.ck(clk),
	.d(n7433));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__28_ (.o(proc_input_NIB_storage_data_f_13__28_),
	.ck(clk),
	.d(n7428));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__29_ (.o(proc_input_NIB_storage_data_f_13__29_),
	.ck(clk),
	.d(n7423));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__30_ (.o(proc_input_NIB_storage_data_f_13__30_),
	.ck(clk),
	.d(n7418));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__31_ (.o(proc_input_NIB_storage_data_f_13__31_),
	.ck(clk),
	.d(n7413));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__32_ (.o(proc_input_NIB_storage_data_f_13__32_),
	.ck(clk),
	.d(n7408));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__33_ (.o(proc_input_NIB_storage_data_f_13__33_),
	.ck(clk),
	.d(n7403));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__34_ (.o(proc_input_NIB_storage_data_f_13__34_),
	.ck(clk),
	.d(n7398));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__35_ (.o(proc_input_NIB_storage_data_f_13__35_),
	.ck(clk),
	.d(n7393));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__36_ (.o(proc_input_NIB_storage_data_f_13__36_),
	.ck(clk),
	.d(n7388));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__37_ (.o(proc_input_NIB_storage_data_f_13__37_),
	.ck(clk),
	.d(n7383));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__38_ (.o(proc_input_NIB_storage_data_f_13__38_),
	.ck(clk),
	.d(n7378));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__39_ (.o(proc_input_NIB_storage_data_f_13__39_),
	.ck(clk),
	.d(n7373));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__40_ (.o(proc_input_NIB_storage_data_f_13__40_),
	.ck(clk),
	.d(n7368));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__41_ (.o(proc_input_NIB_storage_data_f_13__41_),
	.ck(clk),
	.d(n7363));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__42_ (.o(proc_input_NIB_storage_data_f_13__42_),
	.ck(clk),
	.d(n7358));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__43_ (.o(proc_input_NIB_storage_data_f_13__43_),
	.ck(clk),
	.d(n7353));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__44_ (.o(proc_input_NIB_storage_data_f_13__44_),
	.ck(clk),
	.d(n7348));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__45_ (.o(proc_input_NIB_storage_data_f_13__45_),
	.ck(clk),
	.d(n7343));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__46_ (.o(proc_input_NIB_storage_data_f_13__46_),
	.ck(clk),
	.d(n7338));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__47_ (.o(proc_input_NIB_storage_data_f_13__47_),
	.ck(clk),
	.d(n7333));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__48_ (.o(proc_input_NIB_storage_data_f_13__48_),
	.ck(clk),
	.d(n7328));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__49_ (.o(proc_input_NIB_storage_data_f_13__49_),
	.ck(clk),
	.d(n7323));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__50_ (.o(proc_input_NIB_storage_data_f_13__50_),
	.ck(clk),
	.d(n7318));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__51_ (.o(proc_input_NIB_storage_data_f_13__51_),
	.ck(clk),
	.d(n7313));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__52_ (.o(proc_input_NIB_storage_data_f_13__52_),
	.ck(clk),
	.d(n7308));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__53_ (.o(proc_input_NIB_storage_data_f_13__53_),
	.ck(clk),
	.d(n7303));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__54_ (.o(proc_input_NIB_storage_data_f_13__54_),
	.ck(clk),
	.d(n7298));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__55_ (.o(proc_input_NIB_storage_data_f_13__55_),
	.ck(clk),
	.d(n7293));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__56_ (.o(proc_input_NIB_storage_data_f_13__56_),
	.ck(clk),
	.d(n7288));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__57_ (.o(proc_input_NIB_storage_data_f_13__57_),
	.ck(clk),
	.d(n7283));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__58_ (.o(proc_input_NIB_storage_data_f_13__58_),
	.ck(clk),
	.d(n7278));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__59_ (.o(proc_input_NIB_storage_data_f_13__59_),
	.ck(clk),
	.d(n7273));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__60_ (.o(proc_input_NIB_storage_data_f_13__60_),
	.ck(clk),
	.d(n7268));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__61_ (.o(proc_input_NIB_storage_data_f_13__61_),
	.ck(clk),
	.d(n7263));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__62_ (.o(proc_input_NIB_storage_data_f_13__62_),
	.ck(clk),
	.d(n7258));
   ms00f80 proc_input_NIB_storage_data_f_reg_13__63_ (.o(proc_input_NIB_storage_data_f_13__63_),
	.ck(clk),
	.d(n7253));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__0_ (.o(proc_input_NIB_storage_data_f_12__0_),
	.ck(clk),
	.d(n7248));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__1_ (.o(proc_input_NIB_storage_data_f_12__1_),
	.ck(clk),
	.d(n7243));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__2_ (.o(proc_input_NIB_storage_data_f_12__2_),
	.ck(clk),
	.d(n7238));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__3_ (.o(proc_input_NIB_storage_data_f_12__3_),
	.ck(clk),
	.d(n7233));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__4_ (.o(proc_input_NIB_storage_data_f_12__4_),
	.ck(clk),
	.d(n7228));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__5_ (.o(proc_input_NIB_storage_data_f_12__5_),
	.ck(clk),
	.d(n7223));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__6_ (.o(proc_input_NIB_storage_data_f_12__6_),
	.ck(clk),
	.d(n7218));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__7_ (.o(proc_input_NIB_storage_data_f_12__7_),
	.ck(clk),
	.d(n7213));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__8_ (.o(proc_input_NIB_storage_data_f_12__8_),
	.ck(clk),
	.d(n7208));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__9_ (.o(proc_input_NIB_storage_data_f_12__9_),
	.ck(clk),
	.d(n7203));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__10_ (.o(proc_input_NIB_storage_data_f_12__10_),
	.ck(clk),
	.d(n7198));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__11_ (.o(proc_input_NIB_storage_data_f_12__11_),
	.ck(clk),
	.d(n7193));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__12_ (.o(proc_input_NIB_storage_data_f_12__12_),
	.ck(clk),
	.d(n7188));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__13_ (.o(proc_input_NIB_storage_data_f_12__13_),
	.ck(clk),
	.d(n7183));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__14_ (.o(proc_input_NIB_storage_data_f_12__14_),
	.ck(clk),
	.d(n7178));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__15_ (.o(proc_input_NIB_storage_data_f_12__15_),
	.ck(clk),
	.d(n7173));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__16_ (.o(proc_input_NIB_storage_data_f_12__16_),
	.ck(clk),
	.d(n7168));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__17_ (.o(proc_input_NIB_storage_data_f_12__17_),
	.ck(clk),
	.d(n7163));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__18_ (.o(proc_input_NIB_storage_data_f_12__18_),
	.ck(clk),
	.d(n7158));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__19_ (.o(proc_input_NIB_storage_data_f_12__19_),
	.ck(clk),
	.d(n7153));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__20_ (.o(proc_input_NIB_storage_data_f_12__20_),
	.ck(clk),
	.d(n7148));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__21_ (.o(proc_input_NIB_storage_data_f_12__21_),
	.ck(clk),
	.d(n7143));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__22_ (.o(proc_input_NIB_storage_data_f_12__22_),
	.ck(clk),
	.d(n7138));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__23_ (.o(proc_input_NIB_storage_data_f_12__23_),
	.ck(clk),
	.d(n7133));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__24_ (.o(proc_input_NIB_storage_data_f_12__24_),
	.ck(clk),
	.d(n7128));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__25_ (.o(proc_input_NIB_storage_data_f_12__25_),
	.ck(clk),
	.d(n7123));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__26_ (.o(proc_input_NIB_storage_data_f_12__26_),
	.ck(clk),
	.d(n7118));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__27_ (.o(proc_input_NIB_storage_data_f_12__27_),
	.ck(clk),
	.d(n7113));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__28_ (.o(proc_input_NIB_storage_data_f_12__28_),
	.ck(clk),
	.d(n7108));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__29_ (.o(proc_input_NIB_storage_data_f_12__29_),
	.ck(clk),
	.d(n7103));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__30_ (.o(proc_input_NIB_storage_data_f_12__30_),
	.ck(clk),
	.d(n7098));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__31_ (.o(proc_input_NIB_storage_data_f_12__31_),
	.ck(clk),
	.d(n7093));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__32_ (.o(proc_input_NIB_storage_data_f_12__32_),
	.ck(clk),
	.d(n7088));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__33_ (.o(proc_input_NIB_storage_data_f_12__33_),
	.ck(clk),
	.d(n7083));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__34_ (.o(proc_input_NIB_storage_data_f_12__34_),
	.ck(clk),
	.d(n7078));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__35_ (.o(proc_input_NIB_storage_data_f_12__35_),
	.ck(clk),
	.d(n7073));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__36_ (.o(proc_input_NIB_storage_data_f_12__36_),
	.ck(clk),
	.d(n7068));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__37_ (.o(proc_input_NIB_storage_data_f_12__37_),
	.ck(clk),
	.d(n7063));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__38_ (.o(proc_input_NIB_storage_data_f_12__38_),
	.ck(clk),
	.d(n7058));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__39_ (.o(proc_input_NIB_storage_data_f_12__39_),
	.ck(clk),
	.d(n7053));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__40_ (.o(proc_input_NIB_storage_data_f_12__40_),
	.ck(clk),
	.d(n7048));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__41_ (.o(proc_input_NIB_storage_data_f_12__41_),
	.ck(clk),
	.d(n7043));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__42_ (.o(proc_input_NIB_storage_data_f_12__42_),
	.ck(clk),
	.d(n7038));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__43_ (.o(proc_input_NIB_storage_data_f_12__43_),
	.ck(clk),
	.d(n7033));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__44_ (.o(proc_input_NIB_storage_data_f_12__44_),
	.ck(clk),
	.d(n7028));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__45_ (.o(proc_input_NIB_storage_data_f_12__45_),
	.ck(clk),
	.d(n7023));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__46_ (.o(proc_input_NIB_storage_data_f_12__46_),
	.ck(clk),
	.d(n7018));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__47_ (.o(proc_input_NIB_storage_data_f_12__47_),
	.ck(clk),
	.d(n7013));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__48_ (.o(proc_input_NIB_storage_data_f_12__48_),
	.ck(clk),
	.d(n7008));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__49_ (.o(proc_input_NIB_storage_data_f_12__49_),
	.ck(clk),
	.d(n7003));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__50_ (.o(proc_input_NIB_storage_data_f_12__50_),
	.ck(clk),
	.d(n6998));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__51_ (.o(proc_input_NIB_storage_data_f_12__51_),
	.ck(clk),
	.d(n6993));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__52_ (.o(proc_input_NIB_storage_data_f_12__52_),
	.ck(clk),
	.d(n6988));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__53_ (.o(proc_input_NIB_storage_data_f_12__53_),
	.ck(clk),
	.d(n6983));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__54_ (.o(proc_input_NIB_storage_data_f_12__54_),
	.ck(clk),
	.d(n6978));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__55_ (.o(proc_input_NIB_storage_data_f_12__55_),
	.ck(clk),
	.d(n6973));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__56_ (.o(proc_input_NIB_storage_data_f_12__56_),
	.ck(clk),
	.d(n6968));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__57_ (.o(proc_input_NIB_storage_data_f_12__57_),
	.ck(clk),
	.d(n6963));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__58_ (.o(proc_input_NIB_storage_data_f_12__58_),
	.ck(clk),
	.d(n6958));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__59_ (.o(proc_input_NIB_storage_data_f_12__59_),
	.ck(clk),
	.d(n6953));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__60_ (.o(proc_input_NIB_storage_data_f_12__60_),
	.ck(clk),
	.d(n6948));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__61_ (.o(proc_input_NIB_storage_data_f_12__61_),
	.ck(clk),
	.d(n6943));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__62_ (.o(proc_input_NIB_storage_data_f_12__62_),
	.ck(clk),
	.d(n6938));
   ms00f80 proc_input_NIB_storage_data_f_reg_12__63_ (.o(proc_input_NIB_storage_data_f_12__63_),
	.ck(clk),
	.d(n6933));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__0_ (.o(proc_input_NIB_storage_data_f_11__0_),
	.ck(clk),
	.d(n6928));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__1_ (.o(proc_input_NIB_storage_data_f_11__1_),
	.ck(clk),
	.d(n6923));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__2_ (.o(proc_input_NIB_storage_data_f_11__2_),
	.ck(clk),
	.d(n6918));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__3_ (.o(proc_input_NIB_storage_data_f_11__3_),
	.ck(clk),
	.d(n6913));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__4_ (.o(proc_input_NIB_storage_data_f_11__4_),
	.ck(clk),
	.d(n6908));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__5_ (.o(proc_input_NIB_storage_data_f_11__5_),
	.ck(clk),
	.d(n6903));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__6_ (.o(proc_input_NIB_storage_data_f_11__6_),
	.ck(clk),
	.d(n6898));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__7_ (.o(proc_input_NIB_storage_data_f_11__7_),
	.ck(clk),
	.d(n6893));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__8_ (.o(proc_input_NIB_storage_data_f_11__8_),
	.ck(clk),
	.d(n6888));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__9_ (.o(proc_input_NIB_storage_data_f_11__9_),
	.ck(clk),
	.d(n6883));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__10_ (.o(proc_input_NIB_storage_data_f_11__10_),
	.ck(clk),
	.d(n6878));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__11_ (.o(proc_input_NIB_storage_data_f_11__11_),
	.ck(clk),
	.d(n6873));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__12_ (.o(proc_input_NIB_storage_data_f_11__12_),
	.ck(clk),
	.d(n6868));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__13_ (.o(proc_input_NIB_storage_data_f_11__13_),
	.ck(clk),
	.d(n6863));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__14_ (.o(proc_input_NIB_storage_data_f_11__14_),
	.ck(clk),
	.d(n6858));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__15_ (.o(proc_input_NIB_storage_data_f_11__15_),
	.ck(clk),
	.d(n6853));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__16_ (.o(proc_input_NIB_storage_data_f_11__16_),
	.ck(clk),
	.d(n6848));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__17_ (.o(proc_input_NIB_storage_data_f_11__17_),
	.ck(clk),
	.d(n6843));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__18_ (.o(proc_input_NIB_storage_data_f_11__18_),
	.ck(clk),
	.d(n6838));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__19_ (.o(proc_input_NIB_storage_data_f_11__19_),
	.ck(clk),
	.d(n6833));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__20_ (.o(proc_input_NIB_storage_data_f_11__20_),
	.ck(clk),
	.d(n6828));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__21_ (.o(proc_input_NIB_storage_data_f_11__21_),
	.ck(clk),
	.d(n6823));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__22_ (.o(proc_input_NIB_storage_data_f_11__22_),
	.ck(clk),
	.d(n6818));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__23_ (.o(proc_input_NIB_storage_data_f_11__23_),
	.ck(clk),
	.d(n6813));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__24_ (.o(proc_input_NIB_storage_data_f_11__24_),
	.ck(clk),
	.d(n6808));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__25_ (.o(proc_input_NIB_storage_data_f_11__25_),
	.ck(clk),
	.d(n6803));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__26_ (.o(proc_input_NIB_storage_data_f_11__26_),
	.ck(clk),
	.d(n6798));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__27_ (.o(proc_input_NIB_storage_data_f_11__27_),
	.ck(clk),
	.d(n6793));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__28_ (.o(proc_input_NIB_storage_data_f_11__28_),
	.ck(clk),
	.d(n6788));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__29_ (.o(proc_input_NIB_storage_data_f_11__29_),
	.ck(clk),
	.d(n6783));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__30_ (.o(proc_input_NIB_storage_data_f_11__30_),
	.ck(clk),
	.d(n6778));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__31_ (.o(proc_input_NIB_storage_data_f_11__31_),
	.ck(clk),
	.d(n6773));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__32_ (.o(proc_input_NIB_storage_data_f_11__32_),
	.ck(clk),
	.d(n6768));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__33_ (.o(proc_input_NIB_storage_data_f_11__33_),
	.ck(clk),
	.d(n6763));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__34_ (.o(proc_input_NIB_storage_data_f_11__34_),
	.ck(clk),
	.d(n6758));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__35_ (.o(proc_input_NIB_storage_data_f_11__35_),
	.ck(clk),
	.d(n6753));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__36_ (.o(proc_input_NIB_storage_data_f_11__36_),
	.ck(clk),
	.d(n6748));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__37_ (.o(proc_input_NIB_storage_data_f_11__37_),
	.ck(clk),
	.d(n6743));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__38_ (.o(proc_input_NIB_storage_data_f_11__38_),
	.ck(clk),
	.d(n6738));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__39_ (.o(proc_input_NIB_storage_data_f_11__39_),
	.ck(clk),
	.d(n6733));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__40_ (.o(proc_input_NIB_storage_data_f_11__40_),
	.ck(clk),
	.d(n6728));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__41_ (.o(proc_input_NIB_storage_data_f_11__41_),
	.ck(clk),
	.d(n6723));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__42_ (.o(proc_input_NIB_storage_data_f_11__42_),
	.ck(clk),
	.d(n6718));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__43_ (.o(proc_input_NIB_storage_data_f_11__43_),
	.ck(clk),
	.d(n6713));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__44_ (.o(proc_input_NIB_storage_data_f_11__44_),
	.ck(clk),
	.d(n6708));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__45_ (.o(proc_input_NIB_storage_data_f_11__45_),
	.ck(clk),
	.d(n6703));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__46_ (.o(proc_input_NIB_storage_data_f_11__46_),
	.ck(clk),
	.d(n6698));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__47_ (.o(proc_input_NIB_storage_data_f_11__47_),
	.ck(clk),
	.d(n6693));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__48_ (.o(proc_input_NIB_storage_data_f_11__48_),
	.ck(clk),
	.d(n6688));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__49_ (.o(proc_input_NIB_storage_data_f_11__49_),
	.ck(clk),
	.d(n6683));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__50_ (.o(proc_input_NIB_storage_data_f_11__50_),
	.ck(clk),
	.d(n6678));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__51_ (.o(proc_input_NIB_storage_data_f_11__51_),
	.ck(clk),
	.d(n6673));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__52_ (.o(proc_input_NIB_storage_data_f_11__52_),
	.ck(clk),
	.d(n6668));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__53_ (.o(proc_input_NIB_storage_data_f_11__53_),
	.ck(clk),
	.d(n6663));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__54_ (.o(proc_input_NIB_storage_data_f_11__54_),
	.ck(clk),
	.d(n6658));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__55_ (.o(proc_input_NIB_storage_data_f_11__55_),
	.ck(clk),
	.d(n6653));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__56_ (.o(proc_input_NIB_storage_data_f_11__56_),
	.ck(clk),
	.d(n6648));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__57_ (.o(proc_input_NIB_storage_data_f_11__57_),
	.ck(clk),
	.d(n6643));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__58_ (.o(proc_input_NIB_storage_data_f_11__58_),
	.ck(clk),
	.d(n6638));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__59_ (.o(proc_input_NIB_storage_data_f_11__59_),
	.ck(clk),
	.d(n6633));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__60_ (.o(proc_input_NIB_storage_data_f_11__60_),
	.ck(clk),
	.d(n6628));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__61_ (.o(proc_input_NIB_storage_data_f_11__61_),
	.ck(clk),
	.d(n6623));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__62_ (.o(proc_input_NIB_storage_data_f_11__62_),
	.ck(clk),
	.d(n6618));
   ms00f80 proc_input_NIB_storage_data_f_reg_11__63_ (.o(proc_input_NIB_storage_data_f_11__63_),
	.ck(clk),
	.d(n6613));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__0_ (.o(proc_input_NIB_storage_data_f_10__0_),
	.ck(clk),
	.d(n6608));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__1_ (.o(proc_input_NIB_storage_data_f_10__1_),
	.ck(clk),
	.d(n6603));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__2_ (.o(proc_input_NIB_storage_data_f_10__2_),
	.ck(clk),
	.d(n6598));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__3_ (.o(proc_input_NIB_storage_data_f_10__3_),
	.ck(clk),
	.d(n6593));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__4_ (.o(proc_input_NIB_storage_data_f_10__4_),
	.ck(clk),
	.d(n6588));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__5_ (.o(proc_input_NIB_storage_data_f_10__5_),
	.ck(clk),
	.d(n6583));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__6_ (.o(proc_input_NIB_storage_data_f_10__6_),
	.ck(clk),
	.d(n6578));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__7_ (.o(proc_input_NIB_storage_data_f_10__7_),
	.ck(clk),
	.d(n6573));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__8_ (.o(proc_input_NIB_storage_data_f_10__8_),
	.ck(clk),
	.d(n6568));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__9_ (.o(proc_input_NIB_storage_data_f_10__9_),
	.ck(clk),
	.d(n6563));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__10_ (.o(proc_input_NIB_storage_data_f_10__10_),
	.ck(clk),
	.d(n6558));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__11_ (.o(proc_input_NIB_storage_data_f_10__11_),
	.ck(clk),
	.d(n6553));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__12_ (.o(proc_input_NIB_storage_data_f_10__12_),
	.ck(clk),
	.d(n6548));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__13_ (.o(proc_input_NIB_storage_data_f_10__13_),
	.ck(clk),
	.d(n6543));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__14_ (.o(proc_input_NIB_storage_data_f_10__14_),
	.ck(clk),
	.d(n6538));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__15_ (.o(proc_input_NIB_storage_data_f_10__15_),
	.ck(clk),
	.d(n6533));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__16_ (.o(proc_input_NIB_storage_data_f_10__16_),
	.ck(clk),
	.d(n6528));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__17_ (.o(proc_input_NIB_storage_data_f_10__17_),
	.ck(clk),
	.d(n6523));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__18_ (.o(proc_input_NIB_storage_data_f_10__18_),
	.ck(clk),
	.d(n6518));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__19_ (.o(proc_input_NIB_storage_data_f_10__19_),
	.ck(clk),
	.d(n6513));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__20_ (.o(proc_input_NIB_storage_data_f_10__20_),
	.ck(clk),
	.d(n6508));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__21_ (.o(proc_input_NIB_storage_data_f_10__21_),
	.ck(clk),
	.d(n6503));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__22_ (.o(proc_input_NIB_storage_data_f_10__22_),
	.ck(clk),
	.d(n6498));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__23_ (.o(proc_input_NIB_storage_data_f_10__23_),
	.ck(clk),
	.d(n6493));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__24_ (.o(proc_input_NIB_storage_data_f_10__24_),
	.ck(clk),
	.d(n6488));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__25_ (.o(proc_input_NIB_storage_data_f_10__25_),
	.ck(clk),
	.d(n6483));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__26_ (.o(proc_input_NIB_storage_data_f_10__26_),
	.ck(clk),
	.d(n6478));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__27_ (.o(proc_input_NIB_storage_data_f_10__27_),
	.ck(clk),
	.d(n6473));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__28_ (.o(proc_input_NIB_storage_data_f_10__28_),
	.ck(clk),
	.d(n6468));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__29_ (.o(proc_input_NIB_storage_data_f_10__29_),
	.ck(clk),
	.d(n6463));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__30_ (.o(proc_input_NIB_storage_data_f_10__30_),
	.ck(clk),
	.d(n6458));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__31_ (.o(proc_input_NIB_storage_data_f_10__31_),
	.ck(clk),
	.d(n6453));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__32_ (.o(proc_input_NIB_storage_data_f_10__32_),
	.ck(clk),
	.d(n6448));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__33_ (.o(proc_input_NIB_storage_data_f_10__33_),
	.ck(clk),
	.d(n6443));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__34_ (.o(proc_input_NIB_storage_data_f_10__34_),
	.ck(clk),
	.d(n6438));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__35_ (.o(proc_input_NIB_storage_data_f_10__35_),
	.ck(clk),
	.d(n6433));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__36_ (.o(proc_input_NIB_storage_data_f_10__36_),
	.ck(clk),
	.d(n6428));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__37_ (.o(proc_input_NIB_storage_data_f_10__37_),
	.ck(clk),
	.d(n6423));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__38_ (.o(proc_input_NIB_storage_data_f_10__38_),
	.ck(clk),
	.d(n6418));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__39_ (.o(proc_input_NIB_storage_data_f_10__39_),
	.ck(clk),
	.d(n6413));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__40_ (.o(proc_input_NIB_storage_data_f_10__40_),
	.ck(clk),
	.d(n6408));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__41_ (.o(proc_input_NIB_storage_data_f_10__41_),
	.ck(clk),
	.d(n6403));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__42_ (.o(proc_input_NIB_storage_data_f_10__42_),
	.ck(clk),
	.d(n6398));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__43_ (.o(proc_input_NIB_storage_data_f_10__43_),
	.ck(clk),
	.d(n6393));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__44_ (.o(proc_input_NIB_storage_data_f_10__44_),
	.ck(clk),
	.d(n6388));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__45_ (.o(proc_input_NIB_storage_data_f_10__45_),
	.ck(clk),
	.d(n6383));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__46_ (.o(proc_input_NIB_storage_data_f_10__46_),
	.ck(clk),
	.d(n6378));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__47_ (.o(proc_input_NIB_storage_data_f_10__47_),
	.ck(clk),
	.d(n6373));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__48_ (.o(proc_input_NIB_storage_data_f_10__48_),
	.ck(clk),
	.d(n6368));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__49_ (.o(proc_input_NIB_storage_data_f_10__49_),
	.ck(clk),
	.d(n6363));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__50_ (.o(proc_input_NIB_storage_data_f_10__50_),
	.ck(clk),
	.d(n6358));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__51_ (.o(proc_input_NIB_storage_data_f_10__51_),
	.ck(clk),
	.d(n6353));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__52_ (.o(proc_input_NIB_storage_data_f_10__52_),
	.ck(clk),
	.d(n6348));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__53_ (.o(proc_input_NIB_storage_data_f_10__53_),
	.ck(clk),
	.d(n6343));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__54_ (.o(proc_input_NIB_storage_data_f_10__54_),
	.ck(clk),
	.d(n6338));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__55_ (.o(proc_input_NIB_storage_data_f_10__55_),
	.ck(clk),
	.d(n6333));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__56_ (.o(proc_input_NIB_storage_data_f_10__56_),
	.ck(clk),
	.d(n6328));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__57_ (.o(proc_input_NIB_storage_data_f_10__57_),
	.ck(clk),
	.d(n6323));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__58_ (.o(proc_input_NIB_storage_data_f_10__58_),
	.ck(clk),
	.d(n6318));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__59_ (.o(proc_input_NIB_storage_data_f_10__59_),
	.ck(clk),
	.d(n6313));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__60_ (.o(proc_input_NIB_storage_data_f_10__60_),
	.ck(clk),
	.d(n6308));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__61_ (.o(proc_input_NIB_storage_data_f_10__61_),
	.ck(clk),
	.d(n6303));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__62_ (.o(proc_input_NIB_storage_data_f_10__62_),
	.ck(clk),
	.d(n6298));
   ms00f80 proc_input_NIB_storage_data_f_reg_10__63_ (.o(proc_input_NIB_storage_data_f_10__63_),
	.ck(clk),
	.d(n6293));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__0_ (.o(proc_input_NIB_storage_data_f_9__0_),
	.ck(clk),
	.d(n6288));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__1_ (.o(proc_input_NIB_storage_data_f_9__1_),
	.ck(clk),
	.d(n6283));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__2_ (.o(proc_input_NIB_storage_data_f_9__2_),
	.ck(clk),
	.d(n6278));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__3_ (.o(proc_input_NIB_storage_data_f_9__3_),
	.ck(clk),
	.d(n6273));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__4_ (.o(proc_input_NIB_storage_data_f_9__4_),
	.ck(clk),
	.d(n6268));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__5_ (.o(proc_input_NIB_storage_data_f_9__5_),
	.ck(clk),
	.d(n6263));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__6_ (.o(proc_input_NIB_storage_data_f_9__6_),
	.ck(clk),
	.d(n6258));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__7_ (.o(proc_input_NIB_storage_data_f_9__7_),
	.ck(clk),
	.d(n6253));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__8_ (.o(proc_input_NIB_storage_data_f_9__8_),
	.ck(clk),
	.d(n6248));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__9_ (.o(proc_input_NIB_storage_data_f_9__9_),
	.ck(clk),
	.d(n6243));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__10_ (.o(proc_input_NIB_storage_data_f_9__10_),
	.ck(clk),
	.d(n6238));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__11_ (.o(proc_input_NIB_storage_data_f_9__11_),
	.ck(clk),
	.d(n6233));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__12_ (.o(proc_input_NIB_storage_data_f_9__12_),
	.ck(clk),
	.d(n6228));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__13_ (.o(proc_input_NIB_storage_data_f_9__13_),
	.ck(clk),
	.d(n6223));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__14_ (.o(proc_input_NIB_storage_data_f_9__14_),
	.ck(clk),
	.d(n6218));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__15_ (.o(proc_input_NIB_storage_data_f_9__15_),
	.ck(clk),
	.d(n6213));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__16_ (.o(proc_input_NIB_storage_data_f_9__16_),
	.ck(clk),
	.d(n6208));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__17_ (.o(proc_input_NIB_storage_data_f_9__17_),
	.ck(clk),
	.d(n6203));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__18_ (.o(proc_input_NIB_storage_data_f_9__18_),
	.ck(clk),
	.d(n6198));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__19_ (.o(proc_input_NIB_storage_data_f_9__19_),
	.ck(clk),
	.d(n6193));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__20_ (.o(proc_input_NIB_storage_data_f_9__20_),
	.ck(clk),
	.d(n6188));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__21_ (.o(proc_input_NIB_storage_data_f_9__21_),
	.ck(clk),
	.d(n6183));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__22_ (.o(proc_input_NIB_storage_data_f_9__22_),
	.ck(clk),
	.d(n6178));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__23_ (.o(proc_input_NIB_storage_data_f_9__23_),
	.ck(clk),
	.d(n6173));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__24_ (.o(proc_input_NIB_storage_data_f_9__24_),
	.ck(clk),
	.d(n6168));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__25_ (.o(proc_input_NIB_storage_data_f_9__25_),
	.ck(clk),
	.d(n6163));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__26_ (.o(proc_input_NIB_storage_data_f_9__26_),
	.ck(clk),
	.d(n6158));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__27_ (.o(proc_input_NIB_storage_data_f_9__27_),
	.ck(clk),
	.d(n6153));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__28_ (.o(proc_input_NIB_storage_data_f_9__28_),
	.ck(clk),
	.d(n6148));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__29_ (.o(proc_input_NIB_storage_data_f_9__29_),
	.ck(clk),
	.d(n6143));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__30_ (.o(proc_input_NIB_storage_data_f_9__30_),
	.ck(clk),
	.d(n6138));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__31_ (.o(proc_input_NIB_storage_data_f_9__31_),
	.ck(clk),
	.d(n6133));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__32_ (.o(proc_input_NIB_storage_data_f_9__32_),
	.ck(clk),
	.d(n6128));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__33_ (.o(proc_input_NIB_storage_data_f_9__33_),
	.ck(clk),
	.d(n6123));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__34_ (.o(proc_input_NIB_storage_data_f_9__34_),
	.ck(clk),
	.d(n6118));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__35_ (.o(proc_input_NIB_storage_data_f_9__35_),
	.ck(clk),
	.d(n6113));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__36_ (.o(proc_input_NIB_storage_data_f_9__36_),
	.ck(clk),
	.d(n6108));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__37_ (.o(proc_input_NIB_storage_data_f_9__37_),
	.ck(clk),
	.d(n6103));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__38_ (.o(proc_input_NIB_storage_data_f_9__38_),
	.ck(clk),
	.d(n6098));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__39_ (.o(proc_input_NIB_storage_data_f_9__39_),
	.ck(clk),
	.d(n6093));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__40_ (.o(proc_input_NIB_storage_data_f_9__40_),
	.ck(clk),
	.d(n6088));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__41_ (.o(proc_input_NIB_storage_data_f_9__41_),
	.ck(clk),
	.d(n6083));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__42_ (.o(proc_input_NIB_storage_data_f_9__42_),
	.ck(clk),
	.d(n6078));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__43_ (.o(proc_input_NIB_storage_data_f_9__43_),
	.ck(clk),
	.d(n6073));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__44_ (.o(proc_input_NIB_storage_data_f_9__44_),
	.ck(clk),
	.d(n6068));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__45_ (.o(proc_input_NIB_storage_data_f_9__45_),
	.ck(clk),
	.d(n6063));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__46_ (.o(proc_input_NIB_storage_data_f_9__46_),
	.ck(clk),
	.d(n6058));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__47_ (.o(proc_input_NIB_storage_data_f_9__47_),
	.ck(clk),
	.d(n6053));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__48_ (.o(proc_input_NIB_storage_data_f_9__48_),
	.ck(clk),
	.d(n6048));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__49_ (.o(proc_input_NIB_storage_data_f_9__49_),
	.ck(clk),
	.d(n6043));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__50_ (.o(proc_input_NIB_storage_data_f_9__50_),
	.ck(clk),
	.d(n6038));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__51_ (.o(proc_input_NIB_storage_data_f_9__51_),
	.ck(clk),
	.d(n6033));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__52_ (.o(proc_input_NIB_storage_data_f_9__52_),
	.ck(clk),
	.d(n6028));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__53_ (.o(proc_input_NIB_storage_data_f_9__53_),
	.ck(clk),
	.d(n6023));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__54_ (.o(proc_input_NIB_storage_data_f_9__54_),
	.ck(clk),
	.d(n6018));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__55_ (.o(proc_input_NIB_storage_data_f_9__55_),
	.ck(clk),
	.d(n6013));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__56_ (.o(proc_input_NIB_storage_data_f_9__56_),
	.ck(clk),
	.d(n6008));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__57_ (.o(proc_input_NIB_storage_data_f_9__57_),
	.ck(clk),
	.d(n6003));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__58_ (.o(proc_input_NIB_storage_data_f_9__58_),
	.ck(clk),
	.d(n5998));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__59_ (.o(proc_input_NIB_storage_data_f_9__59_),
	.ck(clk),
	.d(n5993));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__60_ (.o(proc_input_NIB_storage_data_f_9__60_),
	.ck(clk),
	.d(n5988));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__61_ (.o(proc_input_NIB_storage_data_f_9__61_),
	.ck(clk),
	.d(n5983));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__62_ (.o(proc_input_NIB_storage_data_f_9__62_),
	.ck(clk),
	.d(n5978));
   ms00f80 proc_input_NIB_storage_data_f_reg_9__63_ (.o(proc_input_NIB_storage_data_f_9__63_),
	.ck(clk),
	.d(n5973));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__0_ (.o(proc_input_NIB_storage_data_f_8__0_),
	.ck(clk),
	.d(n5968));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__1_ (.o(proc_input_NIB_storage_data_f_8__1_),
	.ck(clk),
	.d(n5963));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__2_ (.o(proc_input_NIB_storage_data_f_8__2_),
	.ck(clk),
	.d(n5958));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__3_ (.o(proc_input_NIB_storage_data_f_8__3_),
	.ck(clk),
	.d(n5953));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__4_ (.o(proc_input_NIB_storage_data_f_8__4_),
	.ck(clk),
	.d(n5948));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__5_ (.o(proc_input_NIB_storage_data_f_8__5_),
	.ck(clk),
	.d(n5943));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__6_ (.o(proc_input_NIB_storage_data_f_8__6_),
	.ck(clk),
	.d(n5938));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__7_ (.o(proc_input_NIB_storage_data_f_8__7_),
	.ck(clk),
	.d(n5933));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__8_ (.o(proc_input_NIB_storage_data_f_8__8_),
	.ck(clk),
	.d(n5928));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__9_ (.o(proc_input_NIB_storage_data_f_8__9_),
	.ck(clk),
	.d(n5923));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__10_ (.o(proc_input_NIB_storage_data_f_8__10_),
	.ck(clk),
	.d(n5918));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__11_ (.o(proc_input_NIB_storage_data_f_8__11_),
	.ck(clk),
	.d(n5913));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__12_ (.o(proc_input_NIB_storage_data_f_8__12_),
	.ck(clk),
	.d(n5908));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__13_ (.o(proc_input_NIB_storage_data_f_8__13_),
	.ck(clk),
	.d(n5903));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__14_ (.o(proc_input_NIB_storage_data_f_8__14_),
	.ck(clk),
	.d(n5898));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__15_ (.o(proc_input_NIB_storage_data_f_8__15_),
	.ck(clk),
	.d(n5893));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__16_ (.o(proc_input_NIB_storage_data_f_8__16_),
	.ck(clk),
	.d(n5888));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__17_ (.o(proc_input_NIB_storage_data_f_8__17_),
	.ck(clk),
	.d(n5883));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__18_ (.o(proc_input_NIB_storage_data_f_8__18_),
	.ck(clk),
	.d(n5878));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__19_ (.o(proc_input_NIB_storage_data_f_8__19_),
	.ck(clk),
	.d(n5873));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__20_ (.o(proc_input_NIB_storage_data_f_8__20_),
	.ck(clk),
	.d(n5868));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__21_ (.o(proc_input_NIB_storage_data_f_8__21_),
	.ck(clk),
	.d(n5863));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__22_ (.o(proc_input_NIB_storage_data_f_8__22_),
	.ck(clk),
	.d(n5858));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__23_ (.o(proc_input_NIB_storage_data_f_8__23_),
	.ck(clk),
	.d(n5853));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__24_ (.o(proc_input_NIB_storage_data_f_8__24_),
	.ck(clk),
	.d(n5848));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__25_ (.o(proc_input_NIB_storage_data_f_8__25_),
	.ck(clk),
	.d(n5843));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__26_ (.o(proc_input_NIB_storage_data_f_8__26_),
	.ck(clk),
	.d(n5838));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__27_ (.o(proc_input_NIB_storage_data_f_8__27_),
	.ck(clk),
	.d(n5833));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__28_ (.o(proc_input_NIB_storage_data_f_8__28_),
	.ck(clk),
	.d(n5828));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__29_ (.o(proc_input_NIB_storage_data_f_8__29_),
	.ck(clk),
	.d(n5823));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__30_ (.o(proc_input_NIB_storage_data_f_8__30_),
	.ck(clk),
	.d(n5818));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__31_ (.o(proc_input_NIB_storage_data_f_8__31_),
	.ck(clk),
	.d(n5813));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__32_ (.o(proc_input_NIB_storage_data_f_8__32_),
	.ck(clk),
	.d(n5808));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__33_ (.o(proc_input_NIB_storage_data_f_8__33_),
	.ck(clk),
	.d(n5803));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__34_ (.o(proc_input_NIB_storage_data_f_8__34_),
	.ck(clk),
	.d(n5798));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__35_ (.o(proc_input_NIB_storage_data_f_8__35_),
	.ck(clk),
	.d(n5793));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__36_ (.o(proc_input_NIB_storage_data_f_8__36_),
	.ck(clk),
	.d(n5788));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__37_ (.o(proc_input_NIB_storage_data_f_8__37_),
	.ck(clk),
	.d(n5783));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__38_ (.o(proc_input_NIB_storage_data_f_8__38_),
	.ck(clk),
	.d(n5778));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__39_ (.o(proc_input_NIB_storage_data_f_8__39_),
	.ck(clk),
	.d(n5773));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__40_ (.o(proc_input_NIB_storage_data_f_8__40_),
	.ck(clk),
	.d(n5768));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__41_ (.o(proc_input_NIB_storage_data_f_8__41_),
	.ck(clk),
	.d(n5763));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__42_ (.o(proc_input_NIB_storage_data_f_8__42_),
	.ck(clk),
	.d(n5758));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__43_ (.o(proc_input_NIB_storage_data_f_8__43_),
	.ck(clk),
	.d(n5753));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__44_ (.o(proc_input_NIB_storage_data_f_8__44_),
	.ck(clk),
	.d(n5748));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__45_ (.o(proc_input_NIB_storage_data_f_8__45_),
	.ck(clk),
	.d(n5743));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__46_ (.o(proc_input_NIB_storage_data_f_8__46_),
	.ck(clk),
	.d(n5738));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__47_ (.o(proc_input_NIB_storage_data_f_8__47_),
	.ck(clk),
	.d(n5733));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__48_ (.o(proc_input_NIB_storage_data_f_8__48_),
	.ck(clk),
	.d(n5728));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__49_ (.o(proc_input_NIB_storage_data_f_8__49_),
	.ck(clk),
	.d(n5723));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__50_ (.o(proc_input_NIB_storage_data_f_8__50_),
	.ck(clk),
	.d(n5718));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__51_ (.o(proc_input_NIB_storage_data_f_8__51_),
	.ck(clk),
	.d(n5713));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__52_ (.o(proc_input_NIB_storage_data_f_8__52_),
	.ck(clk),
	.d(n5708));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__53_ (.o(proc_input_NIB_storage_data_f_8__53_),
	.ck(clk),
	.d(n5703));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__54_ (.o(proc_input_NIB_storage_data_f_8__54_),
	.ck(clk),
	.d(n5698));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__55_ (.o(proc_input_NIB_storage_data_f_8__55_),
	.ck(clk),
	.d(n5693));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__56_ (.o(proc_input_NIB_storage_data_f_8__56_),
	.ck(clk),
	.d(n5688));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__57_ (.o(proc_input_NIB_storage_data_f_8__57_),
	.ck(clk),
	.d(n5683));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__58_ (.o(proc_input_NIB_storage_data_f_8__58_),
	.ck(clk),
	.d(n5678));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__59_ (.o(proc_input_NIB_storage_data_f_8__59_),
	.ck(clk),
	.d(n5673));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__60_ (.o(proc_input_NIB_storage_data_f_8__60_),
	.ck(clk),
	.d(n5668));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__61_ (.o(proc_input_NIB_storage_data_f_8__61_),
	.ck(clk),
	.d(n5663));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__62_ (.o(proc_input_NIB_storage_data_f_8__62_),
	.ck(clk),
	.d(n5658));
   ms00f80 proc_input_NIB_storage_data_f_reg_8__63_ (.o(proc_input_NIB_storage_data_f_8__63_),
	.ck(clk),
	.d(n5653));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__0_ (.o(proc_input_NIB_storage_data_f_7__0_),
	.ck(clk),
	.d(n5648));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__1_ (.o(proc_input_NIB_storage_data_f_7__1_),
	.ck(clk),
	.d(n5643));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__2_ (.o(proc_input_NIB_storage_data_f_7__2_),
	.ck(clk),
	.d(n5638));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__3_ (.o(proc_input_NIB_storage_data_f_7__3_),
	.ck(clk),
	.d(n5633));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__4_ (.o(proc_input_NIB_storage_data_f_7__4_),
	.ck(clk),
	.d(n5628));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__5_ (.o(proc_input_NIB_storage_data_f_7__5_),
	.ck(clk),
	.d(n5623));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__6_ (.o(proc_input_NIB_storage_data_f_7__6_),
	.ck(clk),
	.d(n5618));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__7_ (.o(proc_input_NIB_storage_data_f_7__7_),
	.ck(clk),
	.d(n5613));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__8_ (.o(proc_input_NIB_storage_data_f_7__8_),
	.ck(clk),
	.d(n5608));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__9_ (.o(proc_input_NIB_storage_data_f_7__9_),
	.ck(clk),
	.d(n5603));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__10_ (.o(proc_input_NIB_storage_data_f_7__10_),
	.ck(clk),
	.d(n5598));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__11_ (.o(proc_input_NIB_storage_data_f_7__11_),
	.ck(clk),
	.d(n5593));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__12_ (.o(proc_input_NIB_storage_data_f_7__12_),
	.ck(clk),
	.d(n5588));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__13_ (.o(proc_input_NIB_storage_data_f_7__13_),
	.ck(clk),
	.d(n5583));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__14_ (.o(proc_input_NIB_storage_data_f_7__14_),
	.ck(clk),
	.d(n5578));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__15_ (.o(proc_input_NIB_storage_data_f_7__15_),
	.ck(clk),
	.d(n5573));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__16_ (.o(proc_input_NIB_storage_data_f_7__16_),
	.ck(clk),
	.d(n5568));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__17_ (.o(proc_input_NIB_storage_data_f_7__17_),
	.ck(clk),
	.d(n5563));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__18_ (.o(proc_input_NIB_storage_data_f_7__18_),
	.ck(clk),
	.d(n5558));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__19_ (.o(proc_input_NIB_storage_data_f_7__19_),
	.ck(clk),
	.d(n5553));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__20_ (.o(proc_input_NIB_storage_data_f_7__20_),
	.ck(clk),
	.d(n5548));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__21_ (.o(proc_input_NIB_storage_data_f_7__21_),
	.ck(clk),
	.d(n5543));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__22_ (.o(proc_input_NIB_storage_data_f_7__22_),
	.ck(clk),
	.d(n5538));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__23_ (.o(proc_input_NIB_storage_data_f_7__23_),
	.ck(clk),
	.d(n5533));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__24_ (.o(proc_input_NIB_storage_data_f_7__24_),
	.ck(clk),
	.d(n5528));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__25_ (.o(proc_input_NIB_storage_data_f_7__25_),
	.ck(clk),
	.d(n5523));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__26_ (.o(proc_input_NIB_storage_data_f_7__26_),
	.ck(clk),
	.d(n5518));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__27_ (.o(proc_input_NIB_storage_data_f_7__27_),
	.ck(clk),
	.d(n5513));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__28_ (.o(proc_input_NIB_storage_data_f_7__28_),
	.ck(clk),
	.d(n5508));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__29_ (.o(proc_input_NIB_storage_data_f_7__29_),
	.ck(clk),
	.d(n5503));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__30_ (.o(proc_input_NIB_storage_data_f_7__30_),
	.ck(clk),
	.d(n5498));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__31_ (.o(proc_input_NIB_storage_data_f_7__31_),
	.ck(clk),
	.d(n5493));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__32_ (.o(proc_input_NIB_storage_data_f_7__32_),
	.ck(clk),
	.d(n5488));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__33_ (.o(proc_input_NIB_storage_data_f_7__33_),
	.ck(clk),
	.d(n5483));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__34_ (.o(proc_input_NIB_storage_data_f_7__34_),
	.ck(clk),
	.d(n5478));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__35_ (.o(proc_input_NIB_storage_data_f_7__35_),
	.ck(clk),
	.d(n5473));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__36_ (.o(proc_input_NIB_storage_data_f_7__36_),
	.ck(clk),
	.d(n5468));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__37_ (.o(proc_input_NIB_storage_data_f_7__37_),
	.ck(clk),
	.d(n5463));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__38_ (.o(proc_input_NIB_storage_data_f_7__38_),
	.ck(clk),
	.d(n5458));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__39_ (.o(proc_input_NIB_storage_data_f_7__39_),
	.ck(clk),
	.d(n5453));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__40_ (.o(proc_input_NIB_storage_data_f_7__40_),
	.ck(clk),
	.d(n5448));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__41_ (.o(proc_input_NIB_storage_data_f_7__41_),
	.ck(clk),
	.d(n5443));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__42_ (.o(proc_input_NIB_storage_data_f_7__42_),
	.ck(clk),
	.d(n5438));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__43_ (.o(proc_input_NIB_storage_data_f_7__43_),
	.ck(clk),
	.d(n5433));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__44_ (.o(proc_input_NIB_storage_data_f_7__44_),
	.ck(clk),
	.d(n5428));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__45_ (.o(proc_input_NIB_storage_data_f_7__45_),
	.ck(clk),
	.d(n5423));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__46_ (.o(proc_input_NIB_storage_data_f_7__46_),
	.ck(clk),
	.d(n5418));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__47_ (.o(proc_input_NIB_storage_data_f_7__47_),
	.ck(clk),
	.d(n5413));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__48_ (.o(proc_input_NIB_storage_data_f_7__48_),
	.ck(clk),
	.d(n5408));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__49_ (.o(proc_input_NIB_storage_data_f_7__49_),
	.ck(clk),
	.d(n5403));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__50_ (.o(proc_input_NIB_storage_data_f_7__50_),
	.ck(clk),
	.d(n5398));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__51_ (.o(proc_input_NIB_storage_data_f_7__51_),
	.ck(clk),
	.d(n5393));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__52_ (.o(proc_input_NIB_storage_data_f_7__52_),
	.ck(clk),
	.d(n5388));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__53_ (.o(proc_input_NIB_storage_data_f_7__53_),
	.ck(clk),
	.d(n5383));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__54_ (.o(proc_input_NIB_storage_data_f_7__54_),
	.ck(clk),
	.d(n5378));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__55_ (.o(proc_input_NIB_storage_data_f_7__55_),
	.ck(clk),
	.d(n5373));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__56_ (.o(proc_input_NIB_storage_data_f_7__56_),
	.ck(clk),
	.d(n5368));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__57_ (.o(proc_input_NIB_storage_data_f_7__57_),
	.ck(clk),
	.d(n5363));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__58_ (.o(proc_input_NIB_storage_data_f_7__58_),
	.ck(clk),
	.d(n5358));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__59_ (.o(proc_input_NIB_storage_data_f_7__59_),
	.ck(clk),
	.d(n5353));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__60_ (.o(proc_input_NIB_storage_data_f_7__60_),
	.ck(clk),
	.d(n5348));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__61_ (.o(proc_input_NIB_storage_data_f_7__61_),
	.ck(clk),
	.d(n5343));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__62_ (.o(proc_input_NIB_storage_data_f_7__62_),
	.ck(clk),
	.d(n5338));
   ms00f80 proc_input_NIB_storage_data_f_reg_7__63_ (.o(proc_input_NIB_storage_data_f_7__63_),
	.ck(clk),
	.d(n5333));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__0_ (.o(proc_input_NIB_storage_data_f_6__0_),
	.ck(clk),
	.d(n5328));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__1_ (.o(proc_input_NIB_storage_data_f_6__1_),
	.ck(clk),
	.d(n5323));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__2_ (.o(proc_input_NIB_storage_data_f_6__2_),
	.ck(clk),
	.d(n5318));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__3_ (.o(proc_input_NIB_storage_data_f_6__3_),
	.ck(clk),
	.d(n5313));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__4_ (.o(proc_input_NIB_storage_data_f_6__4_),
	.ck(clk),
	.d(n5308));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__5_ (.o(proc_input_NIB_storage_data_f_6__5_),
	.ck(clk),
	.d(n5303));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__6_ (.o(proc_input_NIB_storage_data_f_6__6_),
	.ck(clk),
	.d(n5298));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__7_ (.o(proc_input_NIB_storage_data_f_6__7_),
	.ck(clk),
	.d(n5293));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__8_ (.o(proc_input_NIB_storage_data_f_6__8_),
	.ck(clk),
	.d(n5288));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__9_ (.o(proc_input_NIB_storage_data_f_6__9_),
	.ck(clk),
	.d(n5283));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__10_ (.o(proc_input_NIB_storage_data_f_6__10_),
	.ck(clk),
	.d(n5278));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__11_ (.o(proc_input_NIB_storage_data_f_6__11_),
	.ck(clk),
	.d(n5273));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__12_ (.o(proc_input_NIB_storage_data_f_6__12_),
	.ck(clk),
	.d(n5268));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__13_ (.o(proc_input_NIB_storage_data_f_6__13_),
	.ck(clk),
	.d(n5263));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__14_ (.o(proc_input_NIB_storage_data_f_6__14_),
	.ck(clk),
	.d(n5258));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__15_ (.o(proc_input_NIB_storage_data_f_6__15_),
	.ck(clk),
	.d(n5253));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__16_ (.o(proc_input_NIB_storage_data_f_6__16_),
	.ck(clk),
	.d(n5248));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__17_ (.o(proc_input_NIB_storage_data_f_6__17_),
	.ck(clk),
	.d(n5243));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__18_ (.o(proc_input_NIB_storage_data_f_6__18_),
	.ck(clk),
	.d(n5238));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__19_ (.o(proc_input_NIB_storage_data_f_6__19_),
	.ck(clk),
	.d(n5233));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__20_ (.o(proc_input_NIB_storage_data_f_6__20_),
	.ck(clk),
	.d(n5228));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__21_ (.o(proc_input_NIB_storage_data_f_6__21_),
	.ck(clk),
	.d(n5223));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__22_ (.o(proc_input_NIB_storage_data_f_6__22_),
	.ck(clk),
	.d(n5218));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__23_ (.o(proc_input_NIB_storage_data_f_6__23_),
	.ck(clk),
	.d(n5213));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__24_ (.o(proc_input_NIB_storage_data_f_6__24_),
	.ck(clk),
	.d(n5208));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__25_ (.o(proc_input_NIB_storage_data_f_6__25_),
	.ck(clk),
	.d(n5203));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__26_ (.o(proc_input_NIB_storage_data_f_6__26_),
	.ck(clk),
	.d(n5198));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__27_ (.o(proc_input_NIB_storage_data_f_6__27_),
	.ck(clk),
	.d(n5193));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__28_ (.o(proc_input_NIB_storage_data_f_6__28_),
	.ck(clk),
	.d(n5188));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__29_ (.o(proc_input_NIB_storage_data_f_6__29_),
	.ck(clk),
	.d(n5183));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__30_ (.o(proc_input_NIB_storage_data_f_6__30_),
	.ck(clk),
	.d(n5178));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__31_ (.o(proc_input_NIB_storage_data_f_6__31_),
	.ck(clk),
	.d(n5173));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__32_ (.o(proc_input_NIB_storage_data_f_6__32_),
	.ck(clk),
	.d(n5168));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__33_ (.o(proc_input_NIB_storage_data_f_6__33_),
	.ck(clk),
	.d(n5163));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__34_ (.o(proc_input_NIB_storage_data_f_6__34_),
	.ck(clk),
	.d(n5158));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__35_ (.o(proc_input_NIB_storage_data_f_6__35_),
	.ck(clk),
	.d(n5153));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__36_ (.o(proc_input_NIB_storage_data_f_6__36_),
	.ck(clk),
	.d(n5148));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__37_ (.o(proc_input_NIB_storage_data_f_6__37_),
	.ck(clk),
	.d(n5143));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__38_ (.o(proc_input_NIB_storage_data_f_6__38_),
	.ck(clk),
	.d(n5138));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__39_ (.o(proc_input_NIB_storage_data_f_6__39_),
	.ck(clk),
	.d(n5133));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__40_ (.o(proc_input_NIB_storage_data_f_6__40_),
	.ck(clk),
	.d(n5128));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__41_ (.o(proc_input_NIB_storage_data_f_6__41_),
	.ck(clk),
	.d(n5123));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__42_ (.o(proc_input_NIB_storage_data_f_6__42_),
	.ck(clk),
	.d(n5118));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__43_ (.o(proc_input_NIB_storage_data_f_6__43_),
	.ck(clk),
	.d(n5113));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__44_ (.o(proc_input_NIB_storage_data_f_6__44_),
	.ck(clk),
	.d(n5108));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__45_ (.o(proc_input_NIB_storage_data_f_6__45_),
	.ck(clk),
	.d(n5103));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__46_ (.o(proc_input_NIB_storage_data_f_6__46_),
	.ck(clk),
	.d(n5098));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__47_ (.o(proc_input_NIB_storage_data_f_6__47_),
	.ck(clk),
	.d(n5093));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__48_ (.o(proc_input_NIB_storage_data_f_6__48_),
	.ck(clk),
	.d(n5088));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__49_ (.o(proc_input_NIB_storage_data_f_6__49_),
	.ck(clk),
	.d(n5083));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__50_ (.o(proc_input_NIB_storage_data_f_6__50_),
	.ck(clk),
	.d(n5078));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__51_ (.o(proc_input_NIB_storage_data_f_6__51_),
	.ck(clk),
	.d(n5073));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__52_ (.o(proc_input_NIB_storage_data_f_6__52_),
	.ck(clk),
	.d(n5068));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__53_ (.o(proc_input_NIB_storage_data_f_6__53_),
	.ck(clk),
	.d(n5063));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__54_ (.o(proc_input_NIB_storage_data_f_6__54_),
	.ck(clk),
	.d(n5058));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__55_ (.o(proc_input_NIB_storage_data_f_6__55_),
	.ck(clk),
	.d(n5053));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__56_ (.o(proc_input_NIB_storage_data_f_6__56_),
	.ck(clk),
	.d(n5048));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__57_ (.o(proc_input_NIB_storage_data_f_6__57_),
	.ck(clk),
	.d(n5043));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__58_ (.o(proc_input_NIB_storage_data_f_6__58_),
	.ck(clk),
	.d(n5038));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__59_ (.o(proc_input_NIB_storage_data_f_6__59_),
	.ck(clk),
	.d(n5033));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__60_ (.o(proc_input_NIB_storage_data_f_6__60_),
	.ck(clk),
	.d(n5028));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__61_ (.o(proc_input_NIB_storage_data_f_6__61_),
	.ck(clk),
	.d(n5023));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__62_ (.o(proc_input_NIB_storage_data_f_6__62_),
	.ck(clk),
	.d(n5018));
   ms00f80 proc_input_NIB_storage_data_f_reg_6__63_ (.o(proc_input_NIB_storage_data_f_6__63_),
	.ck(clk),
	.d(n5013));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__0_ (.o(proc_input_NIB_storage_data_f_5__0_),
	.ck(clk),
	.d(n5008));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__1_ (.o(proc_input_NIB_storage_data_f_5__1_),
	.ck(clk),
	.d(n5003));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__2_ (.o(proc_input_NIB_storage_data_f_5__2_),
	.ck(clk),
	.d(n4998));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__3_ (.o(proc_input_NIB_storage_data_f_5__3_),
	.ck(clk),
	.d(n4993));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__4_ (.o(proc_input_NIB_storage_data_f_5__4_),
	.ck(clk),
	.d(n4988));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__5_ (.o(proc_input_NIB_storage_data_f_5__5_),
	.ck(clk),
	.d(n4983));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__6_ (.o(proc_input_NIB_storage_data_f_5__6_),
	.ck(clk),
	.d(n4978));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__7_ (.o(proc_input_NIB_storage_data_f_5__7_),
	.ck(clk),
	.d(n4973));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__8_ (.o(proc_input_NIB_storage_data_f_5__8_),
	.ck(clk),
	.d(n4968));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__9_ (.o(proc_input_NIB_storage_data_f_5__9_),
	.ck(clk),
	.d(n4963));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__10_ (.o(proc_input_NIB_storage_data_f_5__10_),
	.ck(clk),
	.d(n4958));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__11_ (.o(proc_input_NIB_storage_data_f_5__11_),
	.ck(clk),
	.d(n4953));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__12_ (.o(proc_input_NIB_storage_data_f_5__12_),
	.ck(clk),
	.d(n4948));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__13_ (.o(proc_input_NIB_storage_data_f_5__13_),
	.ck(clk),
	.d(n4943));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__14_ (.o(proc_input_NIB_storage_data_f_5__14_),
	.ck(clk),
	.d(n4938));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__15_ (.o(proc_input_NIB_storage_data_f_5__15_),
	.ck(clk),
	.d(n4933));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__16_ (.o(proc_input_NIB_storage_data_f_5__16_),
	.ck(clk),
	.d(n4928));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__17_ (.o(proc_input_NIB_storage_data_f_5__17_),
	.ck(clk),
	.d(n4923));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__18_ (.o(proc_input_NIB_storage_data_f_5__18_),
	.ck(clk),
	.d(n4918));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__19_ (.o(proc_input_NIB_storage_data_f_5__19_),
	.ck(clk),
	.d(n4913));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__20_ (.o(proc_input_NIB_storage_data_f_5__20_),
	.ck(clk),
	.d(n4908));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__21_ (.o(proc_input_NIB_storage_data_f_5__21_),
	.ck(clk),
	.d(n4903));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__22_ (.o(proc_input_NIB_storage_data_f_5__22_),
	.ck(clk),
	.d(n4898));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__23_ (.o(proc_input_NIB_storage_data_f_5__23_),
	.ck(clk),
	.d(n4893));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__24_ (.o(proc_input_NIB_storage_data_f_5__24_),
	.ck(clk),
	.d(n4888));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__25_ (.o(proc_input_NIB_storage_data_f_5__25_),
	.ck(clk),
	.d(n4883));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__26_ (.o(proc_input_NIB_storage_data_f_5__26_),
	.ck(clk),
	.d(n4878));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__27_ (.o(proc_input_NIB_storage_data_f_5__27_),
	.ck(clk),
	.d(n4873));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__28_ (.o(proc_input_NIB_storage_data_f_5__28_),
	.ck(clk),
	.d(n4868));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__29_ (.o(proc_input_NIB_storage_data_f_5__29_),
	.ck(clk),
	.d(n4863));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__30_ (.o(proc_input_NIB_storage_data_f_5__30_),
	.ck(clk),
	.d(n4858));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__31_ (.o(proc_input_NIB_storage_data_f_5__31_),
	.ck(clk),
	.d(n4853));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__32_ (.o(proc_input_NIB_storage_data_f_5__32_),
	.ck(clk),
	.d(n4848));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__33_ (.o(proc_input_NIB_storage_data_f_5__33_),
	.ck(clk),
	.d(n4843));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__34_ (.o(proc_input_NIB_storage_data_f_5__34_),
	.ck(clk),
	.d(n4838));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__35_ (.o(proc_input_NIB_storage_data_f_5__35_),
	.ck(clk),
	.d(n4833));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__36_ (.o(proc_input_NIB_storage_data_f_5__36_),
	.ck(clk),
	.d(n4828));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__37_ (.o(proc_input_NIB_storage_data_f_5__37_),
	.ck(clk),
	.d(n4823));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__38_ (.o(proc_input_NIB_storage_data_f_5__38_),
	.ck(clk),
	.d(n4818));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__39_ (.o(proc_input_NIB_storage_data_f_5__39_),
	.ck(clk),
	.d(n4813));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__40_ (.o(proc_input_NIB_storage_data_f_5__40_),
	.ck(clk),
	.d(n4808));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__41_ (.o(proc_input_NIB_storage_data_f_5__41_),
	.ck(clk),
	.d(n4803));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__42_ (.o(proc_input_NIB_storage_data_f_5__42_),
	.ck(clk),
	.d(n4798));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__43_ (.o(proc_input_NIB_storage_data_f_5__43_),
	.ck(clk),
	.d(n4793));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__44_ (.o(proc_input_NIB_storage_data_f_5__44_),
	.ck(clk),
	.d(n4788));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__45_ (.o(proc_input_NIB_storage_data_f_5__45_),
	.ck(clk),
	.d(n4783));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__46_ (.o(proc_input_NIB_storage_data_f_5__46_),
	.ck(clk),
	.d(n4778));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__47_ (.o(proc_input_NIB_storage_data_f_5__47_),
	.ck(clk),
	.d(n4773));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__48_ (.o(proc_input_NIB_storage_data_f_5__48_),
	.ck(clk),
	.d(n4768));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__49_ (.o(proc_input_NIB_storage_data_f_5__49_),
	.ck(clk),
	.d(n4763));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__50_ (.o(proc_input_NIB_storage_data_f_5__50_),
	.ck(clk),
	.d(n4758));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__51_ (.o(proc_input_NIB_storage_data_f_5__51_),
	.ck(clk),
	.d(n4753));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__52_ (.o(proc_input_NIB_storage_data_f_5__52_),
	.ck(clk),
	.d(n4748));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__53_ (.o(proc_input_NIB_storage_data_f_5__53_),
	.ck(clk),
	.d(n4743));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__54_ (.o(proc_input_NIB_storage_data_f_5__54_),
	.ck(clk),
	.d(n4738));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__55_ (.o(proc_input_NIB_storage_data_f_5__55_),
	.ck(clk),
	.d(n4733));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__56_ (.o(proc_input_NIB_storage_data_f_5__56_),
	.ck(clk),
	.d(n4728));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__57_ (.o(proc_input_NIB_storage_data_f_5__57_),
	.ck(clk),
	.d(n4723));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__58_ (.o(proc_input_NIB_storage_data_f_5__58_),
	.ck(clk),
	.d(n4718));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__59_ (.o(proc_input_NIB_storage_data_f_5__59_),
	.ck(clk),
	.d(n4713));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__60_ (.o(proc_input_NIB_storage_data_f_5__60_),
	.ck(clk),
	.d(n4708));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__61_ (.o(proc_input_NIB_storage_data_f_5__61_),
	.ck(clk),
	.d(n4703));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__62_ (.o(proc_input_NIB_storage_data_f_5__62_),
	.ck(clk),
	.d(n4698));
   ms00f80 proc_input_NIB_storage_data_f_reg_5__63_ (.o(proc_input_NIB_storage_data_f_5__63_),
	.ck(clk),
	.d(n4693));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__0_ (.o(proc_input_NIB_storage_data_f_4__0_),
	.ck(clk),
	.d(n4688));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__1_ (.o(proc_input_NIB_storage_data_f_4__1_),
	.ck(clk),
	.d(n4683));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__2_ (.o(proc_input_NIB_storage_data_f_4__2_),
	.ck(clk),
	.d(n4678));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__3_ (.o(proc_input_NIB_storage_data_f_4__3_),
	.ck(clk),
	.d(n4673));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__4_ (.o(proc_input_NIB_storage_data_f_4__4_),
	.ck(clk),
	.d(n4668));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__5_ (.o(proc_input_NIB_storage_data_f_4__5_),
	.ck(clk),
	.d(n4663));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__6_ (.o(proc_input_NIB_storage_data_f_4__6_),
	.ck(clk),
	.d(n4658));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__7_ (.o(proc_input_NIB_storage_data_f_4__7_),
	.ck(clk),
	.d(n4653));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__8_ (.o(proc_input_NIB_storage_data_f_4__8_),
	.ck(clk),
	.d(n4648));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__9_ (.o(proc_input_NIB_storage_data_f_4__9_),
	.ck(clk),
	.d(n4643));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__10_ (.o(proc_input_NIB_storage_data_f_4__10_),
	.ck(clk),
	.d(n4638));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__11_ (.o(proc_input_NIB_storage_data_f_4__11_),
	.ck(clk),
	.d(n4633));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__12_ (.o(proc_input_NIB_storage_data_f_4__12_),
	.ck(clk),
	.d(n4628));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__13_ (.o(proc_input_NIB_storage_data_f_4__13_),
	.ck(clk),
	.d(n4623));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__14_ (.o(proc_input_NIB_storage_data_f_4__14_),
	.ck(clk),
	.d(n4618));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__15_ (.o(proc_input_NIB_storage_data_f_4__15_),
	.ck(clk),
	.d(n4613));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__16_ (.o(proc_input_NIB_storage_data_f_4__16_),
	.ck(clk),
	.d(n4608));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__17_ (.o(proc_input_NIB_storage_data_f_4__17_),
	.ck(clk),
	.d(n4603));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__18_ (.o(proc_input_NIB_storage_data_f_4__18_),
	.ck(clk),
	.d(n4598));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__19_ (.o(proc_input_NIB_storage_data_f_4__19_),
	.ck(clk),
	.d(n4593));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__20_ (.o(proc_input_NIB_storage_data_f_4__20_),
	.ck(clk),
	.d(n4588));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__21_ (.o(proc_input_NIB_storage_data_f_4__21_),
	.ck(clk),
	.d(n4583));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__22_ (.o(proc_input_NIB_storage_data_f_4__22_),
	.ck(clk),
	.d(n4578));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__23_ (.o(proc_input_NIB_storage_data_f_4__23_),
	.ck(clk),
	.d(n4573));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__24_ (.o(proc_input_NIB_storage_data_f_4__24_),
	.ck(clk),
	.d(n4568));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__25_ (.o(proc_input_NIB_storage_data_f_4__25_),
	.ck(clk),
	.d(n4563));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__26_ (.o(proc_input_NIB_storage_data_f_4__26_),
	.ck(clk),
	.d(n4558));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__27_ (.o(proc_input_NIB_storage_data_f_4__27_),
	.ck(clk),
	.d(n4553));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__28_ (.o(proc_input_NIB_storage_data_f_4__28_),
	.ck(clk),
	.d(n4548));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__29_ (.o(proc_input_NIB_storage_data_f_4__29_),
	.ck(clk),
	.d(n4543));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__30_ (.o(proc_input_NIB_storage_data_f_4__30_),
	.ck(clk),
	.d(n4538));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__31_ (.o(proc_input_NIB_storage_data_f_4__31_),
	.ck(clk),
	.d(n4533));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__32_ (.o(proc_input_NIB_storage_data_f_4__32_),
	.ck(clk),
	.d(n4528));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__33_ (.o(proc_input_NIB_storage_data_f_4__33_),
	.ck(clk),
	.d(n4523));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__34_ (.o(proc_input_NIB_storage_data_f_4__34_),
	.ck(clk),
	.d(n4518));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__35_ (.o(proc_input_NIB_storage_data_f_4__35_),
	.ck(clk),
	.d(n4513));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__36_ (.o(proc_input_NIB_storage_data_f_4__36_),
	.ck(clk),
	.d(n4508));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__37_ (.o(proc_input_NIB_storage_data_f_4__37_),
	.ck(clk),
	.d(n4503));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__38_ (.o(proc_input_NIB_storage_data_f_4__38_),
	.ck(clk),
	.d(n4498));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__39_ (.o(proc_input_NIB_storage_data_f_4__39_),
	.ck(clk),
	.d(n4493));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__40_ (.o(proc_input_NIB_storage_data_f_4__40_),
	.ck(clk),
	.d(n4488));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__41_ (.o(proc_input_NIB_storage_data_f_4__41_),
	.ck(clk),
	.d(n4483));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__42_ (.o(proc_input_NIB_storage_data_f_4__42_),
	.ck(clk),
	.d(n4478));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__43_ (.o(proc_input_NIB_storage_data_f_4__43_),
	.ck(clk),
	.d(n4473));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__44_ (.o(proc_input_NIB_storage_data_f_4__44_),
	.ck(clk),
	.d(n4468));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__45_ (.o(proc_input_NIB_storage_data_f_4__45_),
	.ck(clk),
	.d(n4463));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__46_ (.o(proc_input_NIB_storage_data_f_4__46_),
	.ck(clk),
	.d(n4458));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__47_ (.o(proc_input_NIB_storage_data_f_4__47_),
	.ck(clk),
	.d(n4453));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__48_ (.o(proc_input_NIB_storage_data_f_4__48_),
	.ck(clk),
	.d(n4448));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__49_ (.o(proc_input_NIB_storage_data_f_4__49_),
	.ck(clk),
	.d(n4443));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__50_ (.o(proc_input_NIB_storage_data_f_4__50_),
	.ck(clk),
	.d(n4438));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__51_ (.o(proc_input_NIB_storage_data_f_4__51_),
	.ck(clk),
	.d(n4433));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__52_ (.o(proc_input_NIB_storage_data_f_4__52_),
	.ck(clk),
	.d(n4428));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__53_ (.o(proc_input_NIB_storage_data_f_4__53_),
	.ck(clk),
	.d(n4423));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__54_ (.o(proc_input_NIB_storage_data_f_4__54_),
	.ck(clk),
	.d(n4418));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__55_ (.o(proc_input_NIB_storage_data_f_4__55_),
	.ck(clk),
	.d(n4413));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__56_ (.o(proc_input_NIB_storage_data_f_4__56_),
	.ck(clk),
	.d(n4408));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__57_ (.o(proc_input_NIB_storage_data_f_4__57_),
	.ck(clk),
	.d(n4403));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__58_ (.o(proc_input_NIB_storage_data_f_4__58_),
	.ck(clk),
	.d(n4398));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__59_ (.o(proc_input_NIB_storage_data_f_4__59_),
	.ck(clk),
	.d(n4393));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__60_ (.o(proc_input_NIB_storage_data_f_4__60_),
	.ck(clk),
	.d(n4388));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__61_ (.o(proc_input_NIB_storage_data_f_4__61_),
	.ck(clk),
	.d(n4383));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__62_ (.o(proc_input_NIB_storage_data_f_4__62_),
	.ck(clk),
	.d(n4378));
   ms00f80 proc_input_NIB_storage_data_f_reg_4__63_ (.o(proc_input_NIB_storage_data_f_4__63_),
	.ck(clk),
	.d(n4373));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__0_ (.o(proc_input_NIB_storage_data_f_3__0_),
	.ck(clk),
	.d(n4368));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__1_ (.o(proc_input_NIB_storage_data_f_3__1_),
	.ck(clk),
	.d(n4363));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__2_ (.o(proc_input_NIB_storage_data_f_3__2_),
	.ck(clk),
	.d(n4358));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__3_ (.o(proc_input_NIB_storage_data_f_3__3_),
	.ck(clk),
	.d(n4353));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__4_ (.o(proc_input_NIB_storage_data_f_3__4_),
	.ck(clk),
	.d(n4348));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__5_ (.o(proc_input_NIB_storage_data_f_3__5_),
	.ck(clk),
	.d(n4343));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__6_ (.o(proc_input_NIB_storage_data_f_3__6_),
	.ck(clk),
	.d(n4338));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__7_ (.o(proc_input_NIB_storage_data_f_3__7_),
	.ck(clk),
	.d(n4333));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__8_ (.o(proc_input_NIB_storage_data_f_3__8_),
	.ck(clk),
	.d(n4328));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__9_ (.o(proc_input_NIB_storage_data_f_3__9_),
	.ck(clk),
	.d(n4323));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__10_ (.o(proc_input_NIB_storage_data_f_3__10_),
	.ck(clk),
	.d(n4318));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__11_ (.o(proc_input_NIB_storage_data_f_3__11_),
	.ck(clk),
	.d(n4313));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__12_ (.o(proc_input_NIB_storage_data_f_3__12_),
	.ck(clk),
	.d(n4308));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__13_ (.o(proc_input_NIB_storage_data_f_3__13_),
	.ck(clk),
	.d(n4303));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__14_ (.o(proc_input_NIB_storage_data_f_3__14_),
	.ck(clk),
	.d(n4298));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__15_ (.o(proc_input_NIB_storage_data_f_3__15_),
	.ck(clk),
	.d(n4293));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__16_ (.o(proc_input_NIB_storage_data_f_3__16_),
	.ck(clk),
	.d(n4288));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__17_ (.o(proc_input_NIB_storage_data_f_3__17_),
	.ck(clk),
	.d(n4283));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__18_ (.o(proc_input_NIB_storage_data_f_3__18_),
	.ck(clk),
	.d(n4278));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__19_ (.o(proc_input_NIB_storage_data_f_3__19_),
	.ck(clk),
	.d(n4273));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__20_ (.o(proc_input_NIB_storage_data_f_3__20_),
	.ck(clk),
	.d(n4268));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__21_ (.o(proc_input_NIB_storage_data_f_3__21_),
	.ck(clk),
	.d(n4263));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__22_ (.o(proc_input_NIB_storage_data_f_3__22_),
	.ck(clk),
	.d(n4258));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__23_ (.o(proc_input_NIB_storage_data_f_3__23_),
	.ck(clk),
	.d(n4253));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__24_ (.o(proc_input_NIB_storage_data_f_3__24_),
	.ck(clk),
	.d(n4248));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__25_ (.o(proc_input_NIB_storage_data_f_3__25_),
	.ck(clk),
	.d(n4243));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__26_ (.o(proc_input_NIB_storage_data_f_3__26_),
	.ck(clk),
	.d(n4238));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__27_ (.o(proc_input_NIB_storage_data_f_3__27_),
	.ck(clk),
	.d(n4233));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__28_ (.o(proc_input_NIB_storage_data_f_3__28_),
	.ck(clk),
	.d(n4228));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__29_ (.o(proc_input_NIB_storage_data_f_3__29_),
	.ck(clk),
	.d(n4223));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__30_ (.o(proc_input_NIB_storage_data_f_3__30_),
	.ck(clk),
	.d(n4218));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__31_ (.o(proc_input_NIB_storage_data_f_3__31_),
	.ck(clk),
	.d(n4213));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__32_ (.o(proc_input_NIB_storage_data_f_3__32_),
	.ck(clk),
	.d(n4208));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__33_ (.o(proc_input_NIB_storage_data_f_3__33_),
	.ck(clk),
	.d(n4203));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__34_ (.o(proc_input_NIB_storage_data_f_3__34_),
	.ck(clk),
	.d(n4198));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__35_ (.o(proc_input_NIB_storage_data_f_3__35_),
	.ck(clk),
	.d(n4193));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__36_ (.o(proc_input_NIB_storage_data_f_3__36_),
	.ck(clk),
	.d(n4188));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__37_ (.o(proc_input_NIB_storage_data_f_3__37_),
	.ck(clk),
	.d(n4183));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__38_ (.o(proc_input_NIB_storage_data_f_3__38_),
	.ck(clk),
	.d(n4178));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__39_ (.o(proc_input_NIB_storage_data_f_3__39_),
	.ck(clk),
	.d(n4173));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__40_ (.o(proc_input_NIB_storage_data_f_3__40_),
	.ck(clk),
	.d(n4168));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__41_ (.o(proc_input_NIB_storage_data_f_3__41_),
	.ck(clk),
	.d(n4163));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__42_ (.o(proc_input_NIB_storage_data_f_3__42_),
	.ck(clk),
	.d(n4158));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__43_ (.o(proc_input_NIB_storage_data_f_3__43_),
	.ck(clk),
	.d(n4153));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__44_ (.o(proc_input_NIB_storage_data_f_3__44_),
	.ck(clk),
	.d(n4148));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__45_ (.o(proc_input_NIB_storage_data_f_3__45_),
	.ck(clk),
	.d(n4143));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__46_ (.o(proc_input_NIB_storage_data_f_3__46_),
	.ck(clk),
	.d(n4138));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__47_ (.o(proc_input_NIB_storage_data_f_3__47_),
	.ck(clk),
	.d(n4133));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__48_ (.o(proc_input_NIB_storage_data_f_3__48_),
	.ck(clk),
	.d(n4128));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__49_ (.o(proc_input_NIB_storage_data_f_3__49_),
	.ck(clk),
	.d(n4123));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__50_ (.o(proc_input_NIB_storage_data_f_3__50_),
	.ck(clk),
	.d(n4118));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__51_ (.o(proc_input_NIB_storage_data_f_3__51_),
	.ck(clk),
	.d(n4113));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__52_ (.o(proc_input_NIB_storage_data_f_3__52_),
	.ck(clk),
	.d(n4108));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__53_ (.o(proc_input_NIB_storage_data_f_3__53_),
	.ck(clk),
	.d(n4103));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__54_ (.o(proc_input_NIB_storage_data_f_3__54_),
	.ck(clk),
	.d(n4098));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__55_ (.o(proc_input_NIB_storage_data_f_3__55_),
	.ck(clk),
	.d(n4093));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__56_ (.o(proc_input_NIB_storage_data_f_3__56_),
	.ck(clk),
	.d(n4088));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__57_ (.o(proc_input_NIB_storage_data_f_3__57_),
	.ck(clk),
	.d(n4083));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__58_ (.o(proc_input_NIB_storage_data_f_3__58_),
	.ck(clk),
	.d(n4078));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__59_ (.o(proc_input_NIB_storage_data_f_3__59_),
	.ck(clk),
	.d(n4073));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__60_ (.o(proc_input_NIB_storage_data_f_3__60_),
	.ck(clk),
	.d(n4068));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__61_ (.o(proc_input_NIB_storage_data_f_3__61_),
	.ck(clk),
	.d(n4063));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__62_ (.o(proc_input_NIB_storage_data_f_3__62_),
	.ck(clk),
	.d(n4058));
   ms00f80 proc_input_NIB_storage_data_f_reg_3__63_ (.o(proc_input_NIB_storage_data_f_3__63_),
	.ck(clk),
	.d(n4053));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__0_ (.o(proc_input_NIB_storage_data_f_2__0_),
	.ck(clk),
	.d(n4048));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__1_ (.o(proc_input_NIB_storage_data_f_2__1_),
	.ck(clk),
	.d(n4043));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__2_ (.o(proc_input_NIB_storage_data_f_2__2_),
	.ck(clk),
	.d(n4038));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__3_ (.o(proc_input_NIB_storage_data_f_2__3_),
	.ck(clk),
	.d(n4033));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__4_ (.o(proc_input_NIB_storage_data_f_2__4_),
	.ck(clk),
	.d(n4028));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__5_ (.o(proc_input_NIB_storage_data_f_2__5_),
	.ck(clk),
	.d(n4023));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__6_ (.o(proc_input_NIB_storage_data_f_2__6_),
	.ck(clk),
	.d(n4018));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__7_ (.o(proc_input_NIB_storage_data_f_2__7_),
	.ck(clk),
	.d(n4013));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__8_ (.o(proc_input_NIB_storage_data_f_2__8_),
	.ck(clk),
	.d(n4008));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__9_ (.o(proc_input_NIB_storage_data_f_2__9_),
	.ck(clk),
	.d(n4003));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__10_ (.o(proc_input_NIB_storage_data_f_2__10_),
	.ck(clk),
	.d(n3998));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__11_ (.o(proc_input_NIB_storage_data_f_2__11_),
	.ck(clk),
	.d(n3993));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__12_ (.o(proc_input_NIB_storage_data_f_2__12_),
	.ck(clk),
	.d(n3988));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__13_ (.o(proc_input_NIB_storage_data_f_2__13_),
	.ck(clk),
	.d(n3983));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__14_ (.o(proc_input_NIB_storage_data_f_2__14_),
	.ck(clk),
	.d(n3978));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__15_ (.o(proc_input_NIB_storage_data_f_2__15_),
	.ck(clk),
	.d(n3973));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__16_ (.o(proc_input_NIB_storage_data_f_2__16_),
	.ck(clk),
	.d(n3968));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__17_ (.o(proc_input_NIB_storage_data_f_2__17_),
	.ck(clk),
	.d(n3963));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__18_ (.o(proc_input_NIB_storage_data_f_2__18_),
	.ck(clk),
	.d(n3958));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__19_ (.o(proc_input_NIB_storage_data_f_2__19_),
	.ck(clk),
	.d(n3953));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__20_ (.o(proc_input_NIB_storage_data_f_2__20_),
	.ck(clk),
	.d(n3948));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__21_ (.o(proc_input_NIB_storage_data_f_2__21_),
	.ck(clk),
	.d(n3943));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__22_ (.o(proc_input_NIB_storage_data_f_2__22_),
	.ck(clk),
	.d(n3938));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__23_ (.o(proc_input_NIB_storage_data_f_2__23_),
	.ck(clk),
	.d(n3933));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__24_ (.o(proc_input_NIB_storage_data_f_2__24_),
	.ck(clk),
	.d(n3928));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__25_ (.o(proc_input_NIB_storage_data_f_2__25_),
	.ck(clk),
	.d(n3923));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__26_ (.o(proc_input_NIB_storage_data_f_2__26_),
	.ck(clk),
	.d(n3918));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__27_ (.o(proc_input_NIB_storage_data_f_2__27_),
	.ck(clk),
	.d(n3913));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__28_ (.o(proc_input_NIB_storage_data_f_2__28_),
	.ck(clk),
	.d(n3908));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__29_ (.o(proc_input_NIB_storage_data_f_2__29_),
	.ck(clk),
	.d(n3903));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__30_ (.o(proc_input_NIB_storage_data_f_2__30_),
	.ck(clk),
	.d(n3898));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__31_ (.o(proc_input_NIB_storage_data_f_2__31_),
	.ck(clk),
	.d(n3893));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__32_ (.o(proc_input_NIB_storage_data_f_2__32_),
	.ck(clk),
	.d(n3888));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__33_ (.o(proc_input_NIB_storage_data_f_2__33_),
	.ck(clk),
	.d(n3883));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__34_ (.o(proc_input_NIB_storage_data_f_2__34_),
	.ck(clk),
	.d(n3878));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__35_ (.o(proc_input_NIB_storage_data_f_2__35_),
	.ck(clk),
	.d(n3873));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__36_ (.o(proc_input_NIB_storage_data_f_2__36_),
	.ck(clk),
	.d(n3868));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__37_ (.o(proc_input_NIB_storage_data_f_2__37_),
	.ck(clk),
	.d(n3863));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__38_ (.o(proc_input_NIB_storage_data_f_2__38_),
	.ck(clk),
	.d(n3858));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__39_ (.o(proc_input_NIB_storage_data_f_2__39_),
	.ck(clk),
	.d(n3853));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__40_ (.o(proc_input_NIB_storage_data_f_2__40_),
	.ck(clk),
	.d(n3848));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__41_ (.o(proc_input_NIB_storage_data_f_2__41_),
	.ck(clk),
	.d(n3843));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__42_ (.o(proc_input_NIB_storage_data_f_2__42_),
	.ck(clk),
	.d(n3838));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__43_ (.o(proc_input_NIB_storage_data_f_2__43_),
	.ck(clk),
	.d(n3833));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__44_ (.o(proc_input_NIB_storage_data_f_2__44_),
	.ck(clk),
	.d(n3828));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__45_ (.o(proc_input_NIB_storage_data_f_2__45_),
	.ck(clk),
	.d(n3823));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__46_ (.o(proc_input_NIB_storage_data_f_2__46_),
	.ck(clk),
	.d(n3818));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__47_ (.o(proc_input_NIB_storage_data_f_2__47_),
	.ck(clk),
	.d(n3813));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__48_ (.o(proc_input_NIB_storage_data_f_2__48_),
	.ck(clk),
	.d(n3808));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__49_ (.o(proc_input_NIB_storage_data_f_2__49_),
	.ck(clk),
	.d(n3803));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__50_ (.o(proc_input_NIB_storage_data_f_2__50_),
	.ck(clk),
	.d(n3798));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__51_ (.o(proc_input_NIB_storage_data_f_2__51_),
	.ck(clk),
	.d(n3793));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__52_ (.o(proc_input_NIB_storage_data_f_2__52_),
	.ck(clk),
	.d(n3788));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__53_ (.o(proc_input_NIB_storage_data_f_2__53_),
	.ck(clk),
	.d(n3783));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__54_ (.o(proc_input_NIB_storage_data_f_2__54_),
	.ck(clk),
	.d(n3778));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__55_ (.o(proc_input_NIB_storage_data_f_2__55_),
	.ck(clk),
	.d(n3773));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__56_ (.o(proc_input_NIB_storage_data_f_2__56_),
	.ck(clk),
	.d(n3768));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__57_ (.o(proc_input_NIB_storage_data_f_2__57_),
	.ck(clk),
	.d(n3763));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__58_ (.o(proc_input_NIB_storage_data_f_2__58_),
	.ck(clk),
	.d(n3758));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__59_ (.o(proc_input_NIB_storage_data_f_2__59_),
	.ck(clk),
	.d(n3753));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__60_ (.o(proc_input_NIB_storage_data_f_2__60_),
	.ck(clk),
	.d(n3748));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__61_ (.o(proc_input_NIB_storage_data_f_2__61_),
	.ck(clk),
	.d(n3743));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__62_ (.o(proc_input_NIB_storage_data_f_2__62_),
	.ck(clk),
	.d(n3738));
   ms00f80 proc_input_NIB_storage_data_f_reg_2__63_ (.o(proc_input_NIB_storage_data_f_2__63_),
	.ck(clk),
	.d(n3733));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__0_ (.o(proc_input_NIB_storage_data_f_1__0_),
	.ck(clk),
	.d(n3728));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__1_ (.o(proc_input_NIB_storage_data_f_1__1_),
	.ck(clk),
	.d(n3723));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__2_ (.o(proc_input_NIB_storage_data_f_1__2_),
	.ck(clk),
	.d(n3718));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__3_ (.o(proc_input_NIB_storage_data_f_1__3_),
	.ck(clk),
	.d(n3713));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__4_ (.o(proc_input_NIB_storage_data_f_1__4_),
	.ck(clk),
	.d(n3708));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__5_ (.o(proc_input_NIB_storage_data_f_1__5_),
	.ck(clk),
	.d(n3703));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__6_ (.o(proc_input_NIB_storage_data_f_1__6_),
	.ck(clk),
	.d(n3698));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__7_ (.o(proc_input_NIB_storage_data_f_1__7_),
	.ck(clk),
	.d(n3693));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__8_ (.o(proc_input_NIB_storage_data_f_1__8_),
	.ck(clk),
	.d(n3688));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__9_ (.o(proc_input_NIB_storage_data_f_1__9_),
	.ck(clk),
	.d(n3683));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__10_ (.o(proc_input_NIB_storage_data_f_1__10_),
	.ck(clk),
	.d(n3678));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__11_ (.o(proc_input_NIB_storage_data_f_1__11_),
	.ck(clk),
	.d(n3673));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__12_ (.o(proc_input_NIB_storage_data_f_1__12_),
	.ck(clk),
	.d(n3668));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__13_ (.o(proc_input_NIB_storage_data_f_1__13_),
	.ck(clk),
	.d(n3663));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__14_ (.o(proc_input_NIB_storage_data_f_1__14_),
	.ck(clk),
	.d(n3658));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__15_ (.o(proc_input_NIB_storage_data_f_1__15_),
	.ck(clk),
	.d(n3653));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__16_ (.o(proc_input_NIB_storage_data_f_1__16_),
	.ck(clk),
	.d(n3648));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__17_ (.o(proc_input_NIB_storage_data_f_1__17_),
	.ck(clk),
	.d(n3643));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__18_ (.o(proc_input_NIB_storage_data_f_1__18_),
	.ck(clk),
	.d(n3638));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__19_ (.o(proc_input_NIB_storage_data_f_1__19_),
	.ck(clk),
	.d(n3633));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__20_ (.o(proc_input_NIB_storage_data_f_1__20_),
	.ck(clk),
	.d(n3628));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__21_ (.o(proc_input_NIB_storage_data_f_1__21_),
	.ck(clk),
	.d(n3623));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__22_ (.o(proc_input_NIB_storage_data_f_1__22_),
	.ck(clk),
	.d(n3618));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__23_ (.o(proc_input_NIB_storage_data_f_1__23_),
	.ck(clk),
	.d(n3613));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__24_ (.o(proc_input_NIB_storage_data_f_1__24_),
	.ck(clk),
	.d(n3608));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__25_ (.o(proc_input_NIB_storage_data_f_1__25_),
	.ck(clk),
	.d(n3603));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__26_ (.o(proc_input_NIB_storage_data_f_1__26_),
	.ck(clk),
	.d(n3598));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__27_ (.o(proc_input_NIB_storage_data_f_1__27_),
	.ck(clk),
	.d(n3593));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__28_ (.o(proc_input_NIB_storage_data_f_1__28_),
	.ck(clk),
	.d(n3588));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__29_ (.o(proc_input_NIB_storage_data_f_1__29_),
	.ck(clk),
	.d(n3583));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__30_ (.o(proc_input_NIB_storage_data_f_1__30_),
	.ck(clk),
	.d(n3578));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__31_ (.o(proc_input_NIB_storage_data_f_1__31_),
	.ck(clk),
	.d(n3573));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__32_ (.o(proc_input_NIB_storage_data_f_1__32_),
	.ck(clk),
	.d(n3568));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__33_ (.o(proc_input_NIB_storage_data_f_1__33_),
	.ck(clk),
	.d(n3563));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__34_ (.o(proc_input_NIB_storage_data_f_1__34_),
	.ck(clk),
	.d(n3558));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__35_ (.o(proc_input_NIB_storage_data_f_1__35_),
	.ck(clk),
	.d(n3553));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__36_ (.o(proc_input_NIB_storage_data_f_1__36_),
	.ck(clk),
	.d(n3548));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__37_ (.o(proc_input_NIB_storage_data_f_1__37_),
	.ck(clk),
	.d(n3543));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__38_ (.o(proc_input_NIB_storage_data_f_1__38_),
	.ck(clk),
	.d(n3538));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__39_ (.o(proc_input_NIB_storage_data_f_1__39_),
	.ck(clk),
	.d(n3533));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__40_ (.o(proc_input_NIB_storage_data_f_1__40_),
	.ck(clk),
	.d(n3528));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__41_ (.o(proc_input_NIB_storage_data_f_1__41_),
	.ck(clk),
	.d(n3523));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__42_ (.o(proc_input_NIB_storage_data_f_1__42_),
	.ck(clk),
	.d(n3518));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__43_ (.o(proc_input_NIB_storage_data_f_1__43_),
	.ck(clk),
	.d(n3513));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__44_ (.o(proc_input_NIB_storage_data_f_1__44_),
	.ck(clk),
	.d(n3508));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__45_ (.o(proc_input_NIB_storage_data_f_1__45_),
	.ck(clk),
	.d(n3503));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__46_ (.o(proc_input_NIB_storage_data_f_1__46_),
	.ck(clk),
	.d(n3498));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__47_ (.o(proc_input_NIB_storage_data_f_1__47_),
	.ck(clk),
	.d(n3493));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__48_ (.o(proc_input_NIB_storage_data_f_1__48_),
	.ck(clk),
	.d(n3488));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__49_ (.o(proc_input_NIB_storage_data_f_1__49_),
	.ck(clk),
	.d(n3483));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__50_ (.o(proc_input_NIB_storage_data_f_1__50_),
	.ck(clk),
	.d(n3478));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__51_ (.o(proc_input_NIB_storage_data_f_1__51_),
	.ck(clk),
	.d(n3473));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__52_ (.o(proc_input_NIB_storage_data_f_1__52_),
	.ck(clk),
	.d(n3468));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__53_ (.o(proc_input_NIB_storage_data_f_1__53_),
	.ck(clk),
	.d(n3463));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__54_ (.o(proc_input_NIB_storage_data_f_1__54_),
	.ck(clk),
	.d(n3458));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__55_ (.o(proc_input_NIB_storage_data_f_1__55_),
	.ck(clk),
	.d(n3453));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__56_ (.o(proc_input_NIB_storage_data_f_1__56_),
	.ck(clk),
	.d(n3448));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__57_ (.o(proc_input_NIB_storage_data_f_1__57_),
	.ck(clk),
	.d(n3443));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__58_ (.o(proc_input_NIB_storage_data_f_1__58_),
	.ck(clk),
	.d(n3438));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__59_ (.o(proc_input_NIB_storage_data_f_1__59_),
	.ck(clk),
	.d(n3433));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__60_ (.o(proc_input_NIB_storage_data_f_1__60_),
	.ck(clk),
	.d(n3428));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__61_ (.o(proc_input_NIB_storage_data_f_1__61_),
	.ck(clk),
	.d(n3423));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__62_ (.o(proc_input_NIB_storage_data_f_1__62_),
	.ck(clk),
	.d(n3418));
   ms00f80 proc_input_NIB_storage_data_f_reg_1__63_ (.o(proc_input_NIB_storage_data_f_1__63_),
	.ck(clk),
	.d(n3413));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__0_ (.o(proc_input_NIB_storage_data_f_0__0_),
	.ck(clk),
	.d(n3408));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__1_ (.o(proc_input_NIB_storage_data_f_0__1_),
	.ck(clk),
	.d(n3403));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__2_ (.o(proc_input_NIB_storage_data_f_0__2_),
	.ck(clk),
	.d(n3398));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__3_ (.o(proc_input_NIB_storage_data_f_0__3_),
	.ck(clk),
	.d(n3393));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__4_ (.o(proc_input_NIB_storage_data_f_0__4_),
	.ck(clk),
	.d(n3388));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__5_ (.o(proc_input_NIB_storage_data_f_0__5_),
	.ck(clk),
	.d(n3383));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__6_ (.o(proc_input_NIB_storage_data_f_0__6_),
	.ck(clk),
	.d(n3378));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__7_ (.o(proc_input_NIB_storage_data_f_0__7_),
	.ck(clk),
	.d(n3373));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__8_ (.o(proc_input_NIB_storage_data_f_0__8_),
	.ck(clk),
	.d(n3368));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__9_ (.o(proc_input_NIB_storage_data_f_0__9_),
	.ck(clk),
	.d(n3363));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__10_ (.o(proc_input_NIB_storage_data_f_0__10_),
	.ck(clk),
	.d(n3358));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__11_ (.o(proc_input_NIB_storage_data_f_0__11_),
	.ck(clk),
	.d(n3353));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__12_ (.o(proc_input_NIB_storage_data_f_0__12_),
	.ck(clk),
	.d(n3348));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__13_ (.o(proc_input_NIB_storage_data_f_0__13_),
	.ck(clk),
	.d(n3343));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__14_ (.o(proc_input_NIB_storage_data_f_0__14_),
	.ck(clk),
	.d(n3338));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__15_ (.o(proc_input_NIB_storage_data_f_0__15_),
	.ck(clk),
	.d(n3333));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__16_ (.o(proc_input_NIB_storage_data_f_0__16_),
	.ck(clk),
	.d(n3328));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__17_ (.o(proc_input_NIB_storage_data_f_0__17_),
	.ck(clk),
	.d(n3323));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__18_ (.o(proc_input_NIB_storage_data_f_0__18_),
	.ck(clk),
	.d(n3318));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__19_ (.o(proc_input_NIB_storage_data_f_0__19_),
	.ck(clk),
	.d(n3313));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__20_ (.o(proc_input_NIB_storage_data_f_0__20_),
	.ck(clk),
	.d(n3308));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__21_ (.o(proc_input_NIB_storage_data_f_0__21_),
	.ck(clk),
	.d(n3303));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__22_ (.o(proc_input_NIB_storage_data_f_0__22_),
	.ck(clk),
	.d(n3298));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__23_ (.o(proc_input_NIB_storage_data_f_0__23_),
	.ck(clk),
	.d(n3293));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__24_ (.o(proc_input_NIB_storage_data_f_0__24_),
	.ck(clk),
	.d(n3288));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__25_ (.o(proc_input_NIB_storage_data_f_0__25_),
	.ck(clk),
	.d(n3283));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__26_ (.o(proc_input_NIB_storage_data_f_0__26_),
	.ck(clk),
	.d(n3278));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__27_ (.o(proc_input_NIB_storage_data_f_0__27_),
	.ck(clk),
	.d(n3273));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__28_ (.o(proc_input_NIB_storage_data_f_0__28_),
	.ck(clk),
	.d(n3268));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__29_ (.o(proc_input_NIB_storage_data_f_0__29_),
	.ck(clk),
	.d(n3263));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__30_ (.o(proc_input_NIB_storage_data_f_0__30_),
	.ck(clk),
	.d(n3258));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__31_ (.o(proc_input_NIB_storage_data_f_0__31_),
	.ck(clk),
	.d(n3253));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__32_ (.o(proc_input_NIB_storage_data_f_0__32_),
	.ck(clk),
	.d(n3248));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__33_ (.o(proc_input_NIB_storage_data_f_0__33_),
	.ck(clk),
	.d(n3243));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__34_ (.o(proc_input_NIB_storage_data_f_0__34_),
	.ck(clk),
	.d(n3238));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__35_ (.o(proc_input_NIB_storage_data_f_0__35_),
	.ck(clk),
	.d(n3233));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__36_ (.o(proc_input_NIB_storage_data_f_0__36_),
	.ck(clk),
	.d(n3228));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__37_ (.o(proc_input_NIB_storage_data_f_0__37_),
	.ck(clk),
	.d(n3223));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__38_ (.o(proc_input_NIB_storage_data_f_0__38_),
	.ck(clk),
	.d(n3218));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__39_ (.o(proc_input_NIB_storage_data_f_0__39_),
	.ck(clk),
	.d(n3213));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__40_ (.o(proc_input_NIB_storage_data_f_0__40_),
	.ck(clk),
	.d(n3208));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__41_ (.o(proc_input_NIB_storage_data_f_0__41_),
	.ck(clk),
	.d(n3203));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__42_ (.o(proc_input_NIB_storage_data_f_0__42_),
	.ck(clk),
	.d(n3198));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__43_ (.o(proc_input_NIB_storage_data_f_0__43_),
	.ck(clk),
	.d(n3193));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__44_ (.o(proc_input_NIB_storage_data_f_0__44_),
	.ck(clk),
	.d(n3188));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__45_ (.o(proc_input_NIB_storage_data_f_0__45_),
	.ck(clk),
	.d(n3183));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__46_ (.o(proc_input_NIB_storage_data_f_0__46_),
	.ck(clk),
	.d(n3178));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__47_ (.o(proc_input_NIB_storage_data_f_0__47_),
	.ck(clk),
	.d(n3173));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__48_ (.o(proc_input_NIB_storage_data_f_0__48_),
	.ck(clk),
	.d(n3168));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__49_ (.o(proc_input_NIB_storage_data_f_0__49_),
	.ck(clk),
	.d(n3163));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__50_ (.o(proc_input_NIB_storage_data_f_0__50_),
	.ck(clk),
	.d(n3158));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__51_ (.o(proc_input_NIB_storage_data_f_0__51_),
	.ck(clk),
	.d(n3153));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__52_ (.o(proc_input_NIB_storage_data_f_0__52_),
	.ck(clk),
	.d(n3148));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__53_ (.o(proc_input_NIB_storage_data_f_0__53_),
	.ck(clk),
	.d(n3143));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__54_ (.o(proc_input_NIB_storage_data_f_0__54_),
	.ck(clk),
	.d(n3138));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__55_ (.o(proc_input_NIB_storage_data_f_0__55_),
	.ck(clk),
	.d(n3133));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__56_ (.o(proc_input_NIB_storage_data_f_0__56_),
	.ck(clk),
	.d(n3128));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__57_ (.o(proc_input_NIB_storage_data_f_0__57_),
	.ck(clk),
	.d(n3123));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__58_ (.o(proc_input_NIB_storage_data_f_0__58_),
	.ck(clk),
	.d(n3118));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__59_ (.o(proc_input_NIB_storage_data_f_0__59_),
	.ck(clk),
	.d(n3113));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__60_ (.o(proc_input_NIB_storage_data_f_0__60_),
	.ck(clk),
	.d(n3108));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__61_ (.o(proc_input_NIB_storage_data_f_0__61_),
	.ck(clk),
	.d(n3103));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__62_ (.o(proc_input_NIB_storage_data_f_0__62_),
	.ck(clk),
	.d(n3098));
   ms00f80 proc_input_NIB_storage_data_f_reg_0__63_ (.o(proc_input_NIB_storage_data_f_0__63_),
	.ck(clk),
	.d(n3093));
   ms00f80 north_output_space_yummy_f_reg (.o(north_output_space_yummy_f),
	.ck(clk),
	.d(north_output_space_N45));
   ms00f80 east_output_space_yummy_f_reg (.o(east_output_space_yummy_f),
	.ck(clk),
	.d(east_output_space_N45));
   ms00f80 south_output_space_yummy_f_reg (.o(south_output_space_yummy_f),
	.ck(clk),
	.d(south_output_space_N45));
   ms00f80 west_output_space_yummy_f_reg (.o(west_output_space_yummy_f),
	.ck(clk),
	.d(west_output_space_N45));
   ms00f80 proc_output_space_yummy_f_reg (.o(proc_output_space_yummy_f),
	.ck(clk),
	.d(proc_output_space_N45));
   ms00f80 proc_output_control_current_route_f_reg_2_ (.o(proc_output_current_route_connection_2_),
	.ck(clk),
	.d(proc_output_control_N469));
   ms00f80 proc_output_space_valid_f_reg (.o(proc_output_space_valid_f),
	.ck(clk),
	.d(proc_output_space_N46));
   ms00f80 proc_output_space_count_f_reg_2_ (.o(proc_output_space_count_f_2_),
	.ck(clk),
	.d(proc_output_space_N44));
   ms00f80 proc_output_space_is_two_or_more_f_reg (.o(proc_output_space_is_two_or_more_f),
	.ck(clk),
	.d(proc_output_space_N48));
   ms00f80 proc_output_space_count_f_reg_1_ (.o(proc_output_space_count_f_1_),
	.ck(clk),
	.d(proc_output_space_N43));
   ms00f80 proc_output_space_is_one_f_reg (.o(proc_output_space_is_one_f),
	.ck(clk),
	.d(proc_output_space_N47));
   ms00f80 proc_output_space_count_f_reg_0_ (.o(proc_output_space_count_f_0_),
	.ck(clk),
	.d(proc_output_space_N42));
   ms00f80 ec_thanks_p_to_p_reg_reg (.o(ec_thanks_p_to_p_reg),
	.ck(clk),
	.d(n26006));
   ms00f80 south_input_control_thanks_all_f_reg (.o(south_input_control_thanks_all_f),
	.ck(clk),
	.d(FE_RN_3));
   ms00f80 south_input_NIB_yummy_out_f_reg (.o(yummyOut_S),
	.ck(clk),
	.d(FE_RN_3));
   ms00f80 south_input_NIB_elements_in_array_f_reg_0_ (.o(south_input_NIB_elements_in_array_f_0_),
	.ck(clk),
	.d(n25991));
   ms00f80 south_input_NIB_elements_in_array_f_reg_1_ (.o(south_input_NIB_elements_in_array_f_1_),
	.ck(clk),
	.d(n25990));
   ms00f80 south_input_NIB_elements_in_array_f_reg_2_ (.o(south_input_NIB_elements_in_array_f_2_),
	.ck(clk),
	.d(n3003));
   ms00f80 ec_south_input_valid_reg_reg (.o(ec_south_input_valid_reg),
	.ck(clk),
	.d(south_input_valid));
   ms00f80 south_input_NIB_head_ptr_f_reg_0_ (.o(south_input_NIB_head_ptr_f_0_),
	.ck(clk),
	.d(n2993));
   ms00f80 south_input_NIB_head_ptr_f_reg_1_ (.o(south_input_NIB_head_ptr_f_1_),
	.ck(clk),
	.d(n2988));
   ms00f80 south_input_control_count_zero_f_reg (.o(south_input_control_count_zero_f),
	.ck(clk),
	.d(south_input_control_N51));
   ms00f80 south_input_control_header_last_f_reg (.o(south_input_control_header_last_f),
	.ck(clk),
	.d(south_input_control_N49));
   ms00f80 south_input_control_count_f_reg_0_ (.o(south_input_control_count_f_0_),
	.ck(clk),
	.d(n26026));
   ms00f80 south_input_control_count_f_reg_1_ (.o(south_input_control_count_f_1_),
	.ck(clk),
	.d(south_input_control_N42));
   ms00f80 south_input_control_count_f_reg_2_ (.o(south_input_control_count_f_2_),
	.ck(clk),
	.d(south_input_control_N43));
   ms00f80 south_input_control_count_f_reg_3_ (.o(south_input_control_count_f_3_),
	.ck(clk),
	.d(south_input_control_N44));
   ms00f80 south_input_control_count_f_reg_4_ (.o(south_input_control_count_f_4_),
	.ck(clk),
	.d(south_input_control_N45));
   ms00f80 south_input_control_count_f_reg_5_ (.o(south_input_control_count_f_5_),
	.ck(clk),
	.d(south_input_control_N46));
   ms00f80 south_input_control_count_f_reg_6_ (.o(south_input_control_count_f_6_),
	.ck(clk),
	.d(south_input_control_N47));
   ms00f80 south_input_control_count_f_reg_7_ (.o(south_input_control_count_f_7_),
	.ck(clk),
	.d(south_input_control_N48));
   ms00f80 south_input_control_count_one_f_reg (.o(south_input_control_count_one_f),
	.ck(clk),
	.d(south_input_control_N52));
   ms00f80 south_input_control_tail_last_f_reg (.o(south_input_control_tail_last_f),
	.ck(clk),
	.d(south_input_control_N53));
   ms00f80 north_output_space_valid_f_reg (.o(north_output_space_valid_f),
	.ck(clk),
	.d(north_output_space_N46));
   ms00f80 north_output_space_count_f_reg_2_ (.o(north_output_space_count_f_2_),
	.ck(clk),
	.d(north_output_space_N44));
   ms00f80 north_output_space_is_two_or_more_f_reg (.o(north_output_space_is_two_or_more_f),
	.ck(clk),
	.d(north_output_space_N48));
   ms00f80 north_output_space_count_f_reg_1_ (.o(north_output_space_count_f_1_),
	.ck(clk),
	.d(north_output_space_N43));
   ms00f80 north_output_space_is_one_f_reg (.o(north_output_space_is_one_f),
	.ck(clk),
	.d(north_output_space_N47));
   ms00f80 north_output_space_count_f_reg_0_ (.o(north_output_space_count_f_0_),
	.ck(clk),
	.d(north_output_space_N42));
   ms00f80 north_output_control_ec_wants_to_send_but_cannot_reg (.o(ec_wants_to_send_but_cannot_N),
	.ck(clk),
	.d(north_output_control_N72));
   ms00f80 ec_thanks_n_to_p_reg_reg (.o(ec_thanks_n_to_p_reg),
	.ck(clk),
	.d(n26023));
   ms00f80 proc_input_control_thanks_all_f_reg (.o(proc_input_control_thanks_all_f),
	.ck(clk),
	.d(n25995));
   ms00f80 proc_input_NIB_yummy_out_f_reg (.o(yummyOut_P),
	.ck(clk),
	.d(n25995));
   ms00f80 proc_input_NIB_head_ptr_f_reg_0_ (.o(proc_input_NIB_head_ptr_f_0_),
	.ck(clk),
	.d(n2873));
   ms00f80 proc_input_NIB_head_ptr_f_reg_1_ (.o(proc_input_NIB_head_ptr_f_1_),
	.ck(clk),
	.d(n2868));
   ms00f80 proc_input_NIB_head_ptr_f_reg_2_ (.o(proc_input_NIB_head_ptr_f_2_),
	.ck(clk),
	.d(n2863));
   ms00f80 proc_input_NIB_head_ptr_f_reg_3_ (.o(proc_input_NIB_head_ptr_f_3_),
	.ck(clk),
	.d(n2858));
   ms00f80 proc_input_NIB_elements_in_array_f_reg_0_ (.o(proc_input_NIB_elements_in_array_f_0_),
	.ck(clk),
	.d(n2853));
   ms00f80 proc_input_NIB_elements_in_array_f_reg_1_ (.o(proc_input_NIB_elements_in_array_f_1_),
	.ck(clk),
	.d(n2848));
   ms00f80 proc_input_NIB_elements_in_array_f_reg_2_ (.o(proc_input_NIB_elements_in_array_f_2_),
	.ck(clk),
	.d(n2843));
   ms00f80 proc_input_NIB_elements_in_array_f_reg_3_ (.o(proc_input_NIB_elements_in_array_f_3_),
	.ck(clk),
	.d(n2838));
   ms00f80 proc_input_NIB_elements_in_array_f_reg_4_ (.o(proc_input_NIB_elements_in_array_f_4_),
	.ck(clk),
	.d(n2833));
   ms00f80 ec_proc_input_valid_reg_reg (.o(ec_proc_input_valid_reg),
	.ck(clk),
	.d(proc_input_valid));
   ms00f80 proc_input_control_count_f_reg_0_ (.o(proc_input_control_count_f_0_),
	.ck(clk),
	.d(proc_input_control_N41));
   ms00f80 proc_input_control_count_f_reg_1_ (.o(proc_input_control_count_f_1_),
	.ck(clk),
	.d(proc_input_control_N42));
   ms00f80 proc_input_control_count_f_reg_2_ (.o(proc_input_control_count_f_2_),
	.ck(clk),
	.d(proc_input_control_N43));
   ms00f80 proc_input_control_count_f_reg_3_ (.o(proc_input_control_count_f_3_),
	.ck(clk),
	.d(proc_input_control_N44));
   ms00f80 proc_input_control_count_f_reg_4_ (.o(proc_input_control_count_f_4_),
	.ck(clk),
	.d(proc_input_control_N45));
   ms00f80 proc_input_control_count_f_reg_5_ (.o(proc_input_control_count_f_5_),
	.ck(clk),
	.d(proc_input_control_N46));
   ms00f80 proc_input_control_count_f_reg_6_ (.o(proc_input_control_count_f_6_),
	.ck(clk),
	.d(proc_input_control_N47));
   ms00f80 proc_input_control_count_f_reg_7_ (.o(proc_input_control_count_f_7_),
	.ck(clk),
	.d(proc_input_control_N48));
   ms00f80 proc_input_control_count_one_f_reg (.o(proc_input_control_count_one_f),
	.ck(clk),
	.d(proc_input_control_N52));
   ms00f80 proc_input_control_count_zero_f_reg (.o(proc_input_control_count_zero_f),
	.ck(clk),
	.d(proc_input_control_N51));
   ms00f80 proc_input_control_header_last_f_reg (.o(proc_input_control_header_last_f),
	.ck(clk),
	.d(proc_input_control_N49));
   ms00f80 proc_input_control_tail_last_f_reg (.o(proc_input_control_tail_last_f),
	.ck(clk),
	.d(proc_input_control_N53));
   ms00f80 east_output_space_valid_f_reg (.o(east_output_space_valid_f),
	.ck(clk),
	.d(east_output_space_N46));
   ms00f80 east_output_space_count_f_reg_2_ (.o(east_output_space_count_f_2_),
	.ck(clk),
	.d(east_output_space_N44));
   ms00f80 east_output_space_is_two_or_more_f_reg (.o(east_output_space_is_two_or_more_f),
	.ck(clk),
	.d(east_output_space_N48));
   ms00f80 east_output_space_count_f_reg_1_ (.o(east_output_space_count_f_1_),
	.ck(clk),
	.d(east_output_space_N43));
   ms00f80 east_output_space_is_one_f_reg (.o(east_output_space_is_one_f),
	.ck(clk),
	.d(east_output_space_N47));
   ms00f80 east_output_space_count_f_reg_0_ (.o(east_output_space_count_f_0_),
	.ck(clk),
	.d(east_output_space_N42));
   ms00f80 east_output_control_ec_wants_to_send_but_cannot_reg (.o(ec_wants_to_send_but_cannot_E),
	.ck(clk),
	.d(east_output_control_N72));
   ms00f80 ec_thanks_e_to_w_reg_reg (.o(ec_thanks_e_to_w_reg),
	.ck(clk),
	.d(n25994));
   ms00f80 west_input_control_thanks_all_f_reg (.o(west_input_control_thanks_all_f),
	.ck(clk),
	.d(n26013));
   ms00f80 west_input_NIB_yummy_out_f_reg (.o(yummyOut_W),
	.ck(clk),
	.d(n26013));
   ms00f80 west_input_NIB_elements_in_array_f_reg_0_ (.o(west_input_NIB_elements_in_array_f_0_),
	.ck(clk),
	.d(n25989));
   ms00f80 west_input_NIB_elements_in_array_f_reg_1_ (.o(west_input_NIB_elements_in_array_f_1_),
	.ck(clk),
	.d(n25988));
   ms00f80 west_input_NIB_elements_in_array_f_reg_2_ (.o(west_input_NIB_elements_in_array_f_2_),
	.ck(clk),
	.d(n2703));
   ms00f80 ec_west_input_valid_reg_reg (.o(ec_west_input_valid_reg),
	.ck(clk),
	.d(west_input_valid));
   ms00f80 west_input_NIB_head_ptr_f_reg_0_ (.o(west_input_NIB_head_ptr_f_0_),
	.ck(clk),
	.d(n2693));
   ms00f80 west_input_NIB_head_ptr_f_reg_1_ (.o(west_input_NIB_head_ptr_f_1_),
	.ck(clk),
	.d(n2688));
   ms00f80 west_input_control_count_zero_f_reg (.o(west_input_control_count_zero_f),
	.ck(clk),
	.d(west_input_control_N51));
   ms00f80 west_input_control_header_last_f_reg (.o(west_input_control_header_last_f),
	.ck(clk),
	.d(west_input_control_N49));
   ms00f80 west_input_control_count_f_reg_0_ (.o(west_input_control_count_f_0_),
	.ck(clk),
	.d(n26012));
   ms00f80 west_input_control_count_f_reg_1_ (.o(west_input_control_count_f_1_),
	.ck(clk),
	.d(west_input_control_N42));
   ms00f80 west_input_control_count_f_reg_2_ (.o(west_input_control_count_f_2_),
	.ck(clk),
	.d(west_input_control_N43));
   ms00f80 west_input_control_count_f_reg_3_ (.o(west_input_control_count_f_3_),
	.ck(clk),
	.d(west_input_control_N44));
   ms00f80 west_input_control_count_f_reg_4_ (.o(west_input_control_count_f_4_),
	.ck(clk),
	.d(west_input_control_N45));
   ms00f80 west_input_control_count_f_reg_5_ (.o(west_input_control_count_f_5_),
	.ck(clk),
	.d(west_input_control_N46));
   ms00f80 west_input_control_count_f_reg_6_ (.o(west_input_control_count_f_6_),
	.ck(clk),
	.d(west_input_control_N47));
   ms00f80 west_input_control_count_f_reg_7_ (.o(west_input_control_count_f_7_),
	.ck(clk),
	.d(west_input_control_N48));
   ms00f80 west_input_control_count_one_f_reg (.o(west_input_control_count_one_f),
	.ck(clk),
	.d(west_input_control_N52));
   ms00f80 west_input_control_tail_last_f_reg (.o(west_input_control_tail_last_f),
	.ck(clk),
	.d(west_input_control_N53));
   ms00f80 east_output_control_current_route_f_reg_1_ (.o(east_output_current_route_connection_1_),
	.ck(clk),
	.d(east_output_control_N468));
   ms00f80 east_output_control_current_route_f_reg_0_ (.o(east_output_current_route_connection_0_),
	.ck(clk),
	.d(n26000));
   ms00f80 ec_thanks_e_to_p_reg_reg (.o(ec_thanks_e_to_p_reg),
	.ck(clk),
	.d(n26025));
   ms00f80 east_output_control_current_route_f_reg_2_ (.o(east_output_current_route_connection_2_),
	.ck(clk),
	.d(east_output_control_N469));
   ms00f80 ec_thanks_e_to_e_reg_reg (.o(ec_thanks_e_to_e_reg),
	.ck(clk),
	.d(n25984));
   ms00f80 ec_thanks_e_to_n_reg_reg (.o(ec_thanks_e_to_n_reg),
	.ck(clk),
	.d(n26011));
   ms00f80 north_input_control_thanks_all_f_reg (.o(north_input_control_thanks_all_f),
	.ck(clk),
	.d(n26010));
   ms00f80 north_input_NIB_yummy_out_f_reg (.o(yummyOut_N),
	.ck(clk),
	.d(n26010));
   ms00f80 north_input_NIB_elements_in_array_f_reg_0_ (.o(north_input_NIB_elements_in_array_f_0_),
	.ck(clk),
	.d(n2583));
   ms00f80 north_input_NIB_elements_in_array_f_reg_1_ (.o(north_input_NIB_elements_in_array_f_1_),
	.ck(clk),
	.d(n2578));
   ms00f80 north_input_NIB_elements_in_array_f_reg_2_ (.o(north_input_NIB_elements_in_array_f_2_),
	.ck(clk),
	.d(n2573));
   ms00f80 ec_north_input_valid_reg_reg (.o(ec_north_input_valid_reg),
	.ck(clk),
	.d(north_input_valid));
   ms00f80 north_input_NIB_head_ptr_f_reg_0_ (.o(north_input_NIB_head_ptr_f_0_),
	.ck(clk),
	.d(n2563));
   ms00f80 north_input_NIB_head_ptr_f_reg_1_ (.o(north_input_NIB_head_ptr_f_1_),
	.ck(clk),
	.d(n2558));
   ms00f80 north_input_control_count_zero_f_reg (.o(north_input_control_count_zero_f),
	.ck(clk),
	.d(north_input_control_N51));
   ms00f80 north_input_control_header_last_f_reg (.o(north_input_control_header_last_f),
	.ck(clk),
	.d(north_input_control_N49));
   ms00f80 north_input_control_count_f_reg_0_ (.o(north_input_control_count_f_0_),
	.ck(clk),
	.d(n26009));
   ms00f80 north_input_control_count_f_reg_1_ (.o(north_input_control_count_f_1_),
	.ck(clk),
	.d(north_input_control_N42));
   ms00f80 north_input_control_count_f_reg_2_ (.o(north_input_control_count_f_2_),
	.ck(clk),
	.d(north_input_control_N43));
   ms00f80 north_input_control_count_f_reg_3_ (.o(north_input_control_count_f_3_),
	.ck(clk),
	.d(north_input_control_N44));
   ms00f80 north_input_control_count_f_reg_4_ (.o(north_input_control_count_f_4_),
	.ck(clk),
	.d(north_input_control_N45));
   ms00f80 north_input_control_count_f_reg_5_ (.o(north_input_control_count_f_5_),
	.ck(clk),
	.d(north_input_control_N46));
   ms00f80 north_input_control_count_f_reg_6_ (.o(north_input_control_count_f_6_),
	.ck(clk),
	.d(north_input_control_N47));
   ms00f80 north_input_control_count_f_reg_7_ (.o(north_input_control_count_f_7_),
	.ck(clk),
	.d(north_input_control_N48));
   ms00f80 north_input_control_count_one_f_reg (.o(north_input_control_count_one_f),
	.ck(clk),
	.d(north_input_control_N52));
   ms00f80 north_input_control_tail_last_f_reg (.o(north_input_control_tail_last_f),
	.ck(clk),
	.d(north_input_control_N53));
   ms00f80 south_output_space_valid_f_reg (.o(south_output_space_valid_f),
	.ck(clk),
	.d(south_output_space_N46));
   ms00f80 south_output_space_count_f_reg_2_ (.o(south_output_space_count_f_2_),
	.ck(clk),
	.d(south_output_space_N44));
   ms00f80 south_output_space_is_two_or_more_f_reg (.o(south_output_space_is_two_or_more_f),
	.ck(clk),
	.d(south_output_space_N48));
   ms00f80 south_output_space_count_f_reg_1_ (.o(south_output_space_count_f_1_),
	.ck(clk),
	.d(south_output_space_N43));
   ms00f80 south_output_space_is_one_f_reg (.o(south_output_space_is_one_f),
	.ck(clk),
	.d(south_output_space_N47));
   ms00f80 south_output_space_count_f_reg_0_ (.o(south_output_space_count_f_0_),
	.ck(clk),
	.d(south_output_space_N42));
   ms00f80 south_output_control_ec_wants_to_send_but_cannot_reg (.o(ec_wants_to_send_but_cannot_S),
	.ck(clk),
	.d(south_output_control_N72));
   ms00f80 ec_thanks_s_to_e_reg_reg (.o(ec_thanks_s_to_e_reg),
	.ck(clk),
	.d(n25997));
   ms00f80 east_input_control_thanks_all_f_reg (.o(east_input_control_thanks_all_f),
	.ck(clk),
	.d(n25993));
   ms00f80 east_input_NIB_yummy_out_f_reg (.o(yummyOut_E),
	.ck(clk),
	.d(n25993));
   ms00f80 east_input_NIB_elements_in_array_f_reg_0_ (.o(east_input_NIB_elements_in_array_f_0_),
	.ck(clk),
	.d(n2443));
   ms00f80 east_input_NIB_elements_in_array_f_reg_1_ (.o(east_input_NIB_elements_in_array_f_1_),
	.ck(clk),
	.d(n2438));
   ms00f80 east_input_NIB_elements_in_array_f_reg_2_ (.o(east_input_NIB_elements_in_array_f_2_),
	.ck(clk),
	.d(n2433));
   ms00f80 ec_east_input_valid_reg_reg (.o(ec_east_input_valid_reg),
	.ck(clk),
	.d(east_input_valid));
   ms00f80 east_input_NIB_head_ptr_f_reg_0_ (.o(east_input_NIB_head_ptr_f_0_),
	.ck(clk),
	.d(n2423));
   ms00f80 east_input_NIB_head_ptr_f_reg_1_ (.o(east_input_NIB_head_ptr_f_1_),
	.ck(clk),
	.d(n2418));
   ms00f80 east_input_control_count_zero_f_reg (.o(east_input_control_count_zero_f),
	.ck(clk),
	.d(east_input_control_N51));
   ms00f80 east_input_control_header_last_f_reg (.o(east_input_control_header_last_f),
	.ck(clk),
	.d(east_input_control_N49));
   ms00f80 east_input_control_count_f_reg_0_ (.o(east_input_control_count_f_0_),
	.ck(clk),
	.d(east_input_control_N41));
   ms00f80 east_input_control_count_f_reg_1_ (.o(east_input_control_count_f_1_),
	.ck(clk),
	.d(east_input_control_N42));
   ms00f80 east_input_control_count_f_reg_2_ (.o(east_input_control_count_f_2_),
	.ck(clk),
	.d(east_input_control_N43));
   ms00f80 east_input_control_count_f_reg_3_ (.o(east_input_control_count_f_3_),
	.ck(clk),
	.d(east_input_control_N44));
   ms00f80 east_input_control_count_f_reg_4_ (.o(east_input_control_count_f_4_),
	.ck(clk),
	.d(east_input_control_N45));
   ms00f80 east_input_control_count_f_reg_5_ (.o(east_input_control_count_f_5_),
	.ck(clk),
	.d(east_input_control_N46));
   ms00f80 east_input_control_count_f_reg_6_ (.o(east_input_control_count_f_6_),
	.ck(clk),
	.d(east_input_control_N47));
   ms00f80 east_input_control_count_f_reg_7_ (.o(east_input_control_count_f_7_),
	.ck(clk),
	.d(east_input_control_N48));
   ms00f80 east_input_control_count_one_f_reg (.o(east_input_control_count_one_f),
	.ck(clk),
	.d(east_input_control_N52));
   ms00f80 east_input_control_tail_last_f_reg (.o(east_input_control_tail_last_f),
	.ck(clk),
	.d(east_input_control_N53));
   ms00f80 proc_output_control_current_route_f_reg_1_ (.o(proc_output_current_route_connection_1_),
	.ck(clk),
	.d(proc_output_control_N468));
   ms00f80 ec_thanks_p_to_s_reg_reg (.o(ec_thanks_p_to_s_reg),
	.ck(clk),
	.d(n25986));
   ms00f80 proc_output_control_current_route_f_reg_0_ (.o(proc_output_current_route_connection_0_),
	.ck(clk),
	.d(proc_output_control_N467));
   ms00f80 ec_thanks_p_to_n_reg_reg (.o(ec_thanks_p_to_n_reg),
	.ck(clk),
	.d(n26028));
   ms00f80 ec_thanks_p_to_e_reg_reg (.o(ec_thanks_p_to_e_reg),
	.ck(clk),
	.d(n26008));
   ms00f80 ec_thanks_p_to_w_reg_reg (.o(ec_thanks_p_to_w_reg),
	.ck(clk),
	.d(n25987));
   ms00f80 proc_output_control_planned_f_reg (.o(proc_output_control_planned_f),
	.ck(clk),
	.d(proc_output_control_N470));
   ms00f80 south_output_control_current_route_f_reg_2_ (.o(south_output_current_route_connection_2_),
	.ck(clk),
	.d(south_output_control_N469));
   ms00f80 south_output_control_current_route_f_reg_1_ (.o(south_output_current_route_connection_1_),
	.ck(clk),
	.d(south_output_control_N468));
   ms00f80 south_output_control_current_route_f_reg_0_ (.o(south_output_current_route_connection_0_),
	.ck(clk),
	.d(south_output_control_N467));
   ms00f80 ec_thanks_s_to_n_reg_reg (.o(ec_thanks_s_to_n_reg),
	.ck(clk),
	.d(n25999));
   ms00f80 south_output_control_planned_f_reg (.o(south_output_control_planned_f),
	.ck(clk),
	.d(south_output_control_N470));
   ms00f80 north_output_control_current_route_f_reg_2_ (.o(north_output_current_route_connection_2_),
	.ck(clk),
	.d(north_output_control_N469));
   ms00f80 ec_thanks_n_to_n_reg_reg (.o(ec_thanks_n_to_n_reg),
	.ck(clk),
	.d(n26022));
   ms00f80 north_output_control_current_route_f_reg_1_ (.o(north_output_current_route_connection_1_),
	.ck(clk),
	.d(north_output_control_N468));
   ms00f80 ec_thanks_n_to_s_reg_reg (.o(ec_thanks_n_to_s_reg),
	.ck(clk),
	.d(n26024));
   ms00f80 north_output_control_current_route_f_reg_0_ (.o(north_output_current_route_connection_0_),
	.ck(clk),
	.d(north_output_control_N467));
   ms00f80 ec_thanks_n_to_e_reg_reg (.o(ec_thanks_n_to_e_reg),
	.ck(clk),
	.d(n25985));
   ms00f80 ec_thanks_n_to_w_reg_reg (.o(ec_thanks_n_to_w_reg),
	.ck(clk),
	.d(n26021));
   ms00f80 north_output_control_planned_f_reg (.o(north_output_control_planned_f),
	.ck(clk),
	.d(north_output_control_N470));
   ms00f80 west_output_space_valid_f_reg (.o(west_output_space_valid_f),
	.ck(clk),
	.d(west_output_space_N46));
   ms00f80 west_output_space_count_f_reg_2_ (.o(west_output_space_count_f_2_),
	.ck(clk),
	.d(west_output_space_N44));
   ms00f80 west_output_space_is_two_or_more_f_reg (.o(west_output_space_is_two_or_more_f),
	.ck(clk),
	.d(west_output_space_N48));
   ms00f80 west_output_space_count_f_reg_1_ (.o(west_output_space_count_f_1_),
	.ck(clk),
	.d(west_output_space_N43));
   ms00f80 west_output_space_is_one_f_reg (.o(west_output_space_is_one_f),
	.ck(clk),
	.d(west_output_space_N47));
   ms00f80 west_output_space_count_f_reg_0_ (.o(west_output_space_count_f_0_),
	.ck(clk),
	.d(west_output_space_N42));
   ms00f80 west_output_control_ec_wants_to_send_but_cannot_reg (.o(ec_wants_to_send_but_cannot_W),
	.ck(clk),
	.d(west_output_control_N72));
   ms00f80 west_output_control_current_route_f_reg_2_ (.o(west_output_current_route_connection_2_),
	.ck(clk),
	.d(west_output_control_N469));
   ms00f80 west_output_control_current_route_f_reg_1_ (.o(west_output_current_route_connection_1_),
	.ck(clk),
	.d(west_output_control_N468));
   ms00f80 west_output_control_current_route_f_reg_0_ (.o(west_output_current_route_connection_0_),
	.ck(clk),
	.d(west_output_control_N467));
   ms00f80 west_output_control_planned_f_reg (.o(west_output_control_planned_f),
	.ck(clk),
	.d(west_output_control_N470));
   ms00f80 ec_thanks_w_to_n_reg_reg (.o(ec_thanks_w_to_n_reg),
	.ck(clk),
	.d(n26018));
   ms00f80 ec_thanks_w_to_e_reg_reg (.o(ec_thanks_w_to_e_reg),
	.ck(clk),
	.d(n25998));
   ms00f80 ec_thanks_w_to_w_reg_reg (.o(ec_thanks_w_to_w_reg),
	.ck(clk),
	.d(n26017));
   ms00f80 ec_thanks_w_to_p_reg_reg (.o(ec_thanks_w_to_p_reg),
	.ck(clk),
	.d(n26019));
   ms00f80 ec_thanks_w_to_s_reg_reg (.o(ec_thanks_w_to_s_reg),
	.ck(clk),
	.d(n26020));
   ms00f80 ec_thanks_s_to_w_reg_reg (.o(ec_thanks_s_to_w_reg),
	.ck(clk),
	.d(n26014));
   ms00f80 ec_thanks_s_to_p_reg_reg (.o(ec_thanks_s_to_p_reg),
	.ck(clk),
	.d(n26016));
   ms00f80 ec_thanks_s_to_s_reg_reg (.o(ec_thanks_s_to_s_reg),
	.ck(clk),
	.d(n26015));
   ms00f80 east_output_control_planned_f_reg (.o(east_output_control_planned_f),
	.ck(clk),
	.d(n26003));
   ms00f80 ec_thanks_e_to_s_reg_reg (.o(ec_thanks_e_to_s_reg),
	.ck(clk),
	.d(n25992));
   ms00f80 proc_output_control_ec_wants_to_send_but_cannot_reg (.o(ec_wants_to_send_but_cannot_P),
	.ck(clk),
	.d(proc_output_control_N72));
   ms00f80 REG_reset_fin_q_reg_0_ (.o(reset),
	.ck(clk),
	.d(reset_in));
   oa12m01 U18136 (.o(n11178),
	.a(n24782),
	.b(FE_OFN555_n24761),
	.c(n24783));
   oa12m01 U18137 (.o(n11138),
	.a(n24764),
	.b(FE_OFN555_n24761),
	.c(n24765));
   oa12m01 U18138 (.o(n11788),
	.a(n25201),
	.b(n24921),
	.c(n25202));
   oa12m01 U18139 (.o(n11823),
	.a(n25203),
	.b(FE_OFN943_n24921),
	.c(n25204));
   oa12m01 U18140 (.o(n11928),
	.a(n25221),
	.b(n24921),
	.c(n25222));
   oa12m01 U18141 (.o(n11933),
	.a(n25223),
	.b(n24921),
	.c(n25224));
   oa12m01 U18142 (.o(n11938),
	.a(n25219),
	.b(n24921),
	.c(n25220));
   oa12m01 U18143 (.o(n11953),
	.a(n25264),
	.b(n24921),
	.c(n25265));
   oa12m01 U18144 (.o(n11958),
	.a(n25256),
	.b(n24921),
	.c(n25257));
   oa12m01 U18145 (.o(n11963),
	.a(n25262),
	.b(n24921),
	.c(n25263));
   oa12m01 U18146 (.o(n11778),
	.a(n25217),
	.b(FE_OFN943_n24921),
	.c(n25218));
   oa12m01 U18147 (.o(n11803),
	.a(n25205),
	.b(n24921),
	.c(n25206));
   oa12m01 U18148 (.o(n11883),
	.a(n25189),
	.b(n24921),
	.c(n25190));
   oa12m01 U18149 (.o(n11943),
	.a(n25258),
	.b(n24921),
	.c(n25259));
   oa12m01 U18150 (.o(n11948),
	.a(n25266),
	.b(n24921),
	.c(n25267));
   oa12m01 U18151 (.o(n11973),
	.a(n25254),
	.b(n24921),
	.c(n25255));
   oa12m01 U18152 (.o(n11978),
	.a(n25252),
	.b(n24921),
	.c(n25253));
   oa12m01 U18153 (.o(n11818),
	.a(n25209),
	.b(n24921),
	.c(n25210));
   oa12m01 U18154 (.o(n11893),
	.a(n24932),
	.b(n24921),
	.c(n24933));
   oa12m01 U18155 (.o(n11968),
	.a(n25260),
	.b(n24921),
	.c(n25261));
   oa12m01 U18156 (.o(n11783),
	.a(n25207),
	.b(FE_OFN943_n24921),
	.c(n25208));
   oa12m01 U18157 (.o(n11773),
	.a(n25197),
	.b(FE_OFN943_n24921),
	.c(n25198));
   oa12m01 U18158 (.o(n11793),
	.a(n25191),
	.b(FE_OFN943_n24921),
	.c(n25192));
   oa12m01 U18159 (.o(n11798),
	.a(n25193),
	.b(FE_OFN943_n24921),
	.c(n25194));
   oa12m01 U18160 (.o(n11808),
	.a(n25215),
	.b(FE_OFN943_n24921),
	.c(n25216));
   oa12m01 U18161 (.o(n11833),
	.a(n25213),
	.b(FE_OFN943_n24921),
	.c(n25214));
   oa12m01 U18162 (.o(n11838),
	.a(n25211),
	.b(FE_OFN943_n24921),
	.c(n25212));
   oa12m01 U18163 (.o(n11813),
	.a(n25195),
	.b(FE_OFN943_n24921),
	.c(n25196));
   oa12m01 U18164 (.o(n11828),
	.a(n25199),
	.b(FE_OFN943_n24921),
	.c(n25200));
   oa12m01 U18165 (.o(n11643),
	.a(n22996),
	.b(n25263),
	.c(n22958));
   oa12m01 U18166 (.o(n11638),
	.a(n22995),
	.b(n25257),
	.c(n22958));
   oa12m01 U18167 (.o(n11658),
	.a(n23002),
	.b(n25253),
	.c(n22958));
   oa12m01 U18168 (.o(n11648),
	.a(n22997),
	.b(n25261),
	.c(n22958));
   oa12m01 U18169 (.o(n11653),
	.a(n23000),
	.b(n25255),
	.c(n22958));
   oa12m01 U18170 (.o(n11593),
	.a(n22986),
	.b(n22958),
	.c(n24939));
   oa12m01 U18171 (.o(n11588),
	.a(n22989),
	.b(n24943),
	.c(n22958));
   oa12m01 U18172 (.o(n10913),
	.a(n22953),
	.b(n24923),
	.c(FE_OFN24847_n22945));
   oa12m01 U18173 (.o(n10998),
	.a(n22981),
	.b(FE_OFN24857_n22945),
	.c(n25257));
   oa12m01 U18174 (.o(n11003),
	.a(n23011),
	.b(FE_OFN24860_n22945),
	.c(n25263));
   oa12m01 U18175 (.o(n11008),
	.a(n23016),
	.b(FE_OFN24844_n22945),
	.c(n25261));
   oa12m01 U18176 (.o(n11013),
	.a(n23015),
	.b(FE_OFN24844_n22945),
	.c(n25255));
   oa12m01 U18177 (.o(n11018),
	.a(n23014),
	.b(FE_OFN24844_n22945),
	.c(n25253));
   oa12m01 U18178 (.o(n10918),
	.a(n22954),
	.b(FE_OFN24848_n22945),
	.c(n24937));
   ao22m01 U18179 (.o(n11743),
	.a(FE_OFN435_n22958),
	.b(n25890),
	.c(n25873),
	.d(FE_OFN24810_n22958));
   ao22m01 U18180 (.o(n11753),
	.a(FE_OFN435_n22958),
	.b(n25888),
	.c(n25872),
	.d(FE_OFN24815_n22958));
   ao22m01 U18181 (.o(n11758),
	.a(FE_OFN435_n22958),
	.b(n25886),
	.c(n25871),
	.d(FE_OFN24811_n22958));
   ao22m01 U18182 (.o(n11768),
	.a(FE_OFN435_n22958),
	.b(n25884),
	.c(n25870),
	.d(FE_OFN24813_n22958));
   ao22m01 U18183 (.o(n11103),
	.a(FE_OFN24862_n22945),
	.b(n25890),
	.c(n25889),
	.d(FE_OFN24861_n22945));
   ao22m01 U18184 (.o(n11113),
	.a(FE_OFN24862_n22945),
	.b(n25888),
	.c(n25887),
	.d(FE_OFN24861_n22945));
   ao22m01 U18185 (.o(n11118),
	.a(FE_OFN24862_n22945),
	.b(n25886),
	.c(n25885),
	.d(FE_OFN24861_n22945));
   ao22m01 U18186 (.o(n11128),
	.a(FE_OFN24862_n22945),
	.b(n25884),
	.c(n25883),
	.d(FE_OFN24861_n22945));
   ao12m01 U18187 (.o(west_input_control_N45),
	.a(FE_OFN25647_reset),
	.b(n20730),
	.c(n20729));
   na03s01 U18188 (.o(n13383),
	.a(FE_OFN88_n21220),
	.b(FE_OFN1087_n20656),
	.c(n25831));
   oa12m01 U18189 (.o(n13268),
	.a(n21179),
	.b(n25836),
	.c(n21226));
   oa12m01 U18190 (.o(n13263),
	.a(n21210),
	.b(n25836),
	.c(n21222));
   oa12m01 U18191 (.o(n13238),
	.a(n21211),
	.b(n25836),
	.c(n21243));
   oa12m01 U18192 (.o(n13243),
	.a(n21203),
	.b(n25836),
	.c(n21250));
   oa12m01 U18193 (.o(n13258),
	.a(n21207),
	.b(n25836),
	.c(n21224));
   oa12m01 U18194 (.o(n13093),
	.a(n21176),
	.b(FE_OFN86_n21175),
	.c(n21274));
   oa12m01 U18195 (.o(n13168),
	.a(n21199),
	.b(n25836),
	.c(n22650));
   oa12m01 U18196 (.o(n13088),
	.a(n21185),
	.b(FE_OFN86_n21175),
	.c(n21256));
   oa12m01 U18197 (.o(n13163),
	.a(n21198),
	.b(n25836),
	.c(n22630));
   oa12m01 U18198 (.o(n12618),
	.a(n21223),
	.b(FE_OFN88_n21220),
	.c(n21224));
   oa12m01 U18199 (.o(n12533),
	.a(n21263),
	.b(FE_OFN88_n21220),
	.c(n21264));
   oa12m01 U18200 (.o(n12538),
	.a(n21261),
	.b(FE_OFN88_n21220),
	.c(n21262));
   oa12m01 U18201 (.o(n12583),
	.a(n21236),
	.b(FE_OFN88_n21220),
	.c(n21237));
   oa12m01 U18202 (.o(n12588),
	.a(n21258),
	.b(FE_OFN88_n21220),
	.c(n21259));
   oa12m01 U18203 (.o(n12593),
	.a(n21247),
	.b(FE_OFN88_n21220),
	.c(n21248));
   oa12m01 U18204 (.o(n12608),
	.a(n21265),
	.b(FE_OFN88_n21220),
	.c(n21266));
   oa12m01 U18205 (.o(n12628),
	.a(n21225),
	.b(FE_OFN88_n21220),
	.c(n21226));
   oa12m01 U18206 (.o(n12488),
	.a(n21281),
	.b(FE_OFN88_n21220),
	.c(n21282));
   oa12m01 U18207 (.o(n12498),
	.a(n21267),
	.b(FE_OFN88_n21220),
	.c(n22652));
   oa12m01 U18208 (.o(n12503),
	.a(n21233),
	.b(FE_OFN88_n21220),
	.c(n21234));
   oa12m01 U18209 (.o(n12578),
	.a(n21230),
	.b(FE_OFN88_n21220),
	.c(n22640));
   oa12m01 U18210 (.o(n12598),
	.a(n21242),
	.b(FE_OFN88_n21220),
	.c(n21243));
   oa12m01 U18211 (.o(n12613),
	.a(n21231),
	.b(FE_OFN88_n21220),
	.c(n21232));
   oa12m01 U18212 (.o(n12623),
	.a(n21221),
	.b(FE_OFN88_n21220),
	.c(n21222));
   oa12m01 U18213 (.o(n12543),
	.a(n21228),
	.b(FE_OFN88_n21220),
	.c(n22646));
   oa12m01 U18214 (.o(n12513),
	.a(n21275),
	.b(FE_OFN88_n21220),
	.c(n22632));
   oa12m01 U18215 (.o(n12568),
	.a(n21260),
	.b(FE_OFN88_n21220),
	.c(n22648));
   oa12m01 U18216 (.o(n12603),
	.a(n21249),
	.b(FE_OFN88_n21220),
	.c(n21250));
   oa12m01 U18217 (.o(n12508),
	.a(n21244),
	.b(FE_OFN88_n21220),
	.c(n22636));
   oa12m01 U18218 (.o(n12528),
	.a(n21235),
	.b(FE_OFN88_n21220),
	.c(n22650));
   oa12m01 U18219 (.o(n12553),
	.a(n21257),
	.b(FE_OFN88_n21220),
	.c(n22654));
   oa12m01 U18220 (.o(n12493),
	.a(n21278),
	.b(FE_OFN88_n21220),
	.c(n22634));
   oa12m01 U18221 (.o(n12548),
	.a(n21268),
	.b(FE_OFN88_n21220),
	.c(n22638));
   oa12m01 U18222 (.o(n12558),
	.a(n21227),
	.b(FE_OFN88_n21220),
	.c(n22656));
   oa12m01 U18223 (.o(n12423),
	.a(n21240),
	.b(n25848),
	.c(n21241));
   oa12m01 U18224 (.o(n12428),
	.a(n21245),
	.b(n25848),
	.c(n21246));
   oa12m01 U18225 (.o(n12448),
	.a(n21255),
	.b(n25848),
	.c(n21256));
   oa12m01 U18226 (.o(n12453),
	.a(n21273),
	.b(n25848),
	.c(n21274));
   oa12m01 U18227 (.o(n12458),
	.a(n21276),
	.b(n25848),
	.c(n21277));
   oa12m01 U18228 (.o(n12463),
	.a(n21253),
	.b(n25848),
	.c(n21254));
   oa12m01 U18229 (.o(n12518),
	.a(n21271),
	.b(FE_OFN88_n21220),
	.c(n21272));
   oa12m01 U18230 (.o(n12523),
	.a(n21283),
	.b(FE_OFN88_n21220),
	.c(n22630));
   oa12m01 U18231 (.o(n12563),
	.a(n21252),
	.b(FE_OFN88_n21220),
	.c(n22644));
   oa12m01 U18232 (.o(n12468),
	.a(n21269),
	.b(n25848),
	.c(n21270));
   oa12m01 U18233 (.o(n12443),
	.a(n21251),
	.b(n25848),
	.c(n22642));
   oa12m01 U18234 (.o(n12433),
	.a(n21229),
	.b(n25848),
	.c(n22444));
   oa12m01 U18235 (.o(n12473),
	.a(n21284),
	.b(FE_OFN88_n21220),
	.c(n21285));
   oa12m01 U18236 (.o(n12478),
	.a(n21279),
	.b(n25848),
	.c(n21280));
   oa12m01 U18237 (.o(n12483),
	.a(n21238),
	.b(n25848),
	.c(n21239));
   oa12m01 U18238 (.o(n12438),
	.a(n21286),
	.b(n25848),
	.c(n21287));
   ao22m01 U18239 (.o(n13348),
	.a(n21175),
	.b(n25851),
	.c(n25832),
	.d(FE_OFN86_n21175));
   ao22m01 U18240 (.o(n12643),
	.a(n21220),
	.b(n25857),
	.c(n25847),
	.d(n25848));
   oa12m01 U18241 (.o(n9073),
	.a(n22708),
	.b(n21053),
	.c(n22745));
   oa12m01 U18242 (.o(n9028),
	.a(n22709),
	.b(FE_OFN25792_n21053),
	.c(n22749));
   oa12m01 U18243 (.o(n9053),
	.a(n22707),
	.b(n21053),
	.c(n22728));
   oa12m01 U18244 (.o(n8963),
	.a(n21064),
	.b(n21101),
	.c(FE_OFN25792_n21053));
   oa12m01 U18245 (.o(n9003),
	.a(n21078),
	.b(FE_OFN25792_n21053),
	.c(n21115));
   oa12m01 U18246 (.o(n9013),
	.a(n21062),
	.b(FE_OFN25792_n21053),
	.c(n21119));
   oa12m01 U18247 (.o(n9033),
	.a(n22713),
	.b(FE_OFN25792_n21053),
	.c(n22714));
   oa12m01 U18248 (.o(n9038),
	.a(n22746),
	.b(FE_OFN25792_n21053),
	.c(n22747));
   oa12m01 U18249 (.o(n9048),
	.a(n22711),
	.b(n22712),
	.c(n21053));
   oa12m01 U18250 (.o(n9058),
	.a(n21067),
	.b(n21053),
	.c(n22751));
   oa12m01 U18251 (.o(n9063),
	.a(n22725),
	.b(n21053),
	.c(n22726));
   oa12m01 U18252 (.o(n9068),
	.a(n22715),
	.b(n21053),
	.c(n22736));
   oa12m01 U18253 (.o(n9078),
	.a(n22721),
	.b(n22732),
	.c(n21053));
   oa12m01 U18254 (.o(n8968),
	.a(n22485),
	.b(FE_OFN25792_n21053),
	.c(n22486));
   oa12m01 U18255 (.o(n9043),
	.a(n21066),
	.b(n21053),
	.c(n22739));
   oa12m01 U18256 (.o(n9018),
	.a(n21065),
	.b(n21121),
	.c(FE_OFN25794_n21053));
   oa12m01 U18257 (.o(n9008),
	.a(n21059),
	.b(n21053),
	.c(n21117));
   oa12m01 U18258 (.o(n8893),
	.a(n22733),
	.b(n22734),
	.c(FE_OFN25792_n21053));
   oa12m01 U18259 (.o(n8873),
	.a(n21061),
	.b(FE_OFN25791_n21053),
	.c(n21072));
   oa12m01 U18260 (.o(n8998),
	.a(n21060),
	.b(FE_OFN25794_n21053),
	.c(n21113));
   oa12m01 U18261 (.o(n8888),
	.a(n21054),
	.b(FE_OFN25791_n21053),
	.c(n21097));
   oa12m01 U18262 (.o(n12913),
	.a(n20666),
	.b(FE_OFN1087_n20656),
	.c(n21248));
   oa12m01 U18263 (.o(n12853),
	.a(n20668),
	.b(FE_OFN1087_n20656),
	.c(n21264));
   oa12m01 U18264 (.o(n12858),
	.a(n20692),
	.b(FE_OFN1087_n20656),
	.c(n21262));
   oa12m01 U18265 (.o(n12903),
	.a(n20679),
	.b(FE_OFN1087_n20656),
	.c(n21237));
   oa12m01 U18266 (.o(n12908),
	.a(n20693),
	.b(FE_OFN1087_n20656),
	.c(n21259));
   oa12m01 U18267 (.o(n12928),
	.a(n20684),
	.b(FE_OFN1087_n20656),
	.c(n21266));
   oa12m01 U18268 (.o(n12948),
	.a(n20690),
	.b(FE_OFN1087_n20656),
	.c(n21226));
   oa12m01 U18269 (.o(n12808),
	.a(n20661),
	.b(FE_OFN1087_n20656),
	.c(n21282));
   oa12m01 U18270 (.o(n12818),
	.a(n20688),
	.b(FE_OFN1087_n20656),
	.c(n22652));
   oa12m01 U18271 (.o(n12823),
	.a(n20689),
	.b(FE_OFN1087_n20656),
	.c(n21234));
   oa12m01 U18272 (.o(n12898),
	.a(n20678),
	.b(FE_OFN1087_n20656),
	.c(n22640));
   oa12m01 U18273 (.o(n12918),
	.a(n20682),
	.b(FE_OFN1087_n20656),
	.c(n21243));
   oa12m01 U18274 (.o(n12933),
	.a(n20671),
	.b(FE_OFN1087_n20656),
	.c(n21232));
   oa12m01 U18275 (.o(n12938),
	.a(n20694),
	.b(FE_OFN1087_n20656),
	.c(n21224));
   oa12m01 U18276 (.o(n12943),
	.a(n20695),
	.b(FE_OFN1087_n20656),
	.c(n21222));
   oa12m01 U18277 (.o(n12833),
	.a(n20687),
	.b(FE_OFN1087_n20656),
	.c(n22632));
   oa12m01 U18278 (.o(n12888),
	.a(n20675),
	.b(FE_OFN1087_n20656),
	.c(n22648));
   oa12m01 U18279 (.o(n12923),
	.a(n20683),
	.b(FE_OFN1087_n20656),
	.c(n21250));
   oa12m01 U18280 (.o(n12828),
	.a(n20662),
	.b(FE_OFN1087_n20656),
	.c(n22636));
   oa12m01 U18281 (.o(n12848),
	.a(n20676),
	.b(FE_OFN1087_n20656),
	.c(n22650));
   oa12m01 U18282 (.o(n12873),
	.a(n20669),
	.b(FE_OFN1087_n20656),
	.c(n22654));
   oa12m01 U18283 (.o(n12868),
	.a(n20680),
	.b(FE_OFN1087_n20656),
	.c(n22638));
   oa12m01 U18284 (.o(n12878),
	.a(n20672),
	.b(FE_OFN1087_n20656),
	.c(n22656));
   oa12m01 U18285 (.o(n12838),
	.a(n20674),
	.b(FE_OFN1087_n20656),
	.c(n21272));
   oa12m01 U18286 (.o(n12743),
	.a(n20685),
	.b(FE_OFN25876_n25842),
	.c(n21241));
   oa12m01 U18287 (.o(n12748),
	.a(n20691),
	.b(FE_OFN25876_n25842),
	.c(n21246));
   oa12m01 U18288 (.o(n12768),
	.a(n20670),
	.b(FE_OFN25876_n25842),
	.c(n21256));
   oa12m01 U18289 (.o(n12773),
	.a(n20659),
	.b(FE_OFN25876_n25842),
	.c(n21274));
   oa12m01 U18290 (.o(n12778),
	.a(n20657),
	.b(FE_OFN25876_n25842),
	.c(n21277));
   oa12m01 U18291 (.o(n12783),
	.a(n20663),
	.b(FE_OFN25876_n25842),
	.c(n21254));
   oa12m01 U18292 (.o(n12813),
	.a(n20667),
	.b(FE_OFN1087_n20656),
	.c(n22634));
   oa12m01 U18293 (.o(n12843),
	.a(n20660),
	.b(FE_OFN1087_n20656),
	.c(n22630));
   oa12m01 U18294 (.o(n12863),
	.a(n20664),
	.b(FE_OFN1087_n20656),
	.c(n22646));
   oa12m01 U18295 (.o(n12883),
	.a(n20673),
	.b(FE_OFN1087_n20656),
	.c(n22644));
   oa12m01 U18296 (.o(n12763),
	.a(n20686),
	.b(FE_OFN25876_n25842),
	.c(n22642));
   oa12m01 U18297 (.o(n12753),
	.a(n20681),
	.b(FE_OFN25876_n25842),
	.c(n22444));
   oa12m01 U18298 (.o(n12788),
	.a(n20665),
	.b(FE_OFN25876_n25842),
	.c(n21270));
   oa12m01 U18299 (.o(n12793),
	.a(n20697),
	.b(FE_OFN1087_n20656),
	.c(n21285));
   oa12m01 U18300 (.o(n12798),
	.a(n20658),
	.b(FE_OFN25876_n25842),
	.c(n21280));
   oa12m01 U18301 (.o(n12803),
	.a(n20677),
	.b(FE_OFN25876_n25842),
	.c(n21239));
   oa12m01 U18302 (.o(n12758),
	.a(n20696),
	.b(FE_OFN25876_n25842),
	.c(n21287));
   ao12m01 U18303 (.o(south_input_control_N43),
	.a(FE_OFN5_reset),
	.b(n20640),
	.c(n20639));
   oa12m01 U18304 (.o(n7573),
	.a(n22021),
	.b(FE_OFN25741_FE_OFN25605_n21944),
	.c(n23827));
   oa12m01 U18305 (.o(n7018),
	.a(n21912),
	.b(n21911),
	.c(n23916));
   oa12m01 U18306 (.o(n6043),
	.a(n22191),
	.b(FE_OFN101_n22098),
	.c(n23908));
   oa12m01 U18307 (.o(n6118),
	.a(n22206),
	.b(FE_OFN101_n22098),
	.c(n23816));
   oa12m01 U18308 (.o(n6933),
	.a(n21954),
	.b(FE_OFN25628_n21910),
	.c(n23827));
   oa12m01 U18309 (.o(n6943),
	.a(n21962),
	.b(FE_OFN25628_n21910),
	.c(n23918));
   oa12m01 U18310 (.o(n7768),
	.a(n21978),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23798));
   oa12m01 U18311 (.o(n7693),
	.a(n21993),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23934));
   oa12m01 U18312 (.o(n5973),
	.a(n22129),
	.b(FE_OFN465_n23476),
	.c(n23827));
   oa12m01 U18313 (.o(n7318),
	.a(n21924),
	.b(FE_OFN25781_FE_OFN448_n23236),
	.c(n23903));
   oa12m01 U18314 (.o(n7393),
	.a(n22033),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23944));
   oa12m01 U18315 (.o(n5818),
	.a(n22120),
	.b(n22085),
	.c(n23894));
   oa12m01 U18316 (.o(n6493),
	.a(n22142),
	.b(FE_OFN103_n22140),
	.c(n23793));
   oa12m01 U18317 (.o(n7618),
	.a(n21998),
	.b(FE_OFN25741_FE_OFN25605_n21944),
	.c(n23924));
   oa12m01 U18318 (.o(n7733),
	.a(n21986),
	.b(FE_OFN25605_n21944),
	.c(n23791));
   oa12m01 U18319 (.o(n6293),
	.a(n22185),
	.b(FE_OFN103_n22140),
	.c(n23827));
   oa12m01 U18320 (.o(n6343),
	.a(n22173),
	.b(FE_OFN103_n22140),
	.c(n23922));
   oa12m01 U18321 (.o(n6418),
	.a(n22158),
	.b(FE_OFN103_n22140),
	.c(n23812));
   oa12m01 U18322 (.o(n7253),
	.a(n21926),
	.b(FE_OFN25781_FE_OFN448_n23236),
	.c(n23827));
   oa12m01 U18323 (.o(n5743),
	.a(n22103),
	.b(n22085),
	.c(n23942));
   oa12m01 U18324 (.o(n5653),
	.a(n22156),
	.b(n23471),
	.c(n23827));
   oa12m01 U18325 (.o(n5668),
	.a(n22086),
	.b(n23471),
	.c(n23926));
   oa12m01 U18326 (.o(n6133),
	.a(n22213),
	.b(FE_OFN465_n23476),
	.c(n23791));
   oa12m01 U18327 (.o(n6168),
	.a(n22180),
	.b(FE_OFN101_n22098),
	.c(n23798));
   oa12m01 U18328 (.o(n7093),
	.a(n21965),
	.b(FE_OFN25627_n21910),
	.c(n23791));
   oa12m01 U18329 (.o(n7128),
	.a(n21948),
	.b(FE_OFN25626_n21910),
	.c(n23798));
   oa12m01 U18330 (.o(n7413),
	.a(n22036),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23791));
   oa12m01 U18331 (.o(n7448),
	.a(n22002),
	.b(n23236),
	.c(n23798));
   oa12m01 U18332 (.o(n6093),
	.a(n22192),
	.b(FE_OFN465_n23476),
	.c(n23934));
   oa12m01 U18333 (.o(n7053),
	.a(n21961),
	.b(FE_OFN913_n23246),
	.c(n23934));
   oa12m01 U18334 (.o(n7373),
	.a(n22011),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23934));
   oa12m01 U18335 (.o(n6018),
	.a(n22186),
	.b(FE_OFN465_n23476),
	.c(n23924));
   oa12m01 U18336 (.o(n7298),
	.a(n21917),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23924));
   oa12m01 U18337 (.o(n6978),
	.a(n21951),
	.b(FE_OFN25627_n21910),
	.c(n23924));
   oa12m01 U18338 (.o(n5848),
	.a(n22126),
	.b(n22085),
	.c(n23798));
   oa12m01 U18339 (.o(n6488),
	.a(n22143),
	.b(n23453),
	.c(n23798));
   oa12m01 U18340 (.o(n5773),
	.a(n22109),
	.b(n22085),
	.c(n23934));
   oa12m01 U18341 (.o(n5813),
	.a(n22119),
	.b(n23471),
	.c(n23791));
   oa12m01 U18342 (.o(n6413),
	.a(n22159),
	.b(FE_OFN103_n22140),
	.c(n23934));
   oa12m01 U18343 (.o(n6453),
	.a(n22150),
	.b(FE_OFN103_n22140),
	.c(n23791));
   oa12m01 U18344 (.o(n6338),
	.a(n22174),
	.b(FE_OFN103_n22140),
	.c(n23924));
   oa12m01 U18345 (.o(n5698),
	.a(n22092),
	.b(n23471),
	.c(n23924));
   oa12m01 U18346 (.o(n10308),
	.a(n20989),
	.b(FE_OFN84_n20972),
	.c(n22667));
   oa12m01 U18347 (.o(n10363),
	.a(n21002),
	.b(FE_OFN84_n20972),
	.c(n21046));
   oa12m01 U18348 (.o(n10368),
	.a(n21003),
	.b(FE_OFN84_n20972),
	.c(n21028));
   oa12m01 U18349 (.o(n10353),
	.a(n21000),
	.b(FE_OFN84_n20972),
	.c(n21009));
   oa12m01 U18350 (.o(n10358),
	.a(n21001),
	.b(FE_OFN84_n20972),
	.c(n21044));
   oa12m01 U18351 (.o(n10318),
	.a(n22701),
	.b(FE_OFN84_n20972),
	.c(n22702));
   oa12m01 U18352 (.o(n10238),
	.a(n22678),
	.b(FE_OFN84_n20972),
	.c(n22679));
   oa12m01 U18353 (.o(n10243),
	.a(n22703),
	.b(n22704),
	.c(FE_OFN84_n20972));
   oa12m01 U18354 (.o(n10168),
	.a(n20984),
	.b(n25905),
	.c(n21007));
   oa12m01 U18355 (.o(n10163),
	.a(n20973),
	.b(n25905),
	.c(n22686));
   oa12m01 U18356 (.o(n9353),
	.a(n21122),
	.b(FE_OFN25866_FE_OFN24766_n21069),
	.c(n22714));
   oa12m01 U18357 (.o(n9373),
	.a(n22727),
	.b(n22728),
	.c(FE_OFN25865_FE_OFN24766_n21069));
   oa12m01 U18358 (.o(n9263),
	.a(n21090),
	.b(n21091),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   oa12m01 U18359 (.o(n9268),
	.a(n21098),
	.b(n21099),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   oa12m01 U18360 (.o(n9348),
	.a(n22748),
	.b(n22749),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   oa12m01 U18361 (.o(n9368),
	.a(n22710),
	.b(FE_OFN25862_FE_OFN24766_n21069),
	.c(n22712));
   oa12m01 U18362 (.o(n9378),
	.a(n22750),
	.b(n22751),
	.c(FE_OFN24766_n21069));
   oa12m01 U18363 (.o(n9383),
	.a(n21123),
	.b(n22726),
	.c(FE_OFN24766_n21069));
   oa12m01 U18364 (.o(n9398),
	.a(n22731),
	.b(FE_OFN25866_FE_OFN24766_n21069),
	.c(n22732));
   oa12m01 U18365 (.o(n9193),
	.a(n21071),
	.b(n21072),
	.c(FE_OFN24767_n21069));
   ao22m01 U18366 (.o(n13028),
	.a(n20656),
	.b(n25851),
	.c(n25838),
	.d(FE_OFN25876_n25842));
   ao22m01 U18367 (.o(n10403),
	.a(n20972),
	.b(n25922),
	.c(n25908),
	.d(FE_OFN84_n20972));
   ao22m01 U18368 (.o(n10438),
	.a(n20972),
	.b(n25918),
	.c(n25906),
	.d(FE_OFN84_n20972));
   ao22m01 U18369 (.o(n9133),
	.a(n25945),
	.b(n25967),
	.c(n25946),
	.d(FE_OFN25791_n21053));
   ao22m01 U18370 (.o(n9423),
	.a(n21070),
	.b(n25969),
	.c(n25939),
	.d(FE_OFN24767_n21069));
   ao22m01 U18371 (.o(n9458),
	.a(n21070),
	.b(n25964),
	.c(n25936),
	.d(FE_OFN24767_n21069));
   ao22m01 U18372 (.o(n9463),
	.a(n21070),
	.b(n25962),
	.c(n25935),
	.d(FE_OFN24767_n21069));
   ao22m01 U18373 (.o(n9473),
	.a(n21070),
	.b(n25960),
	.c(n25934),
	.d(FE_OFN24767_n21069));
   ao22m01 U18374 (.o(n9488),
	.a(n21070),
	.b(n25958),
	.c(n25933),
	.d(FE_OFN24767_n21069));
   ao22m01 U18375 (.o(n9503),
	.a(n21070),
	.b(n25956),
	.c(n25932),
	.d(FE_OFN24767_n21069));
   oa12m01 U18376 (.o(n9358),
	.a(n22737),
	.b(n22747),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   oa12m01 U18377 (.o(n9363),
	.a(n22738),
	.b(n22739),
	.c(FE_OFN24766_n21069));
   oa12m01 U18378 (.o(n9388),
	.a(n22735),
	.b(n22736),
	.c(FE_OFN25865_FE_OFN24766_n21069));
   oa12m01 U18379 (.o(n9393),
	.a(n22744),
	.b(n22745),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f02 U18380 (.o(n2703),
	.a(n18547),
	.b(n18546));
   no02m01 U18381 (.o(west_input_control_N48),
	.a(FE_OFN25647_reset),
	.b(n25233));
   na02f02 U18382 (.o(n2993),
	.a(n18591),
	.b(n25071));
   no02m01 U18383 (.o(north_output_space_N47),
	.a(n25814),
	.b(north_output_space_N48));
   no02m01 U18384 (.o(south_output_space_N47),
	.a(n25819),
	.b(south_output_space_N48));
   na03m02 U18385 (.o(FE_OFN747_dataOut_W_46),
	.a(n21726),
	.b(n21725),
	.c(n21724));
   na03m02 U18386 (.o(FE_OFN699_dataOut_S_27),
	.a(n22326),
	.b(n22325),
	.c(n22324));
   na03m02 U18387 (.o(dataOut_E_53_),
	.a(n22494),
	.b(n22493),
	.c(n22492));
   na03m02 U18388 (.o(dataOut_P_50_),
	.a(n23347),
	.b(n23346),
	.c(n23345));
   ao12f02 U18389 (.o(n25074),
	.a(n18105),
	.b(n17789),
	.c(thanksIn_P));
   in01f02 U18390 (.o(n23798),
	.a(dataIn_P_24_));
   in01f02 U18391 (.o(n23934),
	.a(dataIn_P_39_));
   in01m03 U18392 (.o(n23924),
	.a(dataIn_P_54_));
   in01f02 U18393 (.o(n23791),
	.a(dataIn_P_31_));
   oa12f04 U18394 (.o(n25277),
	.a(n25275),
	.b(n25432),
	.c(n25276));
   na02f02 U18396 (.o(n18541),
	.a(n18501),
	.b(n18507));
   na02f02 U18397 (.o(n24966),
	.a(n18397),
	.b(n18399));
   no02f04 U18399 (.o(n25186),
	.a(west_output_current_route_connection_0_),
	.b(n25185));
   na02f02 U18400 (.o(n25146),
	.a(n25145),
	.b(n25147));
   oa22s01 U18402 (.o(n25657),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_8_),
	.c(east_input_NIB_storage_data_f_0__8_),
	.d(FE_OFN24862_n22945));
   oa22s01 U18403 (.o(n25658),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_7_),
	.c(east_input_NIB_storage_data_f_0__7_),
	.d(FE_OFN24862_n22945));
   oa22s01 U18404 (.o(n25659),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_6_),
	.c(east_input_NIB_storage_data_f_0__6_),
	.d(FE_OFN24862_n22945));
   oa22s01 U18405 (.o(n25660),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_4_),
	.c(east_input_NIB_storage_data_f_0__4_),
	.d(FE_OFN24862_n22945));
   oa22s01 U18406 (.o(n25661),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_1_),
	.c(east_input_NIB_storage_data_f_0__1_),
	.d(FE_OFN24862_n22945));
   oa22s01 U18407 (.o(n25688),
	.a(FE_OFN24810_n22958),
	.b(dataIn_E_11_),
	.c(east_input_NIB_storage_data_f_2__11_),
	.d(FE_OFN435_n22958));
   oa22s01 U18408 (.o(n25689),
	.a(FE_OFN437_n22958),
	.b(dataIn_E_10_),
	.c(east_input_NIB_storage_data_f_2__10_),
	.d(FE_OFN435_n22958));
   oa22s01 U18409 (.o(n25693),
	.a(FE_OFN24815_n22958),
	.b(dataIn_E_6_),
	.c(east_input_NIB_storage_data_f_2__6_),
	.d(FE_OFN435_n22958));
   oa22s01 U18410 (.o(n25694),
	.a(FE_OFN24810_n22958),
	.b(dataIn_E_4_),
	.c(east_input_NIB_storage_data_f_2__4_),
	.d(FE_OFN435_n22958));
   oa22s01 U18411 (.o(n25695),
	.a(FE_OFN24814_n22958),
	.b(dataIn_E_1_),
	.c(east_input_NIB_storage_data_f_2__1_),
	.d(FE_OFN435_n22958));
   oa12f02 U18412 (.o(n20560),
	.a(n20557),
	.b(FE_RN_12),
	.c(n20558));
   oa22s01 U18413 (.o(n22459),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_17_),
	.c(north_input_NIB_storage_data_f_3__17_),
	.d(n21175));
   oa22s01 U18414 (.o(n22460),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_11_),
	.c(north_input_NIB_storage_data_f_3__11_),
	.d(n21175));
   oa22s01 U18415 (.o(n22450),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_10_),
	.c(north_input_NIB_storage_data_f_3__10_),
	.d(n21175));
   oa22s01 U18416 (.o(n22457),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_9_),
	.c(north_input_NIB_storage_data_f_3__9_),
	.d(n21175));
   oa22s01 U18417 (.o(n22451),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_8_),
	.c(north_input_NIB_storage_data_f_3__8_),
	.d(n21175));
   oa22s01 U18418 (.o(n22456),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_7_),
	.c(north_input_NIB_storage_data_f_3__7_),
	.d(n21175));
   oa22s01 U18419 (.o(n22452),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_5_),
	.c(north_input_NIB_storage_data_f_3__5_),
	.d(n21175));
   oa22s01 U18420 (.o(n22447),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_4_),
	.c(north_input_NIB_storage_data_f_3__4_),
	.d(n21175));
   oa22s01 U18421 (.o(n22446),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_3_),
	.c(north_input_NIB_storage_data_f_3__3_),
	.d(n21175));
   oa22s01 U18422 (.o(n22445),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_2_),
	.c(north_input_NIB_storage_data_f_3__2_),
	.d(n21175));
   oa22s01 U18423 (.o(n22453),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_1_),
	.c(north_input_NIB_storage_data_f_3__1_),
	.d(n21175));
   oa22s01 U18424 (.o(n22449),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_0_),
	.c(north_input_NIB_storage_data_f_3__0_),
	.d(n21175));
   na02s01 U18425 (.o(n25195),
	.a(east_input_NIB_storage_data_f_3__55_),
	.b(FE_OFN943_n24921));
   na02s01 U18426 (.o(n25260),
	.a(east_input_NIB_storage_data_f_3__24_),
	.b(n24921));
   na02s01 U18427 (.o(n25217),
	.a(east_input_NIB_storage_data_f_3__62_),
	.b(FE_OFN943_n24921));
   na02s01 U18428 (.o(n25221),
	.a(east_input_NIB_storage_data_f_3__32_),
	.b(n24921));
   na02s01 U18429 (.o(n25254),
	.a(east_input_NIB_storage_data_f_3__23_),
	.b(n24921));
   na02s01 U18430 (.o(n25258),
	.a(east_input_NIB_storage_data_f_3__29_),
	.b(n24921));
   na02s01 U18431 (.o(n25266),
	.a(east_input_NIB_storage_data_f_3__28_),
	.b(n24921));
   na02s01 U18432 (.o(n25201),
	.a(east_input_NIB_storage_data_f_3__60_),
	.b(FE_OFN943_n24921));
   na02s01 U18433 (.o(n25203),
	.a(east_input_NIB_storage_data_f_3__53_),
	.b(FE_OFN943_n24921));
   na02s01 U18434 (.o(n25205),
	.a(east_input_NIB_storage_data_f_3__57_),
	.b(n24921));
   no03f02 U18435 (.o(n25325),
	.a(n25997),
	.b(n25319),
	.c(n25338));
   na03f08 U18436 (.o(n25137),
	.a(n18286),
	.b(n20142),
	.c(FE_OFN25598_reset));
   na03f01 U18437 (.o(west_output_space_N48),
	.a(n25822),
	.b(n17888),
	.c(n25823));
   na02f06 U18438 (.o(n24988),
	.a(n20346),
	.b(n20122));
   na02s01 U18439 (.o(n22996),
	.a(east_input_NIB_storage_data_f_2__25_),
	.b(n22958));
   na03s01 U18440 (.o(n25495),
	.a(n25494),
	.b(n25493),
	.c(n25492));
   na02s01 U18441 (.o(n22999),
	.a(east_input_NIB_storage_data_f_0__61_),
	.b(FE_OFN432_n22945));
   na02s01 U18442 (.o(n23020),
	.a(east_input_NIB_storage_data_f_0__46_),
	.b(FE_OFN24851_n22945));
   na02s01 U18443 (.o(n23008),
	.a(east_input_NIB_storage_data_f_0__31_),
	.b(FE_OFN24844_n22945));
   na02s01 U18444 (.o(n23022),
	.a(east_input_NIB_storage_data_f_2__55_),
	.b(FE_OFN436_n22958));
   na02s01 U18445 (.o(n22976),
	.a(east_input_NIB_storage_data_f_2__40_),
	.b(n22958));
   na02f02 U18446 (.o(south_output_space_N48),
	.a(n20490),
	.b(n25820));
   oa22m01 U18447 (.o(n22475),
	.a(n25848),
	.b(dataIn_N_20_),
	.c(north_input_NIB_storage_data_f_1__20_),
	.d(n21220));
   oa22m01 U18448 (.o(n22464),
	.a(n25848),
	.b(dataIn_N_10_),
	.c(north_input_NIB_storage_data_f_1__10_),
	.d(n21220));
   oa22m01 U18449 (.o(n22470),
	.a(n25848),
	.b(dataIn_N_9_),
	.c(north_input_NIB_storage_data_f_1__9_),
	.d(n21220));
   oa22m01 U18450 (.o(n22468),
	.a(n25848),
	.b(dataIn_N_4_),
	.c(north_input_NIB_storage_data_f_1__4_),
	.d(n21220));
   oa22m01 U18451 (.o(n22479),
	.a(n25848),
	.b(dataIn_N_3_),
	.c(north_input_NIB_storage_data_f_1__3_),
	.d(n21220));
   oa22m01 U18452 (.o(n22472),
	.a(n25848),
	.b(dataIn_N_2_),
	.c(north_input_NIB_storage_data_f_1__2_),
	.d(n21220));
   oa22m01 U18453 (.o(n22476),
	.a(n25848),
	.b(dataIn_N_1_),
	.c(north_input_NIB_storage_data_f_1__1_),
	.d(n21220));
   oa22m01 U18454 (.o(n22474),
	.a(n25848),
	.b(dataIn_N_0_),
	.c(north_input_NIB_storage_data_f_1__0_),
	.d(n21220));
   na03f02 U18455 (.o(n25477),
	.a(n25974),
	.b(thanksIn_P),
	.c(n25476));
   no03f04 U18456 (.o(n25490),
	.a(thanksIn_P),
	.b(n25482),
	.c(n25481));
   na02f01 U18457 (.o(n21269),
	.a(north_input_NIB_storage_data_f_1__54_),
	.b(n25848));
   na02f01 U18458 (.o(n21228),
	.a(north_input_NIB_storage_data_f_1__39_),
	.b(FE_OFN88_n21220));
   na02s01 U18459 (.o(n21223),
	.a(north_input_NIB_storage_data_f_1__24_),
	.b(FE_OFN88_n21220));
   na02f04 U18460 (.o(n18591),
	.a(n25070),
	.b(FE_RN_3));
   oa22m01 U18461 (.o(n22047),
	.a(FE_OFN25875_n25842),
	.b(dataIn_N_15_),
	.c(north_input_NIB_storage_data_f_2__15_),
	.d(n20656));
   oa22m01 U18462 (.o(n22046),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_14_),
	.c(north_input_NIB_storage_data_f_2__14_),
	.d(n20656));
   oa22m01 U18463 (.o(n22054),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_5_),
	.c(north_input_NIB_storage_data_f_2__5_),
	.d(n20656));
   oa22m01 U18464 (.o(n22050),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_4_),
	.c(north_input_NIB_storage_data_f_2__4_),
	.d(n20656));
   oa22m01 U18465 (.o(n22042),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_3_),
	.c(north_input_NIB_storage_data_f_2__3_),
	.d(n20656));
   oa22m01 U18466 (.o(n22044),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_2_),
	.c(north_input_NIB_storage_data_f_2__2_),
	.d(n20656));
   oa22m01 U18467 (.o(n22055),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_1_),
	.c(north_input_NIB_storage_data_f_2__1_),
	.d(n20656));
   oa22m01 U18468 (.o(n22045),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_0_),
	.c(north_input_NIB_storage_data_f_2__0_),
	.d(n20656));
   na02s01 U18469 (.o(n20686),
	.a(north_input_NIB_storage_data_f_2__59_),
	.b(FE_OFN25876_n25842));
   na02s01 U18470 (.o(n20666),
	.a(north_input_NIB_storage_data_f_2__29_),
	.b(FE_OFN1087_n20656));
   na02s01 U18471 (.o(n22708),
	.a(west_input_NIB_storage_data_f_2__23_),
	.b(n21053));
   na02f01 U18472 (.o(n21122),
	.a(west_input_NIB_storage_data_f_3__31_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U18473 (.o(n21998),
	.a(proc_input_NIB_storage_data_f_14__54_),
	.b(FE_OFN25741_FE_OFN25605_n21944));
   na02f01 U18474 (.o(n21993),
	.a(proc_input_NIB_storage_data_f_14__39_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa22s01 U18475 (.o(n24846),
	.a(n25905),
	.b(dataIn_S_21_),
	.c(south_input_NIB_storage_data_f_2__21_),
	.d(n20972));
   oa22s01 U18476 (.o(n22414),
	.a(n25905),
	.b(dataIn_S_7_),
	.c(south_input_NIB_storage_data_f_2__7_),
	.d(n20972));
   oa22s01 U18477 (.o(n22393),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_6_),
	.c(south_input_NIB_storage_data_f_2__6_),
	.d(n20972));
   oa22s01 U18478 (.o(n22409),
	.a(n25905),
	.b(dataIn_S_5_),
	.c(south_input_NIB_storage_data_f_2__5_),
	.d(n20972));
   oa22s01 U18479 (.o(n22408),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_4_),
	.c(south_input_NIB_storage_data_f_2__4_),
	.d(n20972));
   oa22s01 U18480 (.o(n22413),
	.a(n25905),
	.b(dataIn_S_3_),
	.c(south_input_NIB_storage_data_f_2__3_),
	.d(n20972));
   oa22s01 U18481 (.o(n22397),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_2_),
	.c(south_input_NIB_storage_data_f_2__2_),
	.d(n20972));
   oa22s01 U18482 (.o(n22410),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_1_),
	.c(south_input_NIB_storage_data_f_2__1_),
	.d(n20972));
   oa22s01 U18483 (.o(n22406),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_0_),
	.c(south_input_NIB_storage_data_f_2__0_),
	.d(n20972));
   oa22m01 U18484 (.o(n24851),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_20_),
	.c(west_input_NIB_storage_data_f_2__20_),
	.d(n25945));
   oa22m01 U18485 (.o(n22423),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_5_),
	.c(west_input_NIB_storage_data_f_2__5_),
	.d(n25945));
   oa22m01 U18486 (.o(n22421),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_0_),
	.c(west_input_NIB_storage_data_f_2__0_),
	.d(n25945));
   oa22m01 U18487 (.o(n23477),
	.a(FE_OFN101_n22098),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_9__14_),
	.d(n22098));
   oa22m01 U18488 (.o(n23475),
	.a(FE_OFN101_n22098),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_9__13_),
	.d(n22098));
   oa22m01 U18489 (.o(n23428),
	.a(FE_OFN101_n22098),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_9__6_),
	.d(n22098));
   oa22m01 U18490 (.o(n23423),
	.a(FE_OFN101_n22098),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_9__5_),
	.d(n22098));
   oa22m01 U18491 (.o(n23421),
	.a(FE_OFN465_n23476),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_9__4_),
	.d(n22098));
   oa22m01 U18492 (.o(n23420),
	.a(FE_OFN465_n23476),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_9__3_),
	.d(n22098));
   oa22m01 U18493 (.o(n23435),
	.a(FE_OFN101_n22098),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_9__2_),
	.d(n22098));
   oa22m01 U18494 (.o(n23418),
	.a(FE_OFN465_n23476),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_9__1_),
	.d(n22098));
   oa22m01 U18495 (.o(n23417),
	.a(FE_OFN465_n23476),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_9__0_),
	.d(n22098));
   oa22m01 U18496 (.o(n23457),
	.a(n23471),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_8__9_),
	.d(FE_OFN416_n22085));
   oa22m01 U18497 (.o(n23456),
	.a(n23471),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_8__8_),
	.d(FE_OFN416_n22085));
   oa22m01 U18498 (.o(n23452),
	.a(n23471),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_8__6_),
	.d(FE_OFN416_n22085));
   oa22m01 U18499 (.o(n23468),
	.a(n22085),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_8__5_),
	.d(FE_OFN416_n22085));
   oa22m01 U18500 (.o(n23450),
	.a(n23471),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_8__4_),
	.d(FE_OFN416_n22085));
   oa22m01 U18501 (.o(n23449),
	.a(n23471),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_8__3_),
	.d(FE_OFN416_n22085));
   oa22m01 U18502 (.o(n23448),
	.a(n23471),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_8__2_),
	.d(FE_OFN416_n22085));
   oa22m01 U18503 (.o(n23447),
	.a(n23471),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_8__1_),
	.d(FE_OFN416_n22085));
   oa22m01 U18504 (.o(n23446),
	.a(n23471),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_8__0_),
	.d(FE_OFN416_n22085));
   oa22m01 U18505 (.o(n23427),
	.a(n23453),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_10__19_),
	.d(n22140));
   oa22m01 U18506 (.o(n23426),
	.a(FE_OFN103_n22140),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_10__18_),
	.d(FE_OFN104_n22140));
   oa22m01 U18507 (.o(n23451),
	.a(n23453),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_10__6_),
	.d(n22140));
   oa22m01 U18508 (.o(n23434),
	.a(n23453),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_10__5_),
	.d(n22140));
   oa22m01 U18509 (.o(n23430),
	.a(FE_OFN103_n22140),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_10__4_),
	.d(FE_OFN104_n22140));
   oa22m01 U18510 (.o(n23415),
	.a(n23453),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_10__3_),
	.d(n22140));
   oa22m01 U18511 (.o(n23422),
	.a(n23453),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_10__2_),
	.d(n22140));
   oa22m01 U18512 (.o(n23424),
	.a(FE_OFN103_n22140),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_10__1_),
	.d(FE_OFN104_n22140));
   oa22m01 U18513 (.o(n23425),
	.a(n23453),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_10__0_),
	.d(n22140));
   oa22m01 U18514 (.o(n23254),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_14__9_),
	.d(n21945));
   oa22m01 U18515 (.o(n23252),
	.a(FE_OFN25605_n21944),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_14__11_),
	.d(n23262));
   oa22m01 U18516 (.o(n23253),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_14__10_),
	.d(n21945));
   oa22m01 U18517 (.o(n23257),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_14__6_),
	.d(n21945));
   oa22m01 U18518 (.o(n23258),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_14__5_),
	.d(n21945));
   oa22m01 U18519 (.o(n23259),
	.a(FE_OFN25605_n21944),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_14__4_),
	.d(n23262));
   oa22m01 U18520 (.o(n23260),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_14__3_),
	.d(n21945));
   oa22m01 U18521 (.o(n23261),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_14__2_),
	.d(n21945));
   oa22m01 U18522 (.o(n23263),
	.a(FE_OFN25605_n21944),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_14__1_),
	.d(n23262));
   oa22m01 U18523 (.o(n23248),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_14__0_),
	.d(n21945));
   oa22m01 U18524 (.o(n23193),
	.a(FE_OFN25626_n21910),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_12__14_),
	.d(n23246));
   oa22m01 U18525 (.o(n23205),
	.a(FE_OFN25628_n21910),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_12__16_),
	.d(FE_OFN912_n23246));
   oa22m01 U18526 (.o(n23204),
	.a(FE_OFN25626_n21910),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_12__15_),
	.d(FE_OFN912_n23246));
   oa22m01 U18527 (.o(n23211),
	.a(FE_OFN25629_n21910),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_12__6_),
	.d(FE_OFN912_n23246));
   oa22m01 U18528 (.o(n23198),
	.a(FE_OFN25626_n21910),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_12__5_),
	.d(FE_OFN912_n23246));
   oa22m01 U18529 (.o(n23202),
	.a(FE_OFN25629_n21910),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_12__4_),
	.d(FE_OFN912_n23246));
   oa22m01 U18530 (.o(n23201),
	.a(FE_OFN25628_n21910),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_12__3_),
	.d(FE_OFN912_n23246));
   oa22m01 U18531 (.o(n23210),
	.a(FE_OFN25629_n21910),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_12__2_),
	.d(FE_OFN912_n23246));
   oa22m01 U18532 (.o(n23220),
	.a(FE_OFN25628_n21910),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_12__1_),
	.d(FE_OFN912_n23246));
   oa22m01 U18533 (.o(n23221),
	.a(FE_OFN25629_n21910),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_12__0_),
	.d(FE_OFN912_n23246));
   oa22m01 U18534 (.o(n23206),
	.a(FE_OFN448_n23236),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_13__33_),
	.d(n21915));
   oa22m01 U18535 (.o(n23225),
	.a(n23236),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_13__19_),
	.d(n21915));
   oa22m01 U18536 (.o(n23207),
	.a(FE_OFN448_n23236),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_13__21_),
	.d(n21915));
   oa22m01 U18537 (.o(n23208),
	.a(FE_OFN448_n23236),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_13__20_),
	.d(n21915));
   oa22m01 U18538 (.o(n23229),
	.a(n23236),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_13__6_),
	.d(n21915));
   oa22m01 U18539 (.o(n23230),
	.a(n23236),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_13__5_),
	.d(n21915));
   oa22m01 U18540 (.o(n23232),
	.a(n23236),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_13__4_),
	.d(n21915));
   oa22m01 U18541 (.o(n23233),
	.a(FE_OFN25781_FE_OFN448_n23236),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_13__3_),
	.d(n21915));
   oa22m01 U18542 (.o(n23234),
	.a(n23236),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_13__2_),
	.d(n21915));
   oa22m01 U18543 (.o(n23235),
	.a(FE_OFN448_n23236),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_13__1_),
	.d(n21915));
   oa22m01 U18544 (.o(n23237),
	.a(n23236),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_13__0_),
	.d(n21915));
   oa22s01 U18545 (.o(n24860),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_21_),
	.c(west_input_NIB_storage_data_f_3__21_),
	.d(n21070));
   oa22s01 U18546 (.o(n22417),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_8_),
	.c(west_input_NIB_storage_data_f_3__8_),
	.d(n21070));
   oa22s01 U18547 (.o(n24850),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_13_),
	.c(west_input_NIB_storage_data_f_3__13_),
	.d(n21070));
   oa22s01 U18548 (.o(n22419),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_3_),
	.c(west_input_NIB_storage_data_f_3__3_),
	.d(n21070));
   oa22s01 U18549 (.o(n22425),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_0_),
	.c(west_input_NIB_storage_data_f_3__0_),
	.d(n21070));
   na02s01 U18550 (.o(n21177),
	.a(north_input_NIB_storage_data_f_3__56_),
	.b(FE_OFN86_n21175));
   na02f04 U18551 (.o(n25060),
	.a(n25059),
	.b(n25058));
   na02s01 U18552 (.o(n22094),
	.a(proc_input_NIB_storage_data_f_8__52_),
	.b(n23471));
   na02s01 U18553 (.o(n22184),
	.a(proc_input_NIB_storage_data_f_10__62_),
	.b(n23453));
   na02s01 U18554 (.o(n22167),
	.a(proc_input_NIB_storage_data_f_10__47_),
	.b(FE_OFN103_n22140));
   na02s01 U18555 (.o(n20993),
	.a(south_input_NIB_storage_data_f_2__27_),
	.b(FE_OFN84_n20972));
   na02s01 U18556 (.o(n20674),
	.a(north_input_NIB_storage_data_f_2__44_),
	.b(FE_OFN1087_n20656));
   na02s01 U18557 (.o(n21978),
	.a(proc_input_NIB_storage_data_f_14__24_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   na02s01 U18558 (.o(n22113),
	.a(proc_input_NIB_storage_data_f_8__37_),
	.b(n22085));
   na02s01 U18559 (.o(n22128),
	.a(proc_input_NIB_storage_data_f_8__22_),
	.b(n22085));
   na02s01 U18560 (.o(n22151),
	.a(proc_input_NIB_storage_data_f_10__32_),
	.b(FE_OFN103_n22140));
   na02s01 U18561 (.o(n21964),
	.a(proc_input_NIB_storage_data_f_12__59_),
	.b(FE_OFN25628_n21910));
   na02f01 U18562 (.o(n21933),
	.a(proc_input_NIB_storage_data_f_12__44_),
	.b(FE_OFN25627_n21910));
   na02f01 U18563 (.o(n21959),
	.a(proc_input_NIB_storage_data_f_12__29_),
	.b(FE_OFN25626_n21910));
   na02s01 U18564 (.o(n21930),
	.a(proc_input_NIB_storage_data_f_13__49_),
	.b(n23236));
   na02f01 U18565 (.o(n22016),
	.a(proc_input_NIB_storage_data_f_13__34_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   na02s01 U18566 (.o(n22135),
	.a(proc_input_NIB_storage_data_f_9__57_),
	.b(FE_OFN465_n23476));
   na02s01 U18567 (.o(n22200),
	.a(proc_input_NIB_storage_data_f_9__42_),
	.b(FE_OFN101_n22098));
   na02s01 U18568 (.o(n22214),
	.a(proc_input_NIB_storage_data_f_9__27_),
	.b(FE_OFN465_n23476));
   in01f04 U18569 (.o(n24728),
	.a(n25301));
   ao12m01 U18570 (.o(n25794),
	.a(n25792),
	.b(ec_thanks_w_to_e_reg),
	.c(n25793));
   ao22s01 U18571 (.o(n25771),
	.a(ec_thanks_w_to_s_reg),
	.b(n25770),
	.c(ec_cfg_8_),
	.d(n25769));
   in01f01 U18572 (.o(n18103),
	.a(n19646));
   no02f04 U18573 (.o(n23585),
	.a(n21778),
	.b(n21777));
   in01f02 U18574 (.o(n20142),
	.a(n25083));
   no02f06 U18575 (.o(n25111),
	.a(thanksIn_P),
	.b(n25971));
   in01f04 U18576 (.o(n25881),
	.a(n24761));
   no02f04 U18579 (.o(n18604),
	.a(n18605),
	.b(n18399));
   in01f01 U18580 (.o(n20345),
	.a(n18057));
   no04f02 U18581 (.o(n25330),
	.a(FE_OFN25601_reset),
	.b(n25984),
	.c(n25985),
	.d(n25327));
   no03f02 U18582 (.o(n25391),
	.a(reset),
	.b(n25386),
	.c(FE_OFN565_n25385));
   no02f04 U18583 (.o(n25993),
	.a(FE_OFN25600_reset),
	.b(n18575));
   na02f04 U18584 (.o(n25099),
	.a(n25098),
	.b(n18274));
   na02f03 U18585 (.o(n20537),
	.a(n25177),
	.b(n25180));
   no02m02 U18586 (.o(n20557),
	.a(reset),
	.b(n20556));
   no04m01 U18587 (.o(n25290),
	.a(north_input_NIB_elements_in_array_f_2_),
	.b(n25289),
	.c(n25288),
	.d(n25287));
   no03s01 U18588 (.o(n22915),
	.a(south_input_control_count_f_7_),
	.b(n23553),
	.c(n25250));
   in01f02 U18589 (.o(n20346),
	.a(n20338));
   no02f04 U18590 (.o(n25485),
	.a(thanksIn_P),
	.b(n25481));
   in01f08 U18591 (.o(n26013),
	.a(n18540));
   ao12f04 U18592 (.o(n24960),
	.a(FE_OFN4_reset),
	.b(n24953),
	.c(n18570));
   no02f08 U18593 (.o(n25105),
	.a(n25083),
	.b(n25082));
   no04f03 U18594 (.o(n25037),
	.a(FE_OFN5_reset),
	.b(n25036),
	.c(n25035),
	.d(n25309));
   no02f01 U18595 (.o(n25399),
	.a(reset),
	.b(n25394));
   ao22f01 U18596 (.o(n21896),
	.a(n20723),
	.b(north_input_control_count_f_6_),
	.c(n20722),
	.d(n20705));
   na03f01 U18597 (.o(n25823),
	.a(n25452),
	.b(n25451),
	.c(n25450));
   na03f01 U18598 (.o(n25816),
	.a(n25366),
	.b(n25365),
	.c(n25364));
   in01f01 U18599 (.o(n18096),
	.a(n22842));
   na04f04 U18600 (.o(n21777),
	.a(n21776),
	.b(n21775),
	.c(n21774),
	.d(n21773));
   na04f04 U18601 (.o(n21778),
	.a(n21772),
	.b(n21771),
	.c(n21770),
	.d(n21769));
   na04f02 U18602 (.o(n24356),
	.a(n24348),
	.b(n24347),
	.c(n24346),
	.d(n24345));
   na04f04 U18603 (.o(n24355),
	.a(n24354),
	.b(n24353),
	.c(n24352),
	.d(n24351));
   na04f04 U18604 (.o(n24094),
	.a(n24087),
	.b(n24086),
	.c(n24085),
	.d(n24084));
   na04f02 U18605 (.o(n24138),
	.a(n24137),
	.b(n24136),
	.c(n24135),
	.d(n24134));
   na04f04 U18606 (.o(n24047),
	.a(n24041),
	.b(n24040),
	.c(n24039),
	.d(n24038));
   na04f02 U18607 (.o(n24071),
	.a(n24064),
	.b(n24063),
	.c(n24062),
	.d(n24061));
   na04f04 U18608 (.o(n21308),
	.a(n21302),
	.b(n21301),
	.c(n21300),
	.d(n21299));
   na04f02 U18609 (.o(n21307),
	.a(n21306),
	.b(n21305),
	.c(n21304),
	.d(n21303));
   na04f03 U18610 (.o(n21358),
	.a(n21352),
	.b(n21351),
	.c(n21350),
	.d(n21349));
   na04f03 U18611 (.o(n21824),
	.a(n21818),
	.b(n21817),
	.c(n21816),
	.d(n21815));
   na04f03 U18612 (.o(n21823),
	.a(n21822),
	.b(n21821),
	.c(n21820),
	.d(n21819));
   na04f03 U18613 (.o(n21754),
	.a(n21753),
	.b(n21752),
	.c(n21751),
	.d(n21750));
   na04f04 U18615 (.o(n24298),
	.a(n24292),
	.b(n24291),
	.c(n24290),
	.d(n24289));
   na04f04 U18616 (.o(n24297),
	.a(n24296),
	.b(n24295),
	.c(n24294),
	.d(n24293));
   na04f02 U18617 (.o(n24275),
	.a(n24274),
	.b(n24273),
	.c(n24272),
	.d(n24271));
   na04f04 U18618 (.o(n24253),
	.a(n24252),
	.b(n24251),
	.c(n24250),
	.d(n24249));
   na04f03 U18619 (.o(n24231),
	.a(n24225),
	.b(n24224),
	.c(n24223),
	.d(n24222));
   na04f02 U18620 (.o(n24207),
	.a(n24201),
	.b(n24200),
	.c(n24199),
	.d(n24198));
   na04f02 U18621 (.o(n21856),
	.a(n21850),
	.b(n21849),
	.c(n21848),
	.d(n21847));
   na04f02 U18623 (.o(n21357),
	.a(n21356),
	.b(n21355),
	.c(n21354),
	.d(n21353));
   na04f04 U18624 (.o(n24139),
	.a(n24133),
	.b(n24132),
	.c(n24131),
	.d(n24130));
   na04f03 U18625 (.o(n24046),
	.a(n24045),
	.b(n24044),
	.c(n24043),
	.d(n24042));
   na04f03 U18626 (.o(n21755),
	.a(n21744),
	.b(n21743),
	.c(n21742),
	.d(n21741));
   na04f03 U18627 (.o(n24161),
	.a(n24160),
	.b(n24159),
	.c(n24158),
	.d(n24157));
   na04f04 U18628 (.o(n21800),
	.a(n21799),
	.b(n21798),
	.c(n21797),
	.d(n21796));
   na04f03 U18629 (.o(n24254),
	.a(n24248),
	.b(n24247),
	.c(n24246),
	.d(n24245));
   na04f02 U18631 (.o(n24461),
	.a(n24452),
	.b(n24451),
	.c(n24450),
	.d(n24449));
   na04f04 U18632 (.o(n24162),
	.a(n24156),
	.b(n24155),
	.c(n24154),
	.d(n24153));
   na04f03 U18633 (.o(n24388),
	.a(n24387),
	.b(n24386),
	.c(n24385),
	.d(n24384));
   na04f02 U18634 (.o(n24184),
	.a(n24183),
	.b(n24182),
	.c(n24181),
	.d(n24180));
   na04f03 U18635 (.o(n24185),
	.a(n24179),
	.b(n24178),
	.c(n24177),
	.d(n24176));
   na04f04 U18636 (.o(n24320),
	.a(n24314),
	.b(n24313),
	.c(n24312),
	.d(n24311));
   na04f02 U18637 (.o(n21855),
	.a(n21854),
	.b(n21853),
	.c(n21852),
	.d(n21851));
   na04f04 U18638 (.o(n24115),
	.a(n24114),
	.b(n24113),
	.c(n24112),
	.d(n24111));
   na04f02 U18639 (.o(n24319),
	.a(n24318),
	.b(n24317),
	.c(n24316),
	.d(n24315));
   na04f04 U18640 (.o(n24070),
	.a(n24069),
	.b(n24068),
	.c(n24067),
	.d(n24066));
   na04f02 U18641 (.o(n24460),
	.a(n24459),
	.b(n24458),
	.c(n24457),
	.d(n24456));
   na04f02 U18642 (.o(n24116),
	.a(n24110),
	.b(n24109),
	.c(n24108),
	.d(n24107));
   na04f03 U18643 (.o(n24276),
	.a(n24270),
	.b(n24269),
	.c(n24268),
	.d(n24267));
   na04f04 U18644 (.o(n24389),
	.a(n24383),
	.b(n24382),
	.c(n24381),
	.d(n24380));
   na04f03 U18645 (.o(n24206),
	.a(n24205),
	.b(n24204),
	.c(n24203),
	.d(n24202));
   no02f08 U18646 (.o(n25184),
	.a(n20541),
	.b(n20530));
   in01f01 U18647 (.o(n25134),
	.a(n25091));
   na02f02 U18648 (.o(n24980),
	.a(n17749),
	.b(n24978));
   in01f04 U18653 (.o(n25395),
	.a(FE_OFN269_n25506));
   na03f10 U18656 (.o(n25384),
	.a(n20553),
	.b(n20326),
	.c(n20551));
   in01f03 U18657 (.o(n20539),
	.a(n20530));
   no04f04 U18658 (.o(n25336),
	.a(n25984),
	.b(n25997),
	.c(n25334),
	.d(n25333));
   na03f06 U18661 (.o(n20532),
	.a(n25170),
	.b(n20531),
	.c(FE_OFN393_n19446));
   na02f10 U18662 (.o(n18057),
	.a(n18012),
	.b(n17749));
   na03f08 U18663 (.o(n20338),
	.a(n20120),
	.b(n18625),
	.c(n18571));
   no03f04 U18664 (.o(n20315),
	.a(n20266),
	.b(n19020),
	.c(n20312));
   na02f06 U18665 (.o(n24990),
	.a(FE_OFN25599_reset),
	.b(n24958));
   na02f08 U18666 (.o(n18540),
	.a(FE_OFN25597_reset),
	.b(n18507));
   no02f02 U18668 (.o(n25394),
	.a(n25393),
	.b(n25392));
   in01s01 U18669 (.o(n25482),
	.a(proc_input_NIB_elements_in_array_f_3_));
   in01f02 U18670 (.o(n18191),
	.a(n18192));
   in01f08 U18671 (.o(n25142),
	.a(thanksIn_P));
   no03f06 U18672 (.o(n18500),
	.a(n25406),
	.b(n25404),
	.c(n25405));
   ao22m02 U18673 (.o(n25305),
	.a(proc_output_control_planned_f),
	.b(n25300),
	.c(n25414),
	.d(n25299));
   in01f04 U18674 (.o(n25178),
	.a(n25177));
   na03f02 U18675 (.o(n18281),
	.a(n25091),
	.b(n25128),
	.c(n19054));
   no02f04 U18677 (.o(n20121),
	.a(south_output_control_planned_f),
	.b(validOut_S));
   in01s01 U18678 (.o(n18083),
	.a(proc_input_NIB_elements_in_array_f_1_));
   na03s01 U18681 (.o(n18398),
	.a(FE_OFN24745_n18648),
	.b(n24965),
	.c(FE_OFN575_n25463));
   no02f04 U18682 (.o(n25311),
	.a(n25036),
	.b(n25031));
   na02s01 U18683 (.o(n18574),
	.a(n20506),
	.b(n20507));
   no02f03 U18684 (.o(n25496),
	.a(west_output_control_planned_f),
	.b(n20534));
   no02m01 U18685 (.o(n25063),
	.a(east_output_current_route_connection_1_),
	.b(n25062));
   na03s01 U18686 (.o(n18506),
	.a(FE_OFN30_n18974),
	.b(n24465),
	.c(FE_OFN573_n25463));
   na02s01 U18687 (.o(n18257),
	.a(n23316),
	.b(n19017));
   na02s01 U18688 (.o(n18260),
	.a(n23316),
	.b(FE_OFN44_n19054));
   na02s01 U18689 (.o(n18269),
	.a(n18670),
	.b(n17787));
   no03f06 U18690 (.o(n25036),
	.a(n25028),
	.b(n17759),
	.c(n25027));
   na02f02 U18691 (.o(n21174),
	.a(n21218),
	.b(n21173));
   in01f04 U18692 (.o(n25169),
	.a(n20534));
   ao22f04 U18693 (.o(n20553),
	.a(n26025),
	.b(n25078),
	.c(n20322),
	.d(n20321));
   in01f08 U18694 (.o(n17858),
	.a(n17859));
   in01f08 U18695 (.o(n17860),
	.a(n20332));
   in01f06 U18696 (.o(n18571),
	.a(n18465));
   no02f06 U18697 (.o(n25180),
	.a(n20413),
	.b(n20412));
   in01f02 U18698 (.o(n18428),
	.a(n25170));
   na03f08 U18699 (.o(n24958),
	.a(n17792),
	.b(n18625),
	.c(n18167));
   in01f02 U18700 (.o(n24959),
	.a(n24973));
   no03f04 U18701 (.o(n25031),
	.a(n25030),
	.b(n17759),
	.c(n25029));
   no02f10 U18702 (.o(n25177),
	.a(n18432),
	.b(n18431));
   ao22f04 U18703 (.o(n25081),
	.a(n25077),
	.b(n25985),
	.c(n26023),
	.d(n25078));
   na03f03 U18704 (.o(n20550),
	.a(n25062),
	.b(n25387),
	.c(n20549));
   na02f06 U18706 (.o(n20551),
	.a(n26011),
	.b(n22216));
   no02f08 U18707 (.o(n20535),
	.a(n20426),
	.b(n22912));
   oa12f08 U18708 (.o(n18287),
	.a(n20141),
	.b(north_output_control_planned_f),
	.c(validOut_N));
   in01f02 U18709 (.o(n25862),
	.a(n24920));
   no02f04 U18710 (.o(validOut_S),
	.a(n18443),
	.b(n19955));
   no02f01 U18711 (.o(n22944),
	.a(east_input_NIB_tail_ptr_f_1_),
	.b(n25316));
   na02f02 U18712 (.o(n25250),
	.a(south_input_control_thanks_all_f),
	.b(n22912));
   na02f06 U18713 (.o(n25085),
	.a(n25128),
	.b(n25132));
   ao22f01 U18714 (.o(n25237),
	.a(south_input_control_count_f_6_),
	.b(n23553),
	.c(n23552),
	.d(n23551));
   in01m04 U18715 (.o(n17888),
	.a(FE_OFN5_reset));
   in01f01 U18716 (.o(n18194),
	.a(n25329));
   na02f02 U18717 (.o(n21069),
	.a(n21068),
	.b(west_input_NIB_tail_ptr_f_0_));
   na02f02 U18718 (.o(n18192),
	.a(n18199),
	.b(n18601));
   na02f02 U18719 (.o(n20814),
	.a(n18644),
	.b(n20813));
   na02f02 U18720 (.o(n23101),
	.a(n23100),
	.b(n23760));
   na02f02 U18721 (.o(n23789),
	.a(n25976),
	.b(n23788));
   no02f08 U18722 (.o(n25302),
	.a(n25406),
	.b(n25404));
   in01f01 U18723 (.o(n25317),
	.a(n25985));
   na02f02 U18724 (.o(n25080),
	.a(n26021),
	.b(n25079));
   no02f06 U18725 (.o(n25389),
	.a(n18206),
	.b(n18200));
   no02f08 U18726 (.o(n20541),
	.a(west_output_control_planned_f),
	.b(validOut_W));
   na02f04 U18727 (.o(n22778),
	.a(n22777),
	.b(n25980));
   na03m02 U18728 (.o(n20469),
	.a(north_output_current_route_connection_2_),
	.b(FE_OFN255_n25247),
	.c(n20471));
   no03f04 U18729 (.o(n25035),
	.a(proc_output_control_planned_f),
	.b(n25024),
	.c(n25023));
   na02f02 U18730 (.o(n20854),
	.a(n18632),
	.b(n20853));
   na02f02 U18731 (.o(n22084),
	.a(n22777),
	.b(n25976));
   na02f02 U18732 (.o(n22097),
	.a(n22777),
	.b(n22096));
   na02f02 U18733 (.o(n22139),
	.a(n22777),
	.b(n22138));
   na02f03 U18734 (.o(n22273),
	.a(n22272),
	.b(n22271));
   na02f03 U18735 (.o(n23050),
	.a(n23100),
	.b(n23736));
   na02f03 U18736 (.o(n21052),
	.a(n21068),
	.b(n25928));
   ao12s01 U18737 (.o(n21685),
	.a(n21684),
	.b(n21686),
	.c(n21687));
   na02f03 U18738 (.o(n20858),
	.a(n18632),
	.b(n20857));
   na02f04 U18739 (.o(n20796),
	.a(n18644),
	.b(n20795));
   na02f01 U18740 (.o(n21219),
	.a(n21218),
	.b(n21217));
   in01f08 U18743 (.o(n17787),
	.a(n25029));
   in01f08 U18744 (.o(n17786),
	.a(FE_OFN110_n22771));
   in01f08 U18745 (.o(n17755),
	.a(n22772));
   in01f02 U18746 (.o(n20321),
	.a(n23400));
   in01f08 U18747 (.o(n18220),
	.a(n18527));
   in01f06 U18748 (.o(n25032),
	.a(n26028));
   in01f06 U18749 (.o(n18207),
	.a(n18208));
   no03f10 U18750 (.o(n20548),
	.a(n23400),
	.b(n25030),
	.c(n20323));
   no02f02 U18751 (.o(n25976),
	.a(proc_input_NIB_tail_ptr_f_1_),
	.b(proc_input_NIB_tail_ptr_f_0_));
   no03f04 U18752 (.o(n20413),
	.a(n20407),
	.b(n20406),
	.c(n20737));
   ao22f08 U18753 (.o(n20360),
	.a(n26019),
	.b(n25078),
	.c(n20519),
	.d(n25077));
   in01m02 U18754 (.o(n20476),
	.a(n25132));
   na02f08 U18755 (.o(n18217),
	.a(n26022),
	.b(n22216));
   no02m02 U18756 (.o(n25408),
	.a(n25007),
	.b(n24994));
   no02f04 U18757 (.o(n22777),
	.a(proc_input_NIB_tail_ptr_f_2_),
	.b(n22270));
   no02f06 U18758 (.o(n18167),
	.a(n18443),
	.b(n18168));
   no02f02 U18760 (.o(n25227),
	.a(west_input_control_count_f_5_),
	.b(n21379));
   no02f01 U18761 (.o(n18601),
	.a(east_input_NIB_elements_in_array_f_1_),
	.b(n25315));
   no02f08 U18762 (.o(validOut_W),
	.a(n20529),
	.b(n20528));
   na02f08 U18765 (.o(n25091),
	.a(FE_OFN255_n25247),
	.b(n20471));
   no02m01 U18767 (.o(n20853),
	.a(west_input_NIB_tail_ptr_f_0_),
	.b(west_input_NIB_tail_ptr_f_1_));
   na02f06 U18768 (.o(n20477),
	.a(FE_OFN428_n22902),
	.b(n25132));
   in01f01 U18769 (.o(n18112),
	.a(n22216));
   no02s02 U18770 (.o(n25370),
	.a(north_output_space_yummy_f),
	.b(n22936));
   no02f02 U18771 (.o(n21943),
	.a(n23733),
	.b(n22270));
   no02f02 U18772 (.o(n25826),
	.a(north_input_NIB_tail_ptr_f_0_),
	.b(n25287));
   ao22f01 U18773 (.o(n24260),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__14_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__14_));
   na02f01 U18774 (.o(n25726),
	.a(ec_cfg_1_),
	.b(n25725));
   no02f10 U18775 (.o(n26011),
	.a(n23400),
	.b(n20214));
   no02f08 U18778 (.o(n18443),
	.a(south_output_control_planned_f),
	.b(n24968));
   no03f08 U18779 (.o(n25062),
	.a(n20311),
	.b(n20310),
	.c(n20309));
   in01f08 U18780 (.o(n21666),
	.a(n25521));
   na02f06 U18781 (.o(n18080),
	.a(n18138),
	.b(n18139));
   na02f02 U18782 (.o(n22270),
	.a(n25979),
	.b(proc_input_NIB_tail_ptr_f_3_));
   na03f08 U18783 (.o(n20471),
	.a(n25115),
	.b(n18353),
	.c(n25114));
   in01f02 U18784 (.o(n24999),
	.a(n25405));
   no02f02 U18785 (.o(n17866),
	.a(n18377),
	.b(FE_OFN946_n25096));
   no02f02 U18786 (.o(n20289),
	.a(n20271),
	.b(n20270));
   no02f20 U18787 (.o(n26028),
	.a(n17759),
	.b(n25411));
   in01f08 U18788 (.o(n25294),
	.a(n25411));
   no02f08 U18789 (.o(n20428),
	.a(n20520),
	.b(n20427));
   in01f02 U18790 (.o(n25030),
	.a(n20352));
   no02f08 U18791 (.o(n25984),
	.a(n23400),
	.b(n20517));
   no02f04 U18792 (.o(n25999),
	.a(n20504),
	.b(n20331));
   in01f06 U18793 (.o(n17794),
	.a(n20115));
   ao12f02 U18794 (.o(n20358),
	.a(n20350),
	.b(n20351),
	.c(n20514));
   no02f02 U18795 (.o(n20522),
	.a(n20518),
	.b(n25985));
   no02f02 U18796 (.o(n24978),
	.a(n20337),
	.b(n22902));
   no02f10 U18797 (.o(n26006),
	.a(n19070),
	.b(n25025));
   na02f06 U18798 (.o(n25287),
	.a(validIn_N),
	.b(FE_OFN25596_reset));
   na02f02 U18799 (.o(n20489),
	.a(n20496),
	.b(south_output_space_count_f_1_));
   na02f01 U18800 (.o(n20287),
	.a(n20286),
	.b(n20285));
   no02f08 U18801 (.o(n25997),
	.a(n20504),
	.b(n20503));
   in01f06 U18802 (.o(n19743),
	.a(n20222));
   na03f02 U18803 (.o(n20472),
	.a(n24998),
	.b(n23482),
	.c(n25405));
   in01f08 U18804 (.o(n17760),
	.a(n25000));
   in01f02 U18805 (.o(n20165),
	.a(n20407));
   oa22f08 U18806 (.o(n20334),
	.a(n17827),
	.b(n20208),
	.c(n19567),
	.d(n19568));
   in01f02 U18807 (.o(n20212),
	.a(n20213));
   na02f01 U18808 (.o(n20135),
	.a(north_output_current_route_connection_2_),
	.b(n20138));
   in01f02 U18809 (.o(n18466),
	.a(n20223));
   no03f04 U18810 (.o(n20309),
	.a(n20308),
	.b(n20403),
	.c(n20737));
   na02f08 U18811 (.o(n20118),
	.a(n25077),
	.b(n19954));
   oa12f03 U18812 (.o(n25025),
	.a(n19068),
	.b(n19069),
	.c(n25020));
   no02f08 U18813 (.o(n20520),
	.a(FE_OFN25676_n20422),
	.b(n20351));
   na02f03 U18814 (.o(n25115),
	.a(n20465),
	.b(n25018));
   no02f02 U18815 (.o(n18556),
	.a(n20381),
	.b(n18557));
   ao12f08 U18816 (.o(n17936),
	.a(n24970),
	.b(n17829),
	.c(n17828));
   in01f01 U18817 (.o(n20264),
	.a(n20448));
   in01f01 U18818 (.o(n20371),
	.a(n20369));
   no02s02 U18819 (.o(n20727),
	.a(west_input_control_count_f_3_),
	.b(n20633));
   in01f01 U18821 (.o(n25010),
	.a(n23035));
   no02f04 U18825 (.o(n23734),
	.a(proc_input_NIB_tail_ptr_f_3_),
	.b(n25971));
   na03m02 U18826 (.o(n22082),
	.a(proc_output_space_count_f_0_),
	.b(proc_output_space_yummy_f),
	.c(n22061));
   in01s01 U18827 (.o(n21151),
	.a(east_input_control_thanks_all_f));
   na03m02 U18828 (.o(n22392),
	.a(east_output_space_count_f_0_),
	.b(east_output_space_yummy_f),
	.c(n22371));
   in01f02 U18829 (.o(n18353),
	.a(n18354));
   na02s06 U18830 (.o(n20137),
	.a(n25521),
	.b(n20138));
   na02f02 U18831 (.o(n20139),
	.a(n19057),
	.b(n20138));
   oa12f02 U18832 (.o(n20111),
	.a(n20108),
	.b(FE_RN_9),
	.c(n20109));
   no03f03 U18833 (.o(n20310),
	.a(n20297),
	.b(n20296),
	.c(n20295));
   na02f08 U18834 (.o(n18642),
	.a(FE_OFN259_n25295),
	.b(validOut_P));
   no02f03 U18835 (.o(n20355),
	.a(n20353),
	.b(n20352));
   na02f01 U18836 (.o(n19471),
	.a(FE_OFN366_n17753),
	.b(n20138));
   no02s02 U18837 (.o(n25459),
	.a(west_output_space_valid_f),
	.b(n25436));
   no02s02 U18838 (.o(n25374),
	.a(north_output_space_valid_f),
	.b(n25351));
   no02f02 U18839 (.o(n23308),
	.a(south_input_control_count_f_4_),
	.b(n23309));
   no02f20 U18840 (.o(n26014),
	.a(n20504),
	.b(n19494));
   no02f04 U18841 (.o(n17831),
	.a(n20450),
	.b(n20448));
   no02f02 U18842 (.o(n17872),
	.a(n20110),
	.b(n17871));
   oa22f10 U18843 (.o(n25000),
	.a(FE_RN_6),
	.b(n19871),
	.c(n19801),
	.d(n19800));
   in01f08 U18844 (.o(n25295),
	.a(n25027));
   no02f10 U18845 (.o(n18212),
	.a(n20222),
	.b(n20221));
   na02f10 U18846 (.o(n19067),
	.a(n19066),
	.b(n20267));
   in01f02 U18847 (.o(n19069),
	.a(n19066));
   no02f10 U18848 (.o(n26015),
	.a(n20504),
	.b(n19473));
   na02f04 U18849 (.o(n20513),
	.a(FE_OFN526_n24731),
	.b(n20349));
   in01f06 U18851 (.o(n17870),
	.a(n20110));
   no02f03 U18852 (.o(n17830),
	.a(n20448),
	.b(n20443));
   na02f02 U18853 (.o(n20438),
	.a(n20437),
	.b(n20436));
   na02f03 U18855 (.o(n20517),
	.a(n20320),
	.b(n23397));
   no03f04 U18856 (.o(n20257),
	.a(n20256),
	.b(n21907),
	.c(FE_OCPN25816_n20147));
   no02m04 U18857 (.o(n25974),
	.a(reset),
	.b(validIn_P));
   no02m01 U18858 (.o(n19068),
	.a(n25019),
	.b(n25061));
   no02m01 U18859 (.o(n18393),
	.a(n21695),
	.b(n20528));
   no03m02 U18860 (.o(n25723),
	.a(ec_thanks_e_to_p_reg),
	.b(ec_thanks_w_to_p_reg),
	.c(n25721));
   na02f10 U18861 (.o(n20267),
	.a(n20464),
	.b(n19065));
   in01f01 U18862 (.o(n20349),
	.a(n20528));
   no03f03 U18864 (.o(n20219),
	.a(n20217),
	.b(n20216),
	.c(n20368));
   na02f08 U18865 (.o(n18395),
	.a(n19474),
	.b(n20377));
   na02f02 U18866 (.o(n17871),
	.a(n18305),
	.b(n19252));
   ao12f08 U18867 (.o(n25017),
	.a(n19952),
	.b(n19953),
	.c(n21908));
   na02f03 U18868 (.o(n25117),
	.a(n20464),
	.b(n20463));
   no02f10 U18869 (.o(n25979),
	.a(reset),
	.b(n25978));
   ao12f20 U18870 (.o(n18074),
	.a(FE_OCPN25816_n20147),
	.b(n19477),
	.c(n19478));
   in01f01 U18872 (.o(n19519),
	.a(n19543));
   na02f02 U18873 (.o(n20218),
	.a(n20381),
	.b(n20369));
   oa22f02 U18874 (.o(n19976),
	.a(south_input_control_thanks_all_f),
	.b(south_input_control_tail_last_f),
	.c(south_input_control_count_one_f),
	.d(n20563));
   no02f03 U18875 (.o(n20630),
	.a(west_input_control_count_f_0_),
	.b(n20566));
   in01f04 U18876 (.o(n20220),
	.a(n20215));
   no02f04 U18877 (.o(n19462),
	.a(FE_OFN393_n19446),
	.b(n20528));
   no02f03 U18878 (.o(n20442),
	.a(n20437),
	.b(n20377));
   na02f01 U18879 (.o(n20446),
	.a(n20444),
	.b(n21426));
   no02m01 U18881 (.o(n20320),
	.a(n23398),
	.b(n20318));
   na02f03 U18882 (.o(n20145),
	.a(n20144),
	.b(n20143));
   in01f03 U18883 (.o(n19480),
	.a(n19479));
   in01f04 U18884 (.o(n20271),
	.a(n20417));
   na02f10 U18885 (.o(n19030),
	.a(n20417),
	.b(n19833));
   na02f10 U18886 (.o(n19029),
	.a(n19028),
	.b(n19027));
   in01f06 U18887 (.o(n25498),
	.a(n22518));
   in01f08 U18888 (.o(n19493),
	.a(FE_OFN247_n24982));
   in01f02 U18889 (.o(n19541),
	.a(n19562));
   no02f06 U18890 (.o(n20217),
	.a(n20365),
	.b(n18629));
   no02f06 U18891 (.o(n20149),
	.a(FE_RN_6),
	.b(n20211));
   no02f01 U18892 (.o(n20156),
	.a(n20167),
	.b(n20155));
   no03f10 U18893 (.o(n19477),
	.a(n19443),
	.b(n19804),
	.c(n19442));
   no02f02 U18894 (.o(n20200),
	.a(n20203),
	.b(n19549));
   in01f01 U18897 (.o(n19565),
	.a(n19738));
   in01s01 U18898 (.o(n20159),
	.a(n20158));
   in01f02 U18899 (.o(n24993),
	.a(n19834));
   in01f01 U18901 (.o(n21688),
	.a(proc_input_control_thanks_all_f));
   ao12f03 U18902 (.o(n20006),
	.a(n20004),
	.b(west_input_control_thanks_all_f),
	.c(n20005));
   in01f06 U18903 (.o(n19478),
	.a(n19476));
   na02f02 U18904 (.o(n17808),
	.a(n17810),
	.b(n17809));
   no04f04 U18905 (.o(n19823),
	.a(n20241),
	.b(n20240),
	.c(n19822),
	.d(n19821));
   no02f02 U18906 (.o(n19065),
	.a(n20463),
	.b(n19064));
   na02f01 U18907 (.o(n19847),
	.a(FE_OFN67_n19548),
	.b(n23968));
   in01f02 U18908 (.o(n22061),
	.a(proc_output_space_valid_f));
   no02f08 U18909 (.o(n18008),
	.a(n20104),
	.b(n20105));
   no02s02 U18910 (.o(n23398),
	.a(n18449),
	.b(n18447));
   no02m02 U18911 (.o(n20350),
	.a(west_output_control_planned_f),
	.b(n20377));
   no03f02 U18913 (.o(n19063),
	.a(n19062),
	.b(north_output_space_is_two_or_more_f),
	.c(north_output_space_yummy_f));
   in01f06 U18914 (.o(n19443),
	.a(n19825));
   na02f06 U18915 (.o(n18137),
	.a(n25020),
	.b(FE_RN_4));
   in01f02 U18916 (.o(n17809),
	.a(n20301));
   in01m06 U18917 (.o(n20343),
	.a(south_output_control_planned_f));
   no02f06 U18918 (.o(n20233),
	.a(n20181),
	.b(n19879));
   oa22f08 U18919 (.o(n19740),
	.a(FE_OFN65_n19542),
	.b(n23189),
	.c(FE_OFN63_n19518),
	.d(n22931));
   no03f06 U18920 (.o(n18885),
	.a(n18964),
	.b(n18967),
	.c(n20439));
   in01f02 U18921 (.o(n19809),
	.a(n19803));
   oa12f08 U18922 (.o(n20251),
	.a(n19785),
	.b(n20241),
	.c(n19329));
   na02f08 U18923 (.o(n20105),
	.a(n23628),
	.b(n23956));
   ao12m02 U18924 (.o(n23711),
	.a(south_output_space_is_two_or_more_f),
	.b(n19251),
	.c(n20493));
   na02f06 U18925 (.o(n19442),
	.a(n19794),
	.b(n19817));
   no02f08 U18926 (.o(n25506),
	.a(n19018),
	.b(n19021));
   no02f01 U18927 (.o(n19062),
	.a(north_output_space_valid_f),
	.b(n19061));
   na02f04 U18928 (.o(n23958),
	.a(n19964),
	.b(n19963));
   oa12f10 U18929 (.o(n20466),
	.a(n19853),
	.b(n19048),
	.c(n19047));
   in01f01 U18930 (.o(n20176),
	.a(n20166));
   no02m02 U18931 (.o(n17810),
	.a(n20299),
	.b(n20394));
   in01f01 U18932 (.o(n20248),
	.a(n20247));
   oa22f01 U18933 (.o(n17865),
	.a(n21864),
	.b(n19890),
	.c(n19225),
	.d(n19891));
   na02f04 U18934 (.o(n23620),
	.a(n19907),
	.b(n19908));
   na02f04 U18935 (.o(n24028),
	.a(n19970),
	.b(n19969));
   na04f04 U18936 (.o(n20017),
	.a(n20016),
	.b(n20015),
	.c(n20014),
	.d(n20013));
   no02f01 U18937 (.o(n18449),
	.a(east_output_space_valid_f),
	.b(n18450));
   in01s01 U18938 (.o(n18447),
	.a(n18448));
   ao22m02 U18939 (.o(n19905),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__26_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__26_));
   ao22m02 U18940 (.o(n19901),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__29_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__29_));
   in01f06 U18941 (.o(n20241),
	.a(n19795));
   ao22m02 U18942 (.o(n19968),
	.a(n24472),
	.b(south_input_NIB_storage_data_f_0__28_),
	.c(FE_RN_17),
	.d(south_input_NIB_storage_data_f_2__28_));
   in01m02 U18943 (.o(n20415),
	.a(n19828));
   na02f01 U18944 (.o(n19893),
	.a(n24364),
	.b(north_input_NIB_storage_data_f_1__22_));
   in01f04 U18945 (.o(n19033),
	.a(n19032));
   na02f01 U18946 (.o(n19892),
	.a(FE_RN_11),
	.b(north_input_NIB_storage_data_f_2__22_));
   na03f06 U18947 (.o(n18386),
	.a(n19716),
	.b(n19715),
	.c(myLocX_f_0_));
   in01f10 U18948 (.o(n18101),
	.a(n18100));
   oa22f08 U18949 (.o(n20240),
	.a(n19725),
	.b(n19413),
	.c(n19729),
	.d(n19412));
   oa12f10 U18950 (.o(n19047),
	.a(FE_RN_22),
	.b(n19043),
	.c(n19042));
   no02f04 U18951 (.o(n25003),
	.a(n19300),
	.b(n19299));
   no02f08 U18952 (.o(n19735),
	.a(myLocX_f_0_),
	.b(n22850));
   na02f02 U18953 (.o(n19459),
	.a(n25152),
	.b(proc_input_valid));
   no02f06 U18954 (.o(n19824),
	.a(n19789),
	.b(n19788));
   na02f10 U18955 (.o(n19630),
	.a(myChipID_f_8_),
	.b(n19629));
   na02f10 U18956 (.o(n23482),
	.a(n19783),
	.b(n19782));
   ao22f02 U18957 (.o(n19024),
	.a(n19017),
	.b(east_input_valid),
	.c(n19019),
	.d(west_input_valid));
   no02f08 U18959 (.o(n24036),
	.a(n20103),
	.b(n20102));
   ao22f01 U18960 (.o(n19978),
	.a(n18959),
	.b(west_input_NIB_storage_data_f_3__22_),
	.c(n18828),
	.d(west_input_NIB_storage_data_f_1__22_));
   ao22f02 U18961 (.o(n19964),
	.a(FE_OCPN25942_n24965),
	.b(south_input_NIB_storage_data_f_3__29_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__29_));
   ao22m02 U18962 (.o(n19902),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__29_),
	.c(FE_OFN24770_n19075),
	.d(north_input_NIB_storage_data_f_0__29_));
   ao22m02 U18963 (.o(n19908),
	.a(FE_OFN51_n19193),
	.b(north_input_NIB_storage_data_f_3__23_),
	.c(FE_OFN24770_n19075),
	.d(north_input_NIB_storage_data_f_0__23_));
   ao22f04 U18964 (.o(n20011),
	.a(proc_input_NIB_storage_data_f_7__22_),
	.b(FE_OFN20_n17779),
	.c(proc_input_NIB_storage_data_f_5__22_),
	.d(FE_RN_49));
   in01f01 U18965 (.o(n19414),
	.a(n19411));
   no02f10 U18966 (.o(n23956),
	.a(n20072),
	.b(n20071));
   ao22m02 U18967 (.o(n20015),
	.a(proc_input_NIB_storage_data_f_11__22_),
	.b(FE_OCPN25909_n19547),
	.c(proc_input_NIB_storage_data_f_15__22_),
	.d(n24065));
   ao22f01 U18968 (.o(n20013),
	.a(n19705),
	.b(proc_input_NIB_storage_data_f_9__22_),
	.c(FE_OFN169_n24343),
	.d(proc_input_NIB_storage_data_f_8__22_));
   no02f10 U18969 (.o(n24998),
	.a(n19767),
	.b(n19766));
   na02f06 U18970 (.o(n19829),
	.a(n20272),
	.b(n20285));
   no02f04 U18971 (.o(n20032),
	.a(n20024),
	.b(n20023));
   no02f04 U18972 (.o(n20062),
	.a(n20053),
	.b(n20052));
   na02f04 U18973 (.o(n19283),
	.a(n20245),
	.b(n19787));
   ao22m02 U18975 (.o(n19913),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__22_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__22_));
   in01f03 U18977 (.o(n20514),
	.a(west_output_control_planned_f));
   ao22f01 U18978 (.o(n20014),
	.a(FE_OFN156_n24129),
	.b(proc_input_NIB_storage_data_f_1__22_),
	.c(n17742),
	.d(proc_input_NIB_storage_data_f_4__22_));
   ao22f02 U18979 (.o(n18550),
	.a(proc_input_valid),
	.b(n25521),
	.c(south_input_valid),
	.d(n19059));
   na02f06 U18980 (.o(n19853),
	.a(n19046),
	.b(n19045));
   no02f02 U18981 (.o(n25020),
	.a(n18813),
	.b(n24992));
   no02f01 U18982 (.o(n19451),
	.a(west_output_space_is_two_or_more_f),
	.b(west_output_space_yummy_f));
   na02f02 U18983 (.o(n18549),
	.a(west_input_valid),
	.b(n19057));
   na02f01 U18984 (.o(n19840),
	.a(n19326),
	.b(n20911));
   na02f02 U18985 (.o(n19450),
	.a(west_output_space_is_one_f),
	.b(n19447));
   ao22m02 U18986 (.o(n19912),
	.a(FE_OFN24777_n19932),
	.b(east_input_NIB_storage_data_f_0__22_),
	.c(n19400),
	.d(east_input_NIB_storage_data_f_3__22_));
   in01s01 U18987 (.o(n18450),
	.a(east_output_space_is_one_f));
   na02s02 U18988 (.o(n20493),
	.a(south_output_space_valid_f),
	.b(n19250));
   no02m01 U18989 (.o(n18448),
	.a(east_output_space_yummy_f),
	.b(east_output_space_is_two_or_more_f));
   in01f08 U18990 (.o(n19042),
	.a(n19041));
   in01f02 U18991 (.o(n19412),
	.a(n22819));
   in01f02 U18992 (.o(n19413),
	.a(n22858));
   oa22f01 U18993 (.o(n19300),
	.a(FE_OFN25664_n19914),
	.b(n19297),
	.c(n20506),
	.d(n19296));
   oa22f01 U18994 (.o(n19299),
	.a(n21858),
	.b(n19298),
	.c(n19435),
	.d(n24787));
   na02f04 U18995 (.o(n24030),
	.a(n19941),
	.b(n19940));
   na02f04 U18996 (.o(n23623),
	.a(n19945),
	.b(n19944));
   no03f10 U18997 (.o(n22826),
	.a(n19728),
	.b(n19727),
	.c(n19726));
   no03f06 U18998 (.o(n18464),
	.a(n21509),
	.b(n19584),
	.c(n21508));
   in01f02 U18999 (.o(n19247),
	.a(n19246));
   ao22m02 U19000 (.o(n19308),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__31_),
	.c(FE_OFN24777_n19932),
	.d(east_input_NIB_storage_data_f_0__31_));
   no02f01 U19001 (.o(n18339),
	.a(FE_OFN24745_n18648),
	.b(n18340));
   no03f06 U19002 (.o(n18024),
	.a(n18076),
	.b(n19600),
	.c(n19617));
   na04f08 U19003 (.o(n19767),
	.a(n19761),
	.b(n19760),
	.c(n19759),
	.d(n19758));
   na04f08 U19004 (.o(n19766),
	.a(n19765),
	.b(n19764),
	.c(n19763),
	.d(n19762));
   no02f08 U19006 (.o(n20160),
	.a(n19137),
	.b(n20173));
   ao22f04 U19007 (.o(n19008),
	.a(myLocY_f_0_),
	.b(FE_OFN25615_n19007),
	.c(n19007),
	.d(n19325));
   no02f10 U19008 (.o(n18104),
	.a(n19546),
	.b(n19545));
   na04f08 U19009 (.o(n20071),
	.a(n20070),
	.b(n20069),
	.c(n20068),
	.d(n20067));
   na02f08 U19010 (.o(n19039),
	.a(n19038),
	.b(n19041));
   na02f02 U19012 (.o(n18813),
	.a(n19834),
	.b(n18803));
   in01f01 U19013 (.o(n18474),
	.a(n20181));
   no02f02 U19014 (.o(n18133),
	.a(n20211),
	.b(n22912));
   in01f01 U19015 (.o(west_input_valid),
	.a(n19453));
   ao22f10 U19016 (.o(n19439),
	.a(myLocY_f_4_),
	.b(n22881),
	.c(myLocY_f_3_),
	.d(n22874));
   no02f20 U19017 (.o(n19057),
	.a(north_output_current_route_connection_2_),
	.b(n25127));
   in01s01 U19018 (.o(n19447),
	.a(west_output_space_valid_f));
   no02f06 U19019 (.o(n20244),
	.a(myLocX_f_1_),
	.b(n21469));
   na02f08 U19020 (.o(n18117),
	.a(n19841),
	.b(n19038));
   no02f20 U19021 (.o(n19019),
	.a(east_output_current_route_connection_0_),
	.b(n19018));
   na02f08 U19022 (.o(n20245),
	.a(myLocX_f_1_),
	.b(n21469));
   na02f04 U19023 (.o(n20166),
	.a(n20158),
	.b(n19129));
   no02m02 U19024 (.o(n19323),
	.a(myLocY_f_0_),
	.b(n22827));
   no03f10 U19025 (.o(n19054),
	.a(north_output_current_route_connection_2_),
	.b(n25130),
	.c(n25138));
   na02f04 U19026 (.o(n19788),
	.a(n19787),
	.b(n19786));
   na02f02 U19027 (.o(n19255),
	.a(n25499),
	.b(proc_input_valid));
   ao22f04 U19028 (.o(n20070),
	.a(FE_OCPN25933_n24342),
	.b(proc_input_NIB_storage_data_f_0__28_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__28_));
   ao22f02 U19029 (.o(n20080),
	.a(FE_OCPN25933_n24342),
	.b(proc_input_NIB_storage_data_f_0__23_),
	.c(FE_OCPN25908_n19547),
	.d(proc_input_NIB_storage_data_f_11__23_));
   ao22m02 U19030 (.o(n20036),
	.a(FE_OCPN25825_n21745),
	.b(proc_input_NIB_storage_data_f_2__25_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__25_));
   na02f01 U19031 (.o(n19981),
	.a(FE_RN_31),
	.b(west_input_NIB_storage_data_f_1__27_));
   ao22f02 U19032 (.o(n19899),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__28_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__28_));
   ao22f02 U19033 (.o(n19900),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__28_),
	.c(FE_OFN24770_n19075),
	.d(north_input_NIB_storage_data_f_0__28_));
   ao22f02 U19034 (.o(n20074),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__23_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__23_));
   ao22m02 U19035 (.o(n20028),
	.a(FE_OFN156_n24129),
	.b(proc_input_NIB_storage_data_f_1__26_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__26_));
   ao22f02 U19036 (.o(n19987),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__25_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__25_));
   ao22m02 U19037 (.o(n20058),
	.a(FE_OFN167_n24343),
	.b(proc_input_NIB_storage_data_f_8__27_),
	.c(n17742),
	.d(proc_input_NIB_storage_data_f_4__27_));
   ao22f02 U19038 (.o(n19895),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__24_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__24_));
   ao22f02 U19039 (.o(n20025),
	.a(proc_input_NIB_storage_data_f_0__26_),
	.b(FE_OCPN25933_n24342),
	.c(proc_input_NIB_storage_data_f_15__26_),
	.d(FE_OFN25637_n19595));
   ao22f02 U19040 (.o(n19898),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__27_),
	.c(FE_OFN24770_n19075),
	.d(north_input_NIB_storage_data_f_0__27_));
   ao22m02 U19041 (.o(n20033),
	.a(FE_RN_35),
	.b(proc_input_NIB_storage_data_f_12__25_),
	.c(FE_OFN191_n24454),
	.d(proc_input_NIB_storage_data_f_13__25_));
   ao22f02 U19042 (.o(n20076),
	.a(proc_input_NIB_storage_data_f_7__23_),
	.b(n17779),
	.c(proc_input_NIB_storage_data_f_5__23_),
	.d(FE_RN_49));
   ao22f02 U19043 (.o(n19761),
	.a(proc_input_NIB_storage_data_f_7__31_),
	.b(FE_OFN20_n17779),
	.c(proc_input_NIB_storage_data_f_5__31_),
	.d(FE_RN_49));
   ao22m02 U19044 (.o(n20021),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__26_),
	.c(n20012),
	.d(proc_input_NIB_storage_data_f_9__26_));
   ao22f02 U19046 (.o(n19764),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__31_),
	.c(FE_OCPN25948_n19595),
	.d(proc_input_NIB_storage_data_f_15__31_));
   ao22f02 U19047 (.o(n19759),
	.a(FE_RN_38),
	.b(proc_input_NIB_storage_data_f_2__31_),
	.c(FE_OCPN25918_n19547),
	.d(proc_input_NIB_storage_data_f_11__31_));
   ao22f02 U19048 (.o(n19989),
	.a(FE_OFN24764_n18960),
	.b(west_input_NIB_storage_data_f_2__26_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__26_));
   ao22f02 U19049 (.o(n20083),
	.a(n18051),
	.b(proc_input_NIB_storage_data_f_10__29_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__29_));
   ao22f02 U19050 (.o(n19896),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__24_),
	.c(FE_OFN24770_n19075),
	.d(north_input_NIB_storage_data_f_0__24_));
   ao22f02 U19052 (.o(n20085),
	.a(proc_input_NIB_storage_data_f_0__29_),
	.b(FE_OCPN25933_n24342),
	.c(proc_input_NIB_storage_data_f_5__29_),
	.d(FE_RN_49));
   na02f06 U19053 (.o(n20272),
	.a(n19720),
	.b(n23293));
   na02f08 U19054 (.o(n19828),
	.a(myLocX_f_7_),
	.b(n22822));
   ao22f08 U19055 (.o(n20303),
	.a(n22860),
	.b(myLocX_f_6_),
	.c(myLocX_f_7_),
	.d(n22821));
   ao22f04 U19056 (.o(n19322),
	.a(n19326),
	.b(n20912),
	.c(FE_OFN67_n19548),
	.d(n23965));
   ao22m02 U19057 (.o(n20050),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__27_),
	.c(FE_OFN25633_n19595),
	.d(proc_input_NIB_storage_data_f_15__27_));
   ao22f08 U19059 (.o(n20279),
	.a(n23303),
	.b(n19719),
	.c(n19706),
	.d(n23503));
   ao22f02 U19060 (.o(n19763),
	.a(FE_OFN161_n24129),
	.b(proc_input_NIB_storage_data_f_1__31_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__31_));
   no02f10 U19061 (.o(n20389),
	.a(n19208),
	.b(n20299));
   na02f08 U19062 (.o(n18388),
	.a(n19711),
	.b(n19717));
   in01m03 U19063 (.o(n18390),
	.a(n19712));
   ao22f02 U19064 (.o(n19765),
	.a(n19707),
	.b(proc_input_NIB_storage_data_f_3__31_),
	.c(n19769),
	.d(proc_input_NIB_storage_data_f_14__31_));
   in01m04 U19065 (.o(n20462),
	.a(n19055));
   in01f02 U19066 (.o(n19128),
	.a(n19127));
   ao22f02 U19067 (.o(n19897),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__27_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__27_));
   na02f10 U19070 (.o(n20263),
	.a(n20444),
	.b(n20196));
   oa22m02 U19071 (.o(n19254),
	.a(n19453),
	.b(n24982),
	.c(n19452),
	.d(n22517));
   na02f06 U19072 (.o(n19329),
	.a(n19720),
	.b(n23292));
   ao22m02 U19073 (.o(n20099),
	.a(n24343),
	.b(proc_input_NIB_storage_data_f_8__24_),
	.c(proc_input_NIB_storage_data_f_3__24_),
	.d(n19709));
   na02f08 U19074 (.o(n19728),
	.a(n19673),
	.b(n19672));
   no02f10 U19075 (.o(n17899),
	.a(n17903),
	.b(n17900));
   ao12f02 U19076 (.o(n20069),
	.a(n17910),
	.b(proc_input_NIB_storage_data_f_1__28_),
	.c(FE_OFN156_n24129));
   na02f06 U19077 (.o(n19724),
	.a(n19681),
	.b(n19680));
   no02f10 U19078 (.o(n17819),
	.a(n17821),
	.b(n17820));
   na03f06 U19079 (.o(n21522),
	.a(n19143),
	.b(n19142),
	.c(n19141));
   ao22f02 U19080 (.o(n20096),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__24_),
	.c(FE_OFN188_n24453),
	.d(proc_input_NIB_storage_data_f_2__24_));
   ao22m02 U19081 (.o(n19941),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__24_),
	.c(n19400),
	.d(east_input_NIB_storage_data_f_3__24_));
   in01f04 U19082 (.o(n18529),
	.a(n19586));
   ao22m02 U19083 (.o(n20089),
	.a(n17747),
	.b(proc_input_NIB_storage_data_f_12__29_),
	.c(FE_OFN25604_n19530),
	.d(proc_input_NIB_storage_data_f_13__29_));
   na02f06 U19084 (.o(n22773),
	.a(n20356),
	.b(n20538));
   no02f08 U19085 (.o(n21469),
	.a(n19262),
	.b(n19261));
   na02f02 U19086 (.o(n19787),
	.a(myLocX_f_0_),
	.b(n22843));
   in01f04 U19087 (.o(n25138),
	.a(north_output_current_route_connection_0_));
   no02f08 U19088 (.o(n19246),
	.a(n23035),
	.b(n20408));
   na02f04 U19089 (.o(n19805),
	.a(n19321),
	.b(n19421));
   na02f01 U19090 (.o(n19982),
	.a(FE_OFN28_n18974),
	.b(west_input_NIB_storage_data_f_0__27_));
   no02f10 U19091 (.o(n20301),
	.a(n19232),
	.b(n20388));
   no02f20 U19092 (.o(n18383),
	.a(n18528),
	.b(n18532));
   in01m04 U19093 (.o(n19021),
	.a(east_output_current_route_connection_0_));
   na02f02 U19094 (.o(n19481),
	.a(west_output_current_route_connection_0_),
	.b(n25176));
   na02f01 U19095 (.o(n19984),
	.a(FE_OFN24764_n18960),
	.b(west_input_NIB_storage_data_f_2__27_));
   ao22f02 U19096 (.o(n20040),
	.a(FE_OCPN25933_n24342),
	.b(proc_input_NIB_storage_data_f_0__25_),
	.c(FE_OCPN25911_n19547),
	.d(proc_input_NIB_storage_data_f_11__25_));
   ao22f02 U19097 (.o(n19990),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__26_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__26_));
   in01f10 U19098 (.o(n19399),
	.a(n23316));
   na02f01 U19099 (.o(n19983),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__27_));
   ao22f02 U19100 (.o(n20027),
	.a(n24343),
	.b(proc_input_NIB_storage_data_f_8__26_),
	.c(n17743),
	.d(proc_input_NIB_storage_data_f_4__26_));
   ao22f02 U19101 (.o(n20048),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__27_),
	.c(FE_OFN20_n17779),
	.d(proc_input_NIB_storage_data_f_7__27_));
   no02f04 U19102 (.o(n19137),
	.a(n19133),
	.b(n20169));
   na02f04 U19103 (.o(n20390),
	.a(n19720),
	.b(n23294));
   na02f08 U19104 (.o(n19280),
	.a(n19719),
	.b(FE_RN_61));
   ao22f03 U19105 (.o(n19762),
	.a(FE_OCPN25955_n18039),
	.b(proc_input_NIB_storage_data_f_10__31_),
	.c(FE_OFN167_n24343),
	.d(proc_input_NIB_storage_data_f_8__31_));
   ao22f02 U19106 (.o(n20077),
	.a(n19705),
	.b(proc_input_NIB_storage_data_f_9__23_),
	.c(FE_OFN25668_n18038),
	.d(proc_input_NIB_storage_data_f_10__23_));
   oa22f08 U19107 (.o(n20173),
	.a(myLocY_f_6_),
	.b(n23185),
	.c(myLocY_f_5_),
	.d(n22853));
   na02f06 U19109 (.o(n20285),
	.a(myLocX_f_6_),
	.b(n22861));
   na02f01 U19110 (.o(n19916),
	.a(FE_RN_69),
	.b(east_input_NIB_storage_data_f_1__26_));
   no02m02 U19111 (.o(n19881),
	.a(myLocY_f_0_),
	.b(FE_OFN25616_n19007));
   ao22f02 U19112 (.o(n20047),
	.a(n21739),
	.b(proc_input_NIB_storage_data_f_12__27_),
	.c(FE_OFN191_n24454),
	.d(proc_input_NIB_storage_data_f_13__27_));
   ao22f02 U19113 (.o(n20090),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__29_),
	.c(FE_OFN156_n24129),
	.d(proc_input_NIB_storage_data_f_1__29_));
   ao22f02 U19114 (.o(n20078),
	.a(FE_OFN169_n24343),
	.b(proc_input_NIB_storage_data_f_8__23_),
	.c(n17744),
	.d(proc_input_NIB_storage_data_f_4__23_));
   ao22m02 U19116 (.o(n19750),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__32_),
	.c(proc_input_NIB_storage_data_f_15__32_),
	.d(FE_OFN25637_n19595));
   ao22f08 U19117 (.o(n19579),
	.a(FE_OCPN25968_n19500),
	.b(proc_input_NIB_storage_data_f_12__61_),
	.c(FE_OCPN25814_FE_OFN186_n24453),
	.d(proc_input_NIB_storage_data_f_2__61_));
   ao22f04 U19118 (.o(n19528),
	.a(FE_OCPN25824_n21745),
	.b(proc_input_NIB_storage_data_f_2__39_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__39_));
   ao22f04 U19119 (.o(n19674),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__49_),
	.c(FE_OFN25637_n19595),
	.d(proc_input_NIB_storage_data_f_15__49_));
   ao22f06 U19120 (.o(n19679),
	.a(FE_OCPN25933_n24342),
	.b(proc_input_NIB_storage_data_f_0__49_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__49_));
   na02f06 U19121 (.o(n18231),
	.a(proc_input_NIB_storage_data_f_2__62_),
	.b(FE_OCPN25814_FE_OFN186_n24453));
   no02f01 U19122 (.o(n17910),
	.a(FE_OFN24806_n19655),
	.b(n17911));
   ao22f06 U19123 (.o(n19532),
	.a(FE_OFN25604_n19530),
	.b(proc_input_NIB_storage_data_f_13__38_),
	.c(FE_OCPN25933_n24342),
	.d(proc_input_NIB_storage_data_f_0__38_));
   ao22f08 U19124 (.o(n18233),
	.a(proc_input_NIB_storage_data_f_6__62_),
	.b(n19503),
	.c(proc_input_NIB_storage_data_f_9__62_),
	.d(FE_OFN25681_n17814));
   ao22f04 U19126 (.o(n19687),
	.a(FE_OCPN25933_n24342),
	.b(proc_input_NIB_storage_data_f_0__48_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__48_));
   ao22f06 U19127 (.o(n19526),
	.a(FE_OFN25633_n19595),
	.b(proc_input_NIB_storage_data_f_15__39_),
	.c(n17744),
	.d(proc_input_NIB_storage_data_f_4__39_));
   ao22f04 U19128 (.o(n19716),
	.a(n17747),
	.b(proc_input_NIB_storage_data_f_12__42_),
	.c(FE_OFN25604_n19530),
	.d(proc_input_NIB_storage_data_f_13__42_));
   ao22f06 U19129 (.o(n19717),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__42_),
	.c(n24343),
	.d(proc_input_NIB_storage_data_f_8__42_));
   oa22f02 U19130 (.o(n19261),
	.a(n21857),
	.b(n24895),
	.c(n20506),
	.d(n19260));
   in01f10 U19131 (.o(n18910),
	.a(n21162));
   in01f08 U19132 (.o(n19364),
	.a(n21288));
   in01f10 U19133 (.o(n19397),
	.a(n21294));
   in01f03 U19134 (.o(n19729),
	.a(myLocX_f_7_));
   in01f10 U19135 (.o(n18176),
	.a(n18177));
   na03f10 U19136 (.o(n23503),
	.a(n18743),
	.b(n18745),
	.c(n18744));
   in01f03 U19137 (.o(n20463),
	.a(n20379));
   in01m03 U19138 (.o(n25163),
	.a(n19454));
   in01f06 U19140 (.o(n17826),
	.a(n19514));
   in01m10 U19141 (.o(n25130),
	.a(north_output_current_route_connection_1_));
   ao22f02 U19142 (.o(n19675),
	.a(n17779),
	.b(proc_input_NIB_storage_data_f_7__49_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__49_));
   ao22f08 U19143 (.o(n18066),
	.a(proc_input_NIB_storage_data_f_2__58_),
	.b(FE_OCPN25814_FE_OFN186_n24453),
	.c(proc_input_NIB_storage_data_f_12__58_),
	.d(FE_OCPN25968_n19500));
   ao22f06 U19144 (.o(n19531),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__38_),
	.c(FE_OFN169_n24343),
	.d(proc_input_NIB_storage_data_f_8__38_));
   no02f01 U19145 (.o(n17908),
	.a(FE_OFN24806_n19655),
	.b(n17909));
   no02f04 U19146 (.o(n19815),
	.a(myLocY_f_4_),
	.b(n22881));
   in01f04 U19147 (.o(n19327),
	.a(n22843));
   ao22f10 U19148 (.o(n18232),
	.a(proc_input_NIB_storage_data_f_0__62_),
	.b(FE_OCPN25970_n24342),
	.c(proc_input_NIB_storage_data_f_13__62_),
	.d(FE_OFN25602_n19530));
   ao22f08 U19149 (.o(n19576),
	.a(n20056),
	.b(proc_input_NIB_storage_data_f_9__61_),
	.c(FE_OFN165_n24129),
	.d(proc_input_NIB_storage_data_f_1__61_));
   ao22f06 U19150 (.o(n19685),
	.a(n24343),
	.b(proc_input_NIB_storage_data_f_8__48_),
	.c(n17743),
	.d(proc_input_NIB_storage_data_f_4__48_));
   ao22f06 U19151 (.o(n19686),
	.a(n19709),
	.b(proc_input_NIB_storage_data_f_3__48_),
	.c(FE_OFN156_n24129),
	.d(proc_input_NIB_storage_data_f_1__48_));
   no02f08 U19152 (.o(n20299),
	.a(n19708),
	.b(n23494));
   ao22f04 U19153 (.o(n19638),
	.a(n18131),
	.b(proc_input_NIB_storage_data_f_0__52_),
	.c(proc_input_NIB_storage_data_f_5__52_),
	.d(FE_RN_49));
   no02f10 U19154 (.o(n22853),
	.a(n18170),
	.b(n18169));
   oa22f08 U19155 (.o(n18586),
	.a(n19617),
	.b(n23509),
	.c(n19387),
	.d(n20745));
   na02f10 U19157 (.o(n18310),
	.a(n19658),
	.b(n19661));
   no02f06 U19158 (.o(n19208),
	.a(n19328),
	.b(n19230));
   oa22f08 U19159 (.o(n18328),
	.a(n23303),
	.b(n19719),
	.c(n19720),
	.d(n23293));
   na02f08 U19161 (.o(n17962),
	.a(n17964),
	.b(n17963));
   ao22f06 U19162 (.o(n19527),
	.a(n21739),
	.b(proc_input_NIB_storage_data_f_12__39_),
	.c(FE_OFN191_n24454),
	.d(proc_input_NIB_storage_data_f_13__39_));
   ao22f04 U19163 (.o(n19642),
	.a(FE_OFN24803_n19500),
	.b(proc_input_NIB_storage_data_f_12__52_),
	.c(n19769),
	.d(proc_input_NIB_storage_data_f_14__52_));
   no02f10 U19164 (.o(n20278),
	.a(myLocX_f_1_),
	.b(n18749));
   ao22f04 U19165 (.o(n19637),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__52_),
	.c(FE_RN_33),
	.d(proc_input_NIB_storage_data_f_3__52_));
   no02f10 U19166 (.o(n17805),
	.a(myLocX_f_5_),
	.b(n19294));
   no02f08 U19167 (.o(n19839),
	.a(FE_OFN67_n19548),
	.b(n23968));
   in01m02 U19168 (.o(n19856),
	.a(n19252));
   na02f02 U19169 (.o(n18792),
	.a(n25301),
	.b(proc_input_valid));
   no02f08 U19170 (.o(n19441),
	.a(myLocY_f_6_),
	.b(n23183));
   no02f06 U19171 (.o(n20266),
	.a(east_output_current_route_connection_2_),
	.b(east_output_current_route_connection_1_));
   no02f08 U19172 (.o(n19229),
	.a(myLocX_f_5_),
	.b(n19237));
   ao22f04 U19173 (.o(n19641),
	.a(FE_OCPN25947_n19595),
	.b(proc_input_NIB_storage_data_f_15__52_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__52_));
   no02f06 U19174 (.o(n19806),
	.a(FE_OFN67_n19548),
	.b(n23965));
   na02f06 U19175 (.o(n18161),
	.a(n18163),
	.b(n18162));
   no02f03 U19176 (.o(n25176),
	.a(west_output_current_route_connection_1_),
	.b(west_output_current_route_connection_2_));
   no02f04 U19177 (.o(n25153),
	.a(west_output_current_route_connection_1_),
	.b(west_output_current_route_connection_0_));
   ao22f06 U19178 (.o(n19535),
	.a(n19705),
	.b(proc_input_NIB_storage_data_f_9__38_),
	.c(n18035),
	.d(proc_input_NIB_storage_data_f_10__38_));
   na02f06 U19179 (.o(n18164),
	.a(n18166),
	.b(n18165));
   no02f08 U19181 (.o(n17839),
	.a(n17841),
	.b(n17840));
   ao22f06 U19182 (.o(n19639),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__52_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__52_));
   na02f08 U19183 (.o(n19036),
	.a(n18296),
	.b(n18294));
   no02f08 U19184 (.o(n18327),
	.a(n19328),
	.b(n18748));
   na02f04 U19185 (.o(n20182),
	.a(myLocY_f_0_),
	.b(FE_OFN25616_n19007));
   no02f01 U19186 (.o(n18425),
	.a(FE_RN_34),
	.b(n18426));
   na02f10 U19187 (.o(n19600),
	.a(n19597),
	.b(n19596));
   oa22f04 U19188 (.o(n18307),
	.a(n24244),
	.b(n17740),
	.c(FE_RN_53),
	.d(n17739));
   ao12f04 U19189 (.o(n20302),
	.a(myLocX_f_7_),
	.b(n19238),
	.c(n19239));
   na02f06 U19190 (.o(n21667),
	.a(n19861),
	.b(n20123));
   ao22f06 U19191 (.o(n19580),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__61_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__61_));
   ao22f04 U19192 (.o(n19715),
	.a(FE_OCPN25933_n24342),
	.b(proc_input_NIB_storage_data_f_0__42_),
	.c(FE_OFN25637_n19595),
	.d(proc_input_NIB_storage_data_f_15__42_));
   ao22f01 U19193 (.o(n19744),
	.a(n17747),
	.b(proc_input_NIB_storage_data_f_12__32_),
	.c(n19769),
	.d(proc_input_NIB_storage_data_f_14__32_));
   ao22f06 U19194 (.o(n19677),
	.a(n24343),
	.b(proc_input_NIB_storage_data_f_8__49_),
	.c(n17743),
	.d(proc_input_NIB_storage_data_f_4__49_));
   ao22f02 U19195 (.o(n19712),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__42_),
	.c(n19709),
	.d(proc_input_NIB_storage_data_f_3__42_));
   ao22f03 U19196 (.o(n19713),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__42_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__42_));
   ao22f04 U19197 (.o(n19533),
	.a(FE_RN_54),
	.b(proc_input_NIB_storage_data_f_12__38_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__38_));
   ao22f06 U19198 (.o(n19643),
	.a(FE_OCPN25814_FE_OFN186_n24453),
	.b(proc_input_NIB_storage_data_f_2__52_),
	.c(FE_OFN165_n24129),
	.d(proc_input_NIB_storage_data_f_1__52_));
   in01f02 U19199 (.o(n19143),
	.a(n19138));
   in01m02 U19200 (.o(n20538),
	.a(west_output_current_route_connection_1_));
   na02f04 U19201 (.o(n18018),
	.a(FE_OCPN25924_n19547),
	.b(proc_input_NIB_storage_data_f_11__62_));
   ao22f02 U19202 (.o(n19711),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__42_),
	.c(n17743),
	.d(proc_input_NIB_storage_data_f_4__42_));
   ao12f01 U19203 (.o(n19777),
	.a(n17928),
	.b(proc_input_NIB_storage_data_f_6__30_),
	.c(n19503));
   na02f04 U19204 (.o(n18227),
	.a(proc_input_NIB_storage_data_f_1__62_),
	.b(FE_OFN165_n24129));
   na02f04 U19205 (.o(n20184),
	.a(myLocY_f_3_),
	.b(n22875));
   no02f06 U19206 (.o(n19119),
	.a(n19326),
	.b(n19123));
   na02f04 U19207 (.o(n18088),
	.a(n23184),
	.b(myLocY_f_6_));
   na02f04 U19208 (.o(n18019),
	.a(FE_OCPN25962_n18039),
	.b(proc_input_NIB_storage_data_f_10__62_));
   ao22f04 U19209 (.o(n19524),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__39_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__39_));
   no02m08 U19210 (.o(n19015),
	.a(east_output_current_route_connection_1_),
	.b(east_output_current_route_connection_0_));
   na02f04 U19211 (.o(n20183),
	.a(myLocY_f_1_),
	.b(n22836));
   oa22f02 U19212 (.o(n19262),
	.a(FE_OFN25664_n19914),
	.b(n19259),
	.c(n21858),
	.d(n19258));
   no02f08 U19213 (.o(n19842),
	.a(n19326),
	.b(n20911));
   na02f20 U19214 (.o(n18530),
	.a(n19590),
	.b(n19593));
   ao22f01 U19215 (.o(n19747),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__32_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__32_));
   na02f08 U19216 (.o(n20737),
	.a(north_input_valid),
	.b(n20618));
   na02f10 U19217 (.o(n20185),
	.a(myLocY_f_2_),
	.b(n19009));
   no02m08 U19218 (.o(n25123),
	.a(north_output_current_route_connection_2_),
	.b(north_output_current_route_connection_0_));
   no02f06 U19219 (.o(n19055),
	.a(north_output_current_route_connection_1_),
	.b(north_output_current_route_connection_0_));
   ao22f06 U19220 (.o(n17898),
	.a(proc_input_NIB_storage_data_f_6__55_),
	.b(n19503),
	.c(proc_input_NIB_storage_data_f_0__55_),
	.d(FE_OCPN25839_n24342));
   na02f08 U19221 (.o(n18412),
	.a(proc_input_NIB_storage_data_f_1__57_),
	.b(FE_OFN161_n24129));
   ao22f04 U19222 (.o(n18486),
	.a(proc_input_NIB_storage_data_f_8__35_),
	.b(FE_OFN169_n24343),
	.c(proc_input_NIB_storage_data_f_9__35_),
	.d(n19705));
   na02f06 U19223 (.o(n17970),
	.a(proc_input_NIB_storage_data_f_3__59_),
	.b(n17754));
   ao22f04 U19224 (.o(n18316),
	.a(proc_input_NIB_storage_data_f_12__41_),
	.b(FE_OCPN25832_n19500),
	.c(proc_input_NIB_storage_data_f_6__41_),
	.d(n19503));
   ao22f04 U19225 (.o(n19316),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__35_),
	.c(FE_OFN24777_n19932),
	.d(east_input_NIB_storage_data_f_0__35_));
   ao22f10 U19226 (.o(n19509),
	.a(FE_OCPN25968_n19500),
	.b(proc_input_NIB_storage_data_f_12__40_),
	.c(n19654),
	.d(proc_input_NIB_storage_data_f_0__40_));
   no02f06 U19227 (.o(n19371),
	.a(FE_RN_57),
	.b(n24785));
   ao22f04 U19228 (.o(n17875),
	.a(FE_OCPN25913_n19547),
	.b(proc_input_NIB_storage_data_f_11__36_),
	.c(FE_OFN20_n17779),
	.d(proc_input_NIB_storage_data_f_7__36_));
   na02f04 U19229 (.o(n17961),
	.a(proc_input_NIB_storage_data_f_9__59_),
	.b(FE_OFN25681_n17814));
   ao22f08 U19230 (.o(n19603),
	.a(FE_RN_33),
	.b(proc_input_NIB_storage_data_f_3__63_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__63_));
   ao22f20 U19231 (.o(n19589),
	.a(n24454),
	.b(proc_input_NIB_storage_data_f_13__51_),
	.c(n17741),
	.d(proc_input_NIB_storage_data_f_4__51_));
   na02f03 U19232 (.o(n17983),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__50_));
   ao22f06 U19233 (.o(n19319),
	.a(FE_OFN24777_n19932),
	.b(east_input_NIB_storage_data_f_0__37_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__37_));
   ao22f10 U19234 (.o(n19362),
	.a(FE_OFN24780_n19932),
	.b(east_input_NIB_storage_data_f_0__61_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__61_));
   in01f10 U19236 (.o(n22884),
	.a(n18716));
   in01f06 U19237 (.o(n19009),
	.a(n23966));
   in01f04 U19239 (.o(n18878),
	.a(n18875));
   ao22f08 U19240 (.o(n18166),
	.a(proc_input_NIB_storage_data_f_4__56_),
	.b(n21749),
	.c(proc_input_NIB_storage_data_f_12__56_),
	.d(FE_OCPN25968_n19500));
   in01f10 U19241 (.o(n19594),
	.a(myChipID_f_1_));
   na02f04 U19242 (.o(n17958),
	.a(proc_input_NIB_storage_data_f_11__59_),
	.b(FE_OFN25673_n18033));
   ao22f10 U19243 (.o(n19510),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__40_),
	.c(FE_OFN20_n17779),
	.d(proc_input_NIB_storage_data_f_7__40_));
   na02f08 U19244 (.o(n23968),
	.a(n18704),
	.b(n18705));
   ao22f06 U19245 (.o(n17901),
	.a(proc_input_NIB_storage_data_f_12__55_),
	.b(FE_OFN24803_n19500),
	.c(proc_input_NIB_storage_data_f_4__55_),
	.d(n21749));
   in01f04 U19246 (.o(n18877),
	.a(n18876));
   in01f04 U19248 (.o(n18414),
	.a(n18423));
   ao22f04 U19249 (.o(n19315),
	.a(FE_OCPN25813_FE_OFN24735_n19306),
	.b(east_input_NIB_storage_data_f_1__35_),
	.c(n19400),
	.d(east_input_NIB_storage_data_f_3__35_));
   ao22f02 U19250 (.o(n18318),
	.a(proc_input_NIB_storage_data_f_7__41_),
	.b(n17779),
	.c(proc_input_NIB_storage_data_f_1__41_),
	.d(FE_OFN161_n24129));
   in01f10 U19251 (.o(n17751),
	.a(n18733));
   ao22f04 U19252 (.o(n18317),
	.a(proc_input_NIB_storage_data_f_5__41_),
	.b(FE_RN_49),
	.c(proc_input_NIB_storage_data_f_14__41_),
	.d(FE_OFN25644_n19504));
   in01f08 U19253 (.o(n25247),
	.a(n22912));
   ao22f04 U19254 (.o(n17902),
	.a(proc_input_NIB_storage_data_f_13__55_),
	.b(FE_OFN25602_n19530),
	.c(proc_input_NIB_storage_data_f_14__55_),
	.d(n19769));
   ao22f08 U19255 (.o(n17948),
	.a(proc_input_NIB_storage_data_f_13__54_),
	.b(FE_OFN25602_n19530),
	.c(proc_input_NIB_storage_data_f_0__54_),
	.d(FE_OCPN25933_n24342));
   ao22f04 U19256 (.o(n18483),
	.a(proc_input_NIB_storage_data_f_7__35_),
	.b(n17779),
	.c(proc_input_NIB_storage_data_f_1__35_),
	.d(FE_OFN161_n24129));
   ao22f04 U19258 (.o(n19558),
	.a(proc_input_NIB_storage_data_f_4__34_),
	.b(n17742),
	.c(proc_input_NIB_storage_data_f_13__34_),
	.d(FE_OFN25604_n19530));
   ao22f10 U19262 (.o(n17943),
	.a(FE_OFN25682_n17814),
	.b(proc_input_NIB_storage_data_f_9__54_),
	.c(proc_input_NIB_storage_data_f_10__54_),
	.d(FE_OCPN25957_n18039));
   na02f08 U19263 (.o(n17843),
	.a(n17845),
	.b(n17844));
   in01m06 U19264 (.o(n19719),
	.a(myLocX_f_3_));
   no02f06 U19265 (.o(n19873),
	.a(n19086),
	.b(n20759));
   no02f08 U19266 (.o(n19376),
	.a(FE_OFN25663_n19914),
	.b(n19373));
   no02f08 U19267 (.o(n19377),
	.a(FE_RN_57),
	.b(n24793));
   no02f06 U19268 (.o(n19384),
	.a(FE_OFN25663_n19914),
	.b(n19380));
   na02f06 U19269 (.o(n18488),
	.a(proc_input_NIB_storage_data_f_2__35_),
	.b(n24453));
   no02f06 U19270 (.o(n19385),
	.a(FE_RN_57),
	.b(n24767));
   na02f03 U19271 (.o(n18224),
	.a(proc_input_NIB_storage_data_f_1__36_),
	.b(FE_OFN161_n24129));
   na02f03 U19272 (.o(n17877),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__36_));
   in01f04 U19273 (.o(n18169),
	.a(n19084));
   ao22f20 U19274 (.o(n19345),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__51_),
	.c(FE_OCPN25813_FE_OFN24735_n19306),
	.d(east_input_NIB_storage_data_f_1__51_));
   no02f10 U19276 (.o(n19878),
	.a(myLocY_f_4_),
	.b(FE_OFN25624_n19003));
   na02f04 U19277 (.o(n17840),
	.a(n17977),
	.b(n17974));
   no02f06 U19278 (.o(n18438),
	.a(myLocY_f_1_),
	.b(n22836));
   no02f06 U19279 (.o(n18840),
	.a(n19328),
	.b(n18843));
   ao22f08 U19280 (.o(n17944),
	.a(n19707),
	.b(proc_input_NIB_storage_data_f_3__54_),
	.c(proc_input_NIB_storage_data_f_7__54_),
	.d(FE_OFN20_n17779));
   na02f04 U19281 (.o(n18371),
	.a(n18373),
	.b(n18372));
   in01f02 U19282 (.o(n19321),
	.a(myLocY_f_3_));
   ao22f08 U19283 (.o(n19515),
	.a(n24454),
	.b(proc_input_NIB_storage_data_f_13__40_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__40_));
   ao22f04 U19284 (.o(n18323),
	.a(proc_input_NIB_storage_data_f_0__41_),
	.b(FE_OCPN25933_n24342),
	.c(proc_input_NIB_storage_data_f_13__41_),
	.d(FE_OFN191_n24454));
   na02f04 U19285 (.o(n17980),
	.a(FE_RN_33),
	.b(proc_input_NIB_storage_data_f_3__50_));
   ao22f04 U19286 (.o(n18750),
	.a(n17782),
	.b(south_input_NIB_storage_data_f_2__31_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__31_));
   no02f03 U19287 (.o(n19314),
	.a(FE_OFN25664_n19914),
	.b(n19309));
   in01f03 U19288 (.o(n19518),
	.a(myLocY_f_7_));
   in01m02 U19289 (.o(n19241),
	.a(n19238));
   oa12f06 U19290 (.o(n19138),
	.a(n19076),
	.b(n19077),
	.c(n19225));
   na02f06 U19291 (.o(n17986),
	.a(proc_input_NIB_storage_data_f_10__50_),
	.b(FE_OCPN25964_n18039));
   na02f04 U19292 (.o(n17972),
	.a(FE_OCPN25962_n18039),
	.b(proc_input_NIB_storage_data_f_10__59_));
   na02f08 U19293 (.o(n18152),
	.a(proc_input_NIB_storage_data_f_10__56_),
	.b(FE_OCPN25959_n18039));
   ao22f04 U19294 (.o(n19516),
	.a(FE_OFN25679_n17814),
	.b(proc_input_NIB_storage_data_f_9__40_),
	.c(FE_OCPN25955_n18039),
	.d(proc_input_NIB_storage_data_f_10__40_));
   na02f04 U19295 (.o(n17904),
	.a(proc_input_NIB_storage_data_f_3__55_),
	.b(n19707));
   no02f03 U19296 (.o(n19139),
	.a(FE_OFN24776_n19073),
	.b(n19074));
   no02f02 U19297 (.o(n19140),
	.a(FE_OFN176_n24364),
	.b(n19072));
   na02f06 U19299 (.o(n18459),
	.a(n19155),
	.b(n19156));
   ao22f08 U19300 (.o(n17922),
	.a(proc_input_NIB_storage_data_f_14__37_),
	.b(FE_OFN25644_n19504),
	.c(proc_input_NIB_storage_data_f_12__37_),
	.d(n17747));
   ao22f08 U19301 (.o(n18491),
	.a(proc_input_NIB_storage_data_f_6__35_),
	.b(n19503),
	.c(proc_input_NIB_storage_data_f_12__35_),
	.d(n17777));
   ao22f08 U19302 (.o(n18490),
	.a(proc_input_NIB_storage_data_f_13__35_),
	.b(FE_OFN191_n24454),
	.c(proc_input_NIB_storage_data_f_0__35_),
	.d(FE_OCPN25933_n24342));
   no02f01 U19303 (.o(n17928),
	.a(n18036),
	.b(n17929));
   na02f20 U19304 (.o(n21162),
	.a(n18906),
	.b(n18905));
   no02f06 U19305 (.o(n19313),
	.a(FE_OFN24733_n19306),
	.b(n24893));
   no02f02 U19306 (.o(n19116),
	.a(FE_OFN176_n24364),
	.b(n19110));
   in01m08 U19307 (.o(n19701),
	.a(myLocX_f_5_));
   na02f04 U19308 (.o(n17960),
	.a(proc_input_NIB_storage_data_f_0__59_),
	.b(FE_OCPN25841_n24342));
   in01m10 U19309 (.o(n19633),
	.a(myChipID_f_5_));
   in01f04 U19311 (.o(n20123),
	.a(south_output_current_route_connection_0_));
   ao22f02 U19312 (.o(n19101),
	.a(FE_RN_11),
	.b(north_input_NIB_storage_data_f_2__32_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__32_));
   in01f06 U19313 (.o(n19720),
	.a(myLocX_f_4_));
   in01f04 U19314 (.o(n19706),
	.a(myLocX_f_2_));
   in01m03 U19315 (.o(n19326),
	.a(myLocY_f_1_));
   in01f02 U19316 (.o(n24895),
	.a(east_input_NIB_storage_data_f_1__43_));
   ao22f02 U19317 (.o(n19102),
	.a(FE_OFN51_n19193),
	.b(north_input_NIB_storage_data_f_3__32_),
	.c(FE_OFN24769_n19075),
	.d(north_input_NIB_storage_data_f_0__32_));
   ao22f06 U19318 (.o(n19662),
	.a(FE_OCPN25829_n21745),
	.b(proc_input_NIB_storage_data_f_2__53_),
	.c(FE_OCPN25947_n19595),
	.d(proc_input_NIB_storage_data_f_15__53_));
   no02f04 U19319 (.o(n19883),
	.a(myLocY_f_7_),
	.b(n22926));
   no02f10 U19320 (.o(n18150),
	.a(n20506),
	.b(n19339));
   ao22f04 U19321 (.o(n19554),
	.a(n17779),
	.b(proc_input_NIB_storage_data_f_7__34_),
	.c(FE_OFN188_n24453),
	.d(proc_input_NIB_storage_data_f_2__34_));
   ao22f06 U19322 (.o(n19551),
	.a(n19709),
	.b(proc_input_NIB_storage_data_f_3__34_),
	.c(FE_OFN169_n24343),
	.d(proc_input_NIB_storage_data_f_8__34_));
   no02m08 U19323 (.o(n19861),
	.a(south_output_current_route_connection_2_),
	.b(south_output_current_route_connection_1_));
   ao22f08 U19325 (.o(n19511),
	.a(FE_OCPN25918_n19547),
	.b(proc_input_NIB_storage_data_f_11__40_),
	.c(FE_OFN167_n24343),
	.d(proc_input_NIB_storage_data_f_8__40_));
   oa12f04 U19326 (.o(n19114),
	.a(n19112),
	.b(n19113),
	.c(n19225));
   ao22f03 U19327 (.o(n18751),
	.a(FE_OCPN25943_n24965),
	.b(south_input_NIB_storage_data_f_3__31_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__31_));
   no02f08 U19328 (.o(n19874),
	.a(myLocY_f_5_),
	.b(n19002));
   na02f03 U19329 (.o(n17966),
	.a(proc_input_NIB_storage_data_f_6__59_),
	.b(n19503));
   na02f04 U19330 (.o(n18165),
	.a(proc_input_NIB_storage_data_f_2__56_),
	.b(FE_RN_38));
   na02f03 U19331 (.o(n18418),
	.a(proc_input_NIB_storage_data_f_2__57_),
	.b(FE_OCPN25829_n21745));
   no02f02 U19332 (.o(n19115),
	.a(FE_OFN24776_n19073),
	.b(n19111));
   na02f08 U19333 (.o(n18737),
	.a(n18745),
	.b(n18743));
   ao22f04 U19334 (.o(n19265),
	.a(FE_OFN24777_n19932),
	.b(east_input_NIB_storage_data_f_0__44_),
	.c(FE_OFN24800_n20506),
	.d(east_input_NIB_storage_data_f_3__44_));
   na02f08 U19335 (.o(n20911),
	.a(n18706),
	.b(n18707));
   no02f04 U19336 (.o(n19001),
	.a(myLocY_f_6_),
	.b(n23184));
   ao22f04 U19337 (.o(n19517),
	.a(n19544),
	.b(proc_input_NIB_storage_data_f_15__40_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__40_));
   na02f06 U19338 (.o(n17969),
	.a(proc_input_NIB_storage_data_f_13__59_),
	.b(n24454));
   no02f02 U19339 (.o(n19109),
	.a(FE_OFN176_n24364),
	.b(n19103));
   no02f02 U19340 (.o(n19108),
	.a(FE_OFN24776_n19073),
	.b(n19104));
   no02m04 U19341 (.o(n24953),
	.a(south_output_current_route_connection_0_),
	.b(south_output_current_route_connection_1_));
   na02f02 U19342 (.o(n18322),
	.a(proc_input_NIB_storage_data_f_2__41_),
	.b(FE_OFN188_n24453));
   na02f02 U19343 (.o(n18315),
	.a(proc_input_NIB_storage_data_f_9__41_),
	.b(n19705));
   na02s04 U19344 (.o(n19454),
	.a(west_output_current_route_connection_1_),
	.b(west_output_current_route_connection_0_));
   no02f03 U19345 (.o(n17846),
	.a(n18036),
	.b(n17847));
   ao22f20 U19346 (.o(n19393),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__52_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__52_));
   in01f02 U19347 (.o(n17740),
	.a(proc_input_NIB_storage_data_f_9__53_));
   oa22f03 U19348 (.o(n19438),
	.a(FE_OFN25664_n19914),
	.b(n19433),
	.c(n20506),
	.d(n19432));
   oa22f04 U19349 (.o(n19437),
	.a(n21858),
	.b(n19436),
	.c(FE_OFN58_n19435),
	.d(n24891));
   oa22f04 U19350 (.o(n19431),
	.a(FE_OFN25664_n19914),
	.b(n19428),
	.c(n20506),
	.d(n19427));
   oa22f04 U19351 (.o(n19430),
	.a(n21858),
	.b(n19429),
	.c(n19933),
	.d(n24777));
   ao22f08 U19352 (.o(n19095),
	.a(FE_RN_11),
	.b(north_input_NIB_storage_data_f_2__36_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__36_));
   ao22f02 U19353 (.o(n18369),
	.a(proc_input_NIB_storage_data_f_8__43_),
	.b(FE_OFN169_n24343),
	.c(proc_input_NIB_storage_data_f_11__43_),
	.d(FE_OCPN25910_n19547));
   ao22f04 U19354 (.o(n19088),
	.a(FE_OFN51_n19193),
	.b(north_input_NIB_storage_data_f_3__38_),
	.c(FE_OFN24769_n19075),
	.d(north_input_NIB_storage_data_f_0__38_));
   oa22f04 U19356 (.o(n19420),
	.a(FE_OFN25664_n19914),
	.b(n19417),
	.c(n20506),
	.d(n19416));
   oa22f04 U19357 (.o(n19425),
	.a(n21858),
	.b(n19424),
	.c(FE_OFN61_n19435),
	.d(n24907));
   ao22f06 U19358 (.o(n17838),
	.a(FE_OFN169_n24343),
	.b(proc_input_NIB_storage_data_f_8__47_),
	.c(proc_input_NIB_storage_data_f_5__47_),
	.d(FE_RN_49));
   ao22f06 U19359 (.o(n17844),
	.a(FE_OCPN25933_n24342),
	.b(proc_input_NIB_storage_data_f_0__47_),
	.c(FE_OCPN25912_n19547),
	.d(proc_input_NIB_storage_data_f_11__47_));
   ao22f06 U19360 (.o(n19318),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__36_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__36_));
   ao22f04 U19361 (.o(n18516),
	.a(proc_input_NIB_storage_data_f_11__45_),
	.b(FE_OCPN25916_n19547),
	.c(proc_input_NIB_storage_data_f_5__45_),
	.d(FE_RN_49));
   ao22f04 U19362 (.o(n19092),
	.a(FE_RN_11),
	.b(north_input_NIB_storage_data_f_2__34_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__34_));
   oa22f04 U19364 (.o(n19426),
	.a(FE_OFN25664_n19914),
	.b(n19423),
	.c(n20506),
	.d(n19422));
   na02f20 U19365 (.o(n18581),
	.a(south_input_NIB_storage_data_f_1__62_),
	.b(n18061));
   ao22f02 U19367 (.o(n19695),
	.a(n19709),
	.b(proc_input_NIB_storage_data_f_3__46_),
	.c(FE_OFN156_n24129),
	.d(proc_input_NIB_storage_data_f_1__46_));
   ao22f02 U19368 (.o(n19691),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__46_),
	.c(FE_OFN25637_n19595),
	.d(proc_input_NIB_storage_data_f_15__46_));
   ao22f20 U19370 (.o(n18686),
	.a(n19973),
	.b(south_input_NIB_storage_data_f_2__50_),
	.c(n18061),
	.d(south_input_NIB_storage_data_f_1__50_));
   ao22f10 U19371 (.o(n18911),
	.a(FE_OFN24763_n18960),
	.b(west_input_NIB_storage_data_f_2__63_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__63_));
   na02f06 U19372 (.o(n18744),
	.a(FE_OCPN25941_n24965),
	.b(south_input_NIB_storage_data_f_3__44_));
   ao22f06 U19373 (.o(n19239),
	.a(FE_OFN24770_n19075),
	.b(north_input_NIB_storage_data_f_0__49_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__49_));
   oa22f04 U19374 (.o(n19419),
	.a(n21858),
	.b(n19418),
	.c(FE_OFN59_n19435),
	.d(n24905));
   na02f02 U19375 (.o(n19112),
	.a(FE_OFN24769_n19075),
	.b(north_input_NIB_storage_data_f_0__30_));
   ao22f04 U19376 (.o(n18007),
	.a(proc_input_NIB_storage_data_f_4__44_),
	.b(n17744),
	.c(proc_input_NIB_storage_data_f_8__44_),
	.d(FE_OFN167_n24343));
   ao22f04 U19377 (.o(n17975),
	.a(proc_input_NIB_storage_data_f_1__47_),
	.b(FE_OFN161_n24129),
	.c(proc_input_NIB_storage_data_f_4__47_),
	.d(n17742));
   ao22f04 U19378 (.o(n17836),
	.a(FE_OFN186_n24453),
	.b(proc_input_NIB_storage_data_f_2__47_),
	.c(n19705),
	.d(proc_input_NIB_storage_data_f_9__47_));
   ao22f02 U19379 (.o(n18961),
	.a(n18960),
	.b(west_input_NIB_storage_data_f_2__31_),
	.c(n18828),
	.d(west_input_NIB_storage_data_f_1__31_));
   in01f03 U19381 (.o(n18836),
	.a(n18835));
   ao22f08 U19382 (.o(n18746),
	.a(n17782),
	.b(south_input_NIB_storage_data_f_2__45_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__45_));
   ao22f06 U19383 (.o(n18004),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__44_),
	.c(proc_input_NIB_storage_data_f_12__44_),
	.d(FE_OCPN25969_n19500));
   oa22f04 U19384 (.o(n19226),
	.a(n19225),
	.b(n19224),
	.c(FE_OFN176_n24364),
	.d(n19222));
   oa22f04 U19385 (.o(n18800),
	.a(n24965),
	.b(n18799),
	.c(FE_OFN24745_n18648),
	.d(n18798));
   oa22f06 U19386 (.o(n18767),
	.a(n24965),
	.b(n18766),
	.c(FE_OFN24745_n18648),
	.d(n18765));
   in01f10 U19387 (.o(n19347),
	.a(myChipID_f_12_));
   oa22f04 U19388 (.o(n19227),
	.a(n19159),
	.b(n19221),
	.c(FE_OFN24776_n19073),
	.d(n19219));
   in01f10 U19389 (.o(n19584),
	.a(myChipID_f_11_));
   ao22f04 U19390 (.o(n19704),
	.a(FE_OCPN25835_n24342),
	.b(proc_input_NIB_storage_data_f_0__44_),
	.c(FE_OCPN25917_n19547),
	.d(proc_input_NIB_storage_data_f_11__44_));
   in01f10 U19391 (.o(n18669),
	.a(n18663));
   in01f06 U19392 (.o(n18801),
	.a(n18797));
   in01f04 U19393 (.o(n19328),
	.a(myLocX_f_0_));
   ao22f04 U19394 (.o(n17845),
	.a(FE_OFN25604_n19530),
	.b(proc_input_NIB_storage_data_f_13__47_),
	.c(FE_OFN25685_n19500),
	.d(proc_input_NIB_storage_data_f_12__47_));
   ao22f04 U19396 (.o(n19087),
	.a(FE_RN_11),
	.b(north_input_NIB_storage_data_f_2__38_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__38_));
   ao22f06 U19397 (.o(n18747),
	.a(FE_OCPN25941_n24965),
	.b(south_input_NIB_storage_data_f_3__45_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__45_));
   ao22f06 U19398 (.o(n19096),
	.a(FE_OFN51_n19193),
	.b(north_input_NIB_storage_data_f_3__36_),
	.c(FE_OFN24769_n19075),
	.d(north_input_NIB_storage_data_f_0__36_));
   ao22f02 U19399 (.o(n19690),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__46_),
	.c(n17779),
	.d(proc_input_NIB_storage_data_f_7__46_));
   ao22f08 U19401 (.o(n19274),
	.a(FE_OFN24777_n19932),
	.b(east_input_NIB_storage_data_f_0__46_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__46_));
   ao22f04 U19402 (.o(n18362),
	.a(proc_input_NIB_storage_data_f_12__43_),
	.b(FE_OFN25686_n19500),
	.c(proc_input_NIB_storage_data_f_14__43_),
	.d(n19769));
   in01f80 U19404 (.o(n19657),
	.a(myChipID_f_0_));
   in01f03 U19405 (.o(n19132),
	.a(myLocY_f_4_));
   no02f08 U19406 (.o(n18854),
	.a(n18997),
	.b(n18850));
   no02f08 U19407 (.o(n18855),
	.a(n18995),
	.b(n18849));
   no02f20 U19408 (.o(n18933),
	.a(FE_OCPN25925_n18828),
	.b(n18929));
   no02f20 U19409 (.o(n18897),
	.a(FE_RN_7),
	.b(n18894));
   no02f20 U19410 (.o(n18926),
	.a(n18995),
	.b(n18921));
   ao22f04 U19411 (.o(n18357),
	.a(proc_input_NIB_storage_data_f_2__44_),
	.b(FE_RN_38),
	.c(proc_input_NIB_storage_data_f_10__44_),
	.d(FE_OCPN25956_n18039));
   ao22f04 U19412 (.o(n18006),
	.a(FE_OFN25634_n19595),
	.b(proc_input_NIB_storage_data_f_15__44_),
	.c(n19769),
	.d(proc_input_NIB_storage_data_f_14__44_));
   no02f10 U19413 (.o(n18659),
	.a(n18754),
	.b(n18143));
   na02f04 U19414 (.o(n18356),
	.a(proc_input_NIB_storage_data_f_9__44_),
	.b(FE_OFN25677_n17814));
   ao22f02 U19415 (.o(n18509),
	.a(proc_input_NIB_storage_data_f_1__45_),
	.b(FE_OFN161_n24129),
	.c(proc_input_NIB_storage_data_f_9__45_),
	.d(n19705));
   na02f03 U19416 (.o(n17974),
	.a(proc_input_NIB_storage_data_f_6__47_),
	.b(n19503));
   ao22f10 U19417 (.o(n18940),
	.a(FE_RN_64),
	.b(west_input_NIB_storage_data_f_3__56_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__56_));
   in01f06 U19418 (.o(n18785),
	.a(n18779));
   na02f08 U19419 (.o(n18460),
	.a(n19156),
	.b(myChipID_f_8_));
   na02f08 U19420 (.o(n18748),
	.a(n18740),
	.b(n18739));
   ao22f04 U19421 (.o(n18366),
	.a(proc_input_NIB_storage_data_f_3__43_),
	.b(n21768),
	.c(proc_input_NIB_storage_data_f_4__43_),
	.d(n17743));
   oa22f04 U19422 (.o(n18759),
	.a(n24965),
	.b(n18758),
	.c(FE_OFN24745_n18648),
	.d(n18757));
   oa22f03 U19423 (.o(n18783),
	.a(n24965),
	.b(n18782),
	.c(FE_OFN24745_n18648),
	.d(n18781));
   in01f06 U19424 (.o(n24989),
	.a(south_output_current_route_connection_1_));
   ao22f03 U19425 (.o(n19696),
	.a(proc_input_NIB_storage_data_f_11__46_),
	.b(n24455),
	.c(proc_input_NIB_storage_data_f_0__46_),
	.d(FE_OCPN25933_n24342));
   ao22f20 U19426 (.o(n18652),
	.a(n19973),
	.b(south_input_NIB_storage_data_f_2__59_),
	.c(n17756),
	.d(south_input_NIB_storage_data_f_1__59_));
   in01m02 U19427 (.o(n24767),
	.a(east_input_NIB_storage_data_f_1__60_));
   no02f04 U19428 (.o(n18875),
	.a(n18995),
	.b(n18863));
   no02f04 U19429 (.o(n18876),
	.a(FE_OCPN25927_n18828),
	.b(n18864));
   no02f06 U19430 (.o(n18862),
	.a(n18995),
	.b(n18856));
   no02f04 U19431 (.o(n19273),
	.a(FE_OFN25664_n19914),
	.b(n19268));
   no02f06 U19432 (.o(n18861),
	.a(FE_OFN183_n24390),
	.b(n18857));
   no02f03 U19433 (.o(n19272),
	.a(FE_RN_57),
	.b(n24911));
   oa12f03 U19434 (.o(n18956),
	.a(n18954),
	.b(n18955),
	.c(n24465));
   ao22f10 U19435 (.o(n19264),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__45_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__45_));
   ao22f06 U19436 (.o(n19718),
	.a(FE_OCPN25967_n19500),
	.b(proc_input_NIB_storage_data_f_12__45_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__45_));
   in01f02 U19437 (.o(n19111),
	.a(north_input_NIB_storage_data_f_2__30_));
   in01f02 U19439 (.o(n19455),
	.a(north_input_valid));
   in01f04 U19441 (.o(n24765),
	.a(east_input_NIB_storage_data_f_1__62_));
   in01m03 U19442 (.o(n24793),
	.a(east_input_NIB_storage_data_f_1__53_));
   in01m03 U19443 (.o(n24785),
	.a(east_input_NIB_storage_data_f_1__57_));
   ao22f06 U19445 (.o(n19263),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__45_),
	.c(FE_OFN24800_n20506),
	.d(east_input_NIB_storage_data_f_3__45_));
   ao22f04 U19446 (.o(n17835),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__47_),
	.c(FE_OFN25632_n19595),
	.d(proc_input_NIB_storage_data_f_15__47_));
   ao22f04 U19447 (.o(n17887),
	.a(north_input_NIB_storage_data_f_2__46_),
	.b(FE_RN_11),
	.c(north_input_NIB_storage_data_f_0__46_),
	.d(FE_OFN24770_n19075));
   ao22f04 U19448 (.o(n18373),
	.a(proc_input_NIB_storage_data_f_6__43_),
	.b(n19503),
	.c(proc_input_NIB_storage_data_f_9__43_),
	.d(n19705));
   in01f06 U19449 (.o(n19708),
	.a(myLocX_f_1_));
   ao22m02 U19451 (.o(n18962),
	.a(FE_RN_5),
	.b(west_input_NIB_storage_data_f_3__31_),
	.c(FE_OFN27_n18974),
	.d(west_input_NIB_storage_data_f_0__31_));
   no02f03 U19452 (.o(n18565),
	.a(FE_OFN24806_n19655),
	.b(n18566));
   na02f04 U19453 (.o(n17886),
	.a(north_input_NIB_storage_data_f_3__46_),
	.b(FE_OFN51_n19193));
   no02f10 U19454 (.o(n19352),
	.a(FE_OFN25663_n19914),
	.b(n19348));
   no02f10 U19455 (.o(n19353),
	.a(FE_RN_57),
	.b(n24783));
   ao22f04 U19456 (.o(n18510),
	.a(proc_input_NIB_storage_data_f_7__45_),
	.b(FE_OFN20_n17779),
	.c(proc_input_NIB_storage_data_f_3__45_),
	.d(n21768));
   in01f04 U19457 (.o(n18461),
	.a(n19155));
   na02f10 U19458 (.o(n18000),
	.a(proc_input_NIB_storage_data_f_13__44_),
	.b(n24454));
   na02f06 U19459 (.o(n18355),
	.a(proc_input_NIB_storage_data_f_1__44_),
	.b(FE_OFN161_n24129));
   na02f08 U19460 (.o(n18183),
	.a(n18960),
	.b(west_input_NIB_storage_data_f_2__55_));
   in01m02 U19461 (.o(n19373),
	.a(east_input_NIB_storage_data_f_2__53_));
   in01f03 U19462 (.o(n19337),
	.a(east_input_NIB_storage_data_f_2__62_));
   in01f03 U19463 (.o(n19366),
	.a(east_input_NIB_storage_data_f_2__57_));
   in01m02 U19464 (.o(n19380),
	.a(east_input_NIB_storage_data_f_2__60_));
   in01m02 U19465 (.o(n19339),
	.a(east_input_NIB_storage_data_f_3__62_));
   na02f02 U19466 (.o(n17976),
	.a(proc_input_NIB_storage_data_f_3__47_),
	.b(n21768));
   ao22f10 U19467 (.o(n18915),
	.a(FE_OFN24763_n18960),
	.b(west_input_NIB_storage_data_f_2__62_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__62_));
   ao22f04 U19468 (.o(n19093),
	.a(FE_OFN51_n19193),
	.b(north_input_NIB_storage_data_f_3__34_),
	.c(FE_OFN24769_n19075),
	.d(north_input_NIB_storage_data_f_0__34_));
   no02f08 U19469 (.o(n17804),
	.a(myLocX_f_6_),
	.b(n22858));
   na02f04 U19470 (.o(n18361),
	.a(proc_input_NIB_storage_data_f_7__43_),
	.b(FE_OFN20_n17779));
   na02f03 U19471 (.o(n17885),
	.a(north_input_NIB_storage_data_f_1__46_),
	.b(n24364));
   in01f02 U19472 (.o(n19086),
	.a(myLocY_f_5_));
   in01f03 U19473 (.o(n19368),
	.a(east_input_NIB_storage_data_f_3__57_));
   na02f04 U19474 (.o(n18519),
	.a(proc_input_NIB_storage_data_f_2__45_),
	.b(FE_OCPN25823_n21745));
   no02m02 U19475 (.o(n18295),
	.a(n18706),
	.b(myLocY_f_1_));
   ao22f08 U19476 (.o(n18753),
	.a(n24472),
	.b(south_input_NIB_storage_data_f_0__46_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__46_));
   na02f10 U19477 (.o(n22912),
	.a(south_input_valid),
	.b(n20590));
   ao22f02 U19478 (.o(n19689),
	.a(n17747),
	.b(proc_input_NIB_storage_data_f_12__46_),
	.c(FE_OFN25604_n19530),
	.d(proc_input_NIB_storage_data_f_13__46_));
   in01f02 U19479 (.o(n19100),
	.a(north_input_control_header_last_f));
   ao22f02 U19480 (.o(n19698),
	.a(n24343),
	.b(proc_input_NIB_storage_data_f_8__46_),
	.c(n17742),
	.d(proc_input_NIB_storage_data_f_4__46_));
   in01f03 U19481 (.o(n19081),
	.a(north_input_NIB_storage_data_f_3__40_));
   ao22f06 U19482 (.o(n18712),
	.a(FE_OCPN25939_n24965),
	.b(south_input_NIB_storage_data_f_3__34_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__34_));
   in01f02 U19483 (.o(n24893),
	.a(east_input_NIB_storage_data_f_1__34_));
   na02f04 U19484 (.o(n17997),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__44_));
   in01f02 U19487 (.o(n19311),
	.a(east_input_NIB_storage_data_f_3__34_));
   no02f02 U19488 (.o(n18958),
	.a(n18995),
	.b(n18952));
   no02m02 U19489 (.o(n18957),
	.a(FE_OFN24748_n18828),
	.b(n18953));
   na02f02 U19490 (.o(n18372),
	.a(proc_input_NIB_storage_data_f_2__43_),
	.b(FE_OFN188_n24453));
   no02f02 U19491 (.o(n18298),
	.a(n18707),
	.b(myLocY_f_1_));
   na02f04 U19492 (.o(n18365),
	.a(proc_input_NIB_storage_data_f_10__43_),
	.b(n18034));
   na02m06 U19493 (.o(n19099),
	.a(north_input_control_thanks_all_f),
	.b(north_input_control_count_zero_f));
   ao22f08 U19494 (.o(n18707),
	.a(FE_OCPN25943_n24965),
	.b(south_input_NIB_storage_data_f_3__35_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__35_));
   oa22f04 U19495 (.o(n18973),
	.a(FE_OFN30_n18974),
	.b(n18969),
	.c(FE_RN_7),
	.d(n18968));
   oa22f04 U19496 (.o(n18972),
	.a(n24465),
	.b(n18971),
	.c(n18995),
	.d(n18970));
   ao22f04 U19497 (.o(n19205),
	.a(FE_OFN51_n19193),
	.b(north_input_NIB_storage_data_f_3__42_),
	.c(FE_OFN24770_n19075),
	.d(north_input_NIB_storage_data_f_0__42_));
   ao22f08 U19498 (.o(n18742),
	.a(n24472),
	.b(south_input_NIB_storage_data_f_0__43_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__43_));
   no02f10 U19499 (.o(n18993),
	.a(n18997),
	.b(n18990));
   no02f06 U19500 (.o(n18983),
	.a(n18995),
	.b(n18977));
   ao22f06 U19501 (.o(n19212),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__45_),
	.c(FE_OFN24770_n19075),
	.d(north_input_NIB_storage_data_f_0__45_));
   no02f06 U19502 (.o(n18982),
	.a(FE_OCPN25925_n18828),
	.b(n18978));
   ao22f08 U19503 (.o(n18703),
	.a(FE_OCPN25943_n24965),
	.b(south_input_NIB_storage_data_f_3__37_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__37_));
   no02f10 U19505 (.o(n18333),
	.a(n18334),
	.b(FE_OFN24745_n18648));
   na02m04 U19506 (.o(n18780),
	.a(FE_OFN24741_n18683),
	.b(south_input_NIB_storage_data_f_1__32_));
   no02f10 U19507 (.o(n18790),
	.a(proc_output_current_route_connection_1_),
	.b(proc_output_current_route_connection_0_));
   ao22f08 U19508 (.o(n19177),
	.a(FE_RN_10),
	.b(north_input_NIB_storage_data_f_3__62_),
	.c(FE_OFN24773_n19075),
	.d(north_input_NIB_storage_data_f_0__62_));
   na02f03 U19509 (.o(n18954),
	.a(FE_OFN27_n18974),
	.b(west_input_NIB_storage_data_f_0__32_));
   oa22f02 U19510 (.o(n19217),
	.a(n19225),
	.b(n19216),
	.c(FE_OFN176_n24364),
	.d(n19215));
   oa22f10 U19511 (.o(n18728),
	.a(n24965),
	.b(n18727),
	.c(n24964),
	.d(n18726));
   ao22f08 U19512 (.o(n18706),
	.a(n21365),
	.b(south_input_NIB_storage_data_f_2__35_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__35_));
   oa22f04 U19513 (.o(n19218),
	.a(FE_OFN264_n25427),
	.b(n19214),
	.c(FE_OFN24776_n19073),
	.d(n19213));
   in01f10 U19514 (.o(n19622),
	.a(myChipID_f_9_));
   in01f10 U19515 (.o(n18729),
	.a(n18725));
   in01f10 U19516 (.o(n18723),
	.a(n18719));
   in01f10 U19517 (.o(n18085),
	.a(n18998));
   ao22f06 U19518 (.o(n18976),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__36_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__36_));
   in01f04 U19519 (.o(n18347),
	.a(n18348));
   in01m10 U19520 (.o(south_input_valid),
	.a(n19452));
   ao22f08 U19521 (.o(n18709),
	.a(n24165),
	.b(south_input_NIB_storage_data_f_2__38_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__38_));
   oa22f03 U19522 (.o(n18832),
	.a(west_input_NIB_head_ptr_f_1_),
	.b(n18819),
	.c(n18818),
	.d(FE_OCPN25820_west_input_NIB_head_ptr_f_1));
   ao22f08 U19523 (.o(n18741),
	.a(FE_OCPN25941_n24965),
	.b(south_input_NIB_storage_data_f_3__43_),
	.c(n24165),
	.d(south_input_NIB_storage_data_f_2__43_));
   no02f10 U19524 (.o(n19000),
	.a(n24390),
	.b(n18996));
   no02f10 U19525 (.o(n18086),
	.a(n18995),
	.b(n18994));
   no02f08 U19526 (.o(n18087),
	.a(n24465),
	.b(n18999));
   in01m04 U19527 (.o(n24783),
	.a(east_input_NIB_storage_data_f_1__54_));
   na02f06 U19528 (.o(n18763),
	.a(FE_OFN25648_n18762),
	.b(south_input_NIB_storage_data_f_2__48_));
   na03f10 U19530 (.o(n18252),
	.a(n19154),
	.b(n19153),
	.c(n19647));
   ao22f20 U19531 (.o(n19175),
	.a(FE_OFN96_n21865),
	.b(north_input_NIB_storage_data_f_2__61_),
	.c(FE_OFN25610_n19071),
	.d(north_input_NIB_storage_data_f_1__61_));
   in01m03 U19532 (.o(n24907),
	.a(east_input_NIB_storage_data_f_1__39_));
   no04f10 U19533 (.o(n18804),
	.a(myLocX_f_0_),
	.b(myLocX_f_7_),
	.c(myLocX_f_5_),
	.d(myLocX_f_6_));
   no04f10 U19534 (.o(n18805),
	.a(myLocX_f_1_),
	.b(myLocX_f_2_),
	.c(myLocX_f_3_),
	.d(myLocX_f_4_));
   in01f02 U19535 (.o(n18856),
	.a(west_input_NIB_storage_data_f_2__49_));
   in01f02 U19536 (.o(n18921),
	.a(west_input_NIB_storage_data_f_2__61_));
   in01m02 U19537 (.o(n18781),
	.a(south_input_NIB_storage_data_f_0__32_));
   in01f03 U19538 (.o(n18666),
	.a(south_input_NIB_storage_data_f_3__55_));
   in01f03 U19539 (.o(n18655),
	.a(south_input_NIB_storage_data_f_0__58_));
   in01f04 U19540 (.o(n19348),
	.a(east_input_NIB_storage_data_f_2__54_));
   in01f03 U19541 (.o(n18852),
	.a(west_input_NIB_storage_data_f_3__48_));
   in01f04 U19542 (.o(n18126),
	.a(west_input_NIB_storage_data_f_0__54_));
   in01f04 U19543 (.o(n18895),
	.a(west_input_NIB_storage_data_f_3__54_));
   ao22f06 U19544 (.o(n19210),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__44_),
	.c(FE_OFN24770_n19075),
	.d(north_input_NIB_storage_data_f_0__44_));
   ao22f20 U19545 (.o(n18619),
	.a(south_input_NIB_storage_data_f_1__39_),
	.b(FE_OFN24742_n18683),
	.c(south_input_NIB_storage_data_f_3__39_),
	.d(FE_OCPN25944_n24965));
   in01f02 U19546 (.o(n24911),
	.a(east_input_NIB_storage_data_f_1__42_));
   na02f08 U19547 (.o(n18764),
	.a(FE_OFN24741_n18683),
	.b(south_input_NIB_storage_data_f_1__48_));
   in01m06 U19548 (.o(n25061),
	.a(proc_output_current_route_connection_2_));
   in01m06 U19549 (.o(n18931),
	.a(west_input_NIB_storage_data_f_3__50_));
   oa22f08 U19550 (.o(n18722),
	.a(n24965),
	.b(n18721),
	.c(FE_OFN24745_n18648),
	.d(n18720));
   na02f06 U19551 (.o(n18756),
	.a(FE_OFN24742_n18683),
	.b(south_input_NIB_storage_data_f_1__49_));
   in01m03 U19552 (.o(n24777),
	.a(east_input_NIB_storage_data_f_1__41_));
   in01m03 U19553 (.o(n24891),
	.a(east_input_NIB_storage_data_f_1__40_));
   na02f10 U19555 (.o(n18663),
	.a(FE_RN_41),
	.b(south_input_NIB_storage_data_f_2__55_));
   ao12f06 U19556 (.o(n18740),
	.a(n18341),
	.b(FE_OCPN25941_n24965),
	.c(south_input_NIB_storage_data_f_3__42_));
   na02f10 U19557 (.o(n18617),
	.a(south_input_NIB_storage_data_f_0__39_),
	.b(n24472));
   in01m02 U19558 (.o(n19268),
	.a(east_input_NIB_storage_data_f_2__42_));
   in01f02 U19559 (.o(n18864),
	.a(west_input_NIB_storage_data_f_1__46_));
   in01f03 U19560 (.o(n18928),
	.a(west_input_NIB_storage_data_f_2__50_));
   in01m02 U19561 (.o(n18929),
	.a(west_input_NIB_storage_data_f_1__50_));
   in01m02 U19562 (.o(n18894),
	.a(west_input_NIB_storage_data_f_1__54_));
   in01f02 U19563 (.o(n18863),
	.a(west_input_NIB_storage_data_f_2__46_));
   in01m02 U19564 (.o(n18849),
	.a(west_input_NIB_storage_data_f_2__48_));
   in01m02 U19565 (.o(n18850),
	.a(west_input_NIB_storage_data_f_1__48_));
   in01f02 U19566 (.o(n18857),
	.a(west_input_NIB_storage_data_f_1__49_));
   in01m02 U19567 (.o(n18782),
	.a(south_input_NIB_storage_data_f_3__32_));
   in01m02 U19568 (.o(n18757),
	.a(south_input_NIB_storage_data_f_0__49_));
   in01m02 U19569 (.o(n18758),
	.a(south_input_NIB_storage_data_f_3__49_));
   in01m02 U19570 (.o(n19219),
	.a(north_input_NIB_storage_data_f_2__48_));
   in01m02 U19571 (.o(n19427),
	.a(east_input_NIB_storage_data_f_3__41_));
   in01m02 U19572 (.o(n19428),
	.a(east_input_NIB_storage_data_f_2__41_));
   in01m02 U19573 (.o(n19422),
	.a(east_input_NIB_storage_data_f_3__39_));
   in01m02 U19574 (.o(n19423),
	.a(east_input_NIB_storage_data_f_2__39_));
   in01m02 U19575 (.o(n19432),
	.a(east_input_NIB_storage_data_f_3__40_));
   in01m02 U19576 (.o(n19433),
	.a(east_input_NIB_storage_data_f_2__40_));
   in01f03 U19577 (.o(n18125),
	.a(west_input_NIB_storage_data_f_0__61_));
   in01f03 U19578 (.o(n18923),
	.a(west_input_NIB_storage_data_f_3__61_));
   in01f03 U19579 (.o(n18665),
	.a(south_input_NIB_storage_data_f_0__55_));
   in01f03 U19580 (.o(n18656),
	.a(south_input_NIB_storage_data_f_3__58_));
   in01m02 U19581 (.o(n18798),
	.a(south_input_NIB_storage_data_f_0__30_));
   in01m02 U19582 (.o(n18799),
	.a(south_input_NIB_storage_data_f_3__30_));
   in01m02 U19583 (.o(n18765),
	.a(south_input_NIB_storage_data_f_0__48_));
   in01m02 U19584 (.o(n18766),
	.a(south_input_NIB_storage_data_f_3__48_));
   in01m02 U19585 (.o(n19222),
	.a(north_input_NIB_storage_data_f_1__48_));
   in01m02 U19586 (.o(n19224),
	.a(north_input_NIB_storage_data_f_3__48_));
   in01m02 U19587 (.o(n18955),
	.a(west_input_NIB_storage_data_f_3__32_));
   in01f03 U19588 (.o(n18859),
	.a(west_input_NIB_storage_data_f_3__49_));
   in01f03 U19589 (.o(n18866),
	.a(west_input_NIB_storage_data_f_3__46_));
   na02f10 U19590 (.o(n18755),
	.a(FE_RN_17),
	.b(south_input_NIB_storage_data_f_2__49_));
   in01f03 U19591 (.o(n19350),
	.a(east_input_NIB_storage_data_f_3__54_));
   na02f10 U19592 (.o(east_input_valid),
	.a(n18787),
	.b(n25315));
   in01m02 U19593 (.o(n19221),
	.a(north_input_NIB_storage_data_f_0__48_));
   in01m02 U19594 (.o(n19424),
	.a(east_input_NIB_storage_data_f_0__39_));
   in01m02 U19595 (.o(n19429),
	.a(east_input_NIB_storage_data_f_0__41_));
   in01m02 U19596 (.o(n19436),
	.a(east_input_NIB_storage_data_f_0__40_));
   in01f02 U19597 (.o(n18953),
	.a(west_input_NIB_storage_data_f_1__32_));
   in01f02 U19599 (.o(n18922),
	.a(west_input_NIB_storage_data_f_1__61_));
   ao22f06 U19600 (.o(n19206),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__43_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__43_));
   ao22f08 U19601 (.o(n19209),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__44_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__44_));
   in01f02 U19602 (.o(n19416),
	.a(east_input_NIB_storage_data_f_3__38_));
   in01f02 U19603 (.o(n19417),
	.a(east_input_NIB_storage_data_f_2__38_));
   in01f02 U19604 (.o(n19418),
	.a(east_input_NIB_storage_data_f_0__38_));
   in01f02 U19606 (.o(n19270),
	.a(east_input_NIB_storage_data_f_3__42_));
   no02f02 U19607 (.o(n18349),
	.a(n18762),
	.b(n18350));
   na02f10 U19608 (.o(north_input_valid),
	.a(n18786),
	.b(n25288));
   no04f10 U19609 (.o(n18808),
	.a(myLocY_f_7_),
	.b(myLocY_f_6_),
	.c(myLocY_f_5_),
	.d(myLocY_f_4_));
   no04f10 U19610 (.o(n18809),
	.a(myLocY_f_1_),
	.b(myLocY_f_0_),
	.c(myLocY_f_2_),
	.d(myLocY_f_3_));
   no03f20 U19611 (.o(n19453),
	.a(west_input_NIB_elements_in_array_f_2_),
	.b(west_input_NIB_elements_in_array_f_1_),
	.c(west_input_NIB_elements_in_array_f_0_));
   na02f10 U19612 (.o(n18998),
	.a(FE_OFN27_n18974),
	.b(west_input_NIB_storage_data_f_0__41_));
   na02f06 U19613 (.o(n18772),
	.a(FE_OCPN25941_n24965),
	.b(south_input_NIB_storage_data_f_3__47_));
   na02f06 U19614 (.o(n18773),
	.a(FE_OFN24742_n18683),
	.b(south_input_NIB_storage_data_f_1__47_));
   no02f06 U19616 (.o(n18341),
	.a(FE_OFN24745_n18648),
	.b(n18342));
   na02f08 U19617 (.o(n18991),
	.a(n18127),
	.b(west_input_NIB_storage_data_f_0__40_));
   in01f10 U19618 (.o(n24165),
	.a(n18754));
   in01f04 U19620 (.o(n18771),
	.a(n18331));
   na02f20 U19621 (.o(n18794),
	.a(south_input_control_thanks_all_f),
	.b(south_input_control_count_zero_f));
   in01m02 U19622 (.o(n18334),
	.a(south_input_NIB_storage_data_f_0__54_));
   in01m10 U19623 (.o(n25422),
	.a(proc_output_current_route_connection_0_));
   in01m08 U19624 (.o(n25315),
	.a(east_input_NIB_elements_in_array_f_0_));
   ao22f08 U19625 (.o(n18986),
	.a(FE_OFN24764_n18960),
	.b(west_input_NIB_storage_data_f_2__38_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__38_));
   in01s10 U19626 (.o(n18795),
	.a(south_input_control_header_last_f));
   no02f02 U19627 (.o(n18818),
	.a(west_input_NIB_head_ptr_f_0_),
	.b(n18817));
   in01m02 U19628 (.o(n18822),
	.a(west_input_NIB_storage_data_f_2__45_));
   in01m02 U19629 (.o(n18989),
	.a(west_input_NIB_storage_data_f_2__40_));
   ao22f06 U19630 (.o(n18985),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__39_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__39_));
   no02m20 U19631 (.o(n18786),
	.a(north_input_NIB_elements_in_array_f_0_),
	.b(north_input_NIB_elements_in_array_f_2_));
   in01m02 U19632 (.o(n19216),
	.a(north_input_NIB_storage_data_f_3__47_));
   in01m02 U19633 (.o(n18820),
	.a(west_input_NIB_storage_data_f_3__45_));
   in01m02 U19634 (.o(n18823),
	.a(west_input_NIB_storage_data_f_0__45_));
   na02f06 U19635 (.o(n18348),
	.a(south_input_NIB_storage_data_f_3__46_),
	.b(FE_OCPN25939_n24965));
   in01f04 U19636 (.o(n18980),
	.a(west_input_NIB_storage_data_f_3__37_));
   in01m10 U19637 (.o(n25288),
	.a(north_input_NIB_elements_in_array_f_1_));
   no02m10 U19638 (.o(n18791),
	.a(proc_input_NIB_elements_in_array_f_2_),
	.b(proc_input_NIB_elements_in_array_f_3_));
   in01m02 U19639 (.o(n18994),
	.a(west_input_NIB_storage_data_f_2__41_));
   in01m02 U19640 (.o(n18999),
	.a(west_input_NIB_storage_data_f_3__41_));
   in01m02 U19641 (.o(n18996),
	.a(west_input_NIB_storage_data_f_1__41_));
   in01f03 U19642 (.o(n18992),
	.a(west_input_NIB_storage_data_f_3__40_));
   in01m02 U19643 (.o(n18990),
	.a(west_input_NIB_storage_data_f_1__40_));
   in01m02 U19644 (.o(n18977),
	.a(west_input_NIB_storage_data_f_2__37_));
   in01m02 U19645 (.o(n18978),
	.a(west_input_NIB_storage_data_f_1__37_));
   in01m02 U19646 (.o(n18971),
	.a(west_input_NIB_storage_data_f_3__35_));
   in01m02 U19647 (.o(n18970),
	.a(west_input_NIB_storage_data_f_2__35_));
   in01m02 U19648 (.o(n19213),
	.a(north_input_NIB_storage_data_f_2__47_));
   in01m02 U19649 (.o(n18968),
	.a(west_input_NIB_storage_data_f_1__35_));
   in01f03 U19650 (.o(n18839),
	.a(west_input_NIB_storage_data_f_3__42_));
   in01f03 U19651 (.o(n18838),
	.a(west_input_NIB_storage_data_f_1__42_));
   in01m02 U19652 (.o(n18726),
	.a(south_input_NIB_storage_data_f_0__40_));
   in01m02 U19653 (.o(n18727),
	.a(south_input_NIB_storage_data_f_3__40_));
   in01m02 U19654 (.o(n18720),
	.a(south_input_NIB_storage_data_f_0__41_));
   in01m02 U19655 (.o(n18721),
	.a(south_input_NIB_storage_data_f_3__41_));
   in01m02 U19656 (.o(n19215),
	.a(north_input_NIB_storage_data_f_1__47_));
   in01m02 U19657 (.o(n18821),
	.a(west_input_NIB_storage_data_f_1__45_));
   in01m02 U19658 (.o(n18969),
	.a(west_input_NIB_storage_data_f_0__35_));
   in01m02 U19659 (.o(n19214),
	.a(north_input_NIB_storage_data_f_0__47_));
   no02m10 U19660 (.o(n18787),
	.a(east_input_NIB_elements_in_array_f_1_),
	.b(east_input_NIB_elements_in_array_f_2_));
   in01f02 U19661 (.o(n18350),
	.a(south_input_NIB_storage_data_f_2__46_));
   no03f20 U19662 (.o(n19452),
	.a(south_input_NIB_elements_in_array_f_2_),
	.b(south_input_NIB_elements_in_array_f_0_),
	.c(south_input_NIB_elements_in_array_f_1_));
   na02f10 U19664 (.o(n18770),
	.a(n19973),
	.b(south_input_NIB_storage_data_f_2__47_));
   no02m10 U19665 (.o(n25475),
	.a(proc_input_NIB_elements_in_array_f_1_),
	.b(proc_input_NIB_elements_in_array_f_0_));
   no02f06 U19667 (.o(n18331),
	.a(FE_OFN24745_n18648),
	.b(n18332));
   in01f04 U19668 (.o(n19161),
	.a(north_input_NIB_storage_data_f_3__50_));
   in01f04 U19669 (.o(n24919),
	.a(east_input_NIB_storage_data_f_1__49_));
   in01f04 U19670 (.o(n24909),
	.a(east_input_NIB_storage_data_f_1__48_));
   in01f03 U19671 (.o(n18344),
	.a(south_input_NIB_storage_data_f_0__38_));
   in01m02 U19672 (.o(n18342),
	.a(south_input_NIB_storage_data_f_0__42_));
   in01f03 U19673 (.o(n19158),
	.a(north_input_NIB_storage_data_f_1__50_));
   in01f03 U19674 (.o(n19157),
	.a(north_input_NIB_storage_data_f_2__50_));
   in01f04 U19675 (.o(n19289),
	.a(east_input_NIB_storage_data_f_3__48_));
   in01m02 U19676 (.o(n19290),
	.a(east_input_NIB_storage_data_f_2__48_));
   in01m02 U19677 (.o(n19284),
	.a(east_input_NIB_storage_data_f_3__49_));
   in01m02 U19678 (.o(n19285),
	.a(east_input_NIB_storage_data_f_2__49_));
   in01f02 U19679 (.o(n18817),
	.a(west_input_NIB_storage_data_f_2__44_));
   in01f03 U19680 (.o(n19286),
	.a(east_input_NIB_storage_data_f_0__49_));
   in01f03 U19681 (.o(n19291),
	.a(east_input_NIB_storage_data_f_0__48_));
   in01f02 U19682 (.o(n18332),
	.a(south_input_NIB_storage_data_f_0__47_));
   no02f06 U19683 (.o(n20177),
	.a(n20297),
	.b(n20296));
   na02f10 U19684 (.o(n20366),
	.a(n19702),
	.b(n20370));
   na02f10 U19685 (.o(n20370),
	.a(n19701),
	.b(n23326));
   na02f10 U19686 (.o(n23292),
	.a(n19275),
	.b(n19274));
   no02f10 U19687 (.o(n18012),
	.a(n25406),
	.b(n18013));
   no02f10 U19688 (.o(n18014),
	.a(n24977),
	.b(n25406));
   in01f20 U19689 (.o(n17759),
	.a(validOut_P));
   oa22f02 U19690 (.o(north_output_control_N467),
	.a(n25139),
	.b(n17889),
	.c(n25138),
	.d(n25137));
   ao22f02 U19691 (.o(n25139),
	.a(n25135),
	.b(n18275),
	.c(n25136),
	.d(n18274));
   in01f02 U19692 (.o(n18200),
	.a(n18201));
   oa12f08 U19693 (.o(n17889),
	.a(n17888),
	.b(n18287),
	.c(n25083));
   no04f04 U19694 (.o(n20533),
	.a(n25177),
	.b(n20535),
	.c(n20534),
	.d(n20532));
   ao12f02 U19695 (.o(n20456),
	.a(n25177),
	.b(FE_OFN250_n25152),
	.c(n20530));
   no02f10 U19696 (.o(n18434),
	.a(n19739),
	.b(n19740));
   ao22f08 U19697 (.o(n19601),
	.a(FE_OCPN25968_n19500),
	.b(proc_input_NIB_storage_data_f_12__63_),
	.c(n19769),
	.d(proc_input_NIB_storage_data_f_14__63_));
   na02f10 U19699 (.o(n18253),
	.a(n21865),
	.b(north_input_NIB_storage_data_f_2__59_));
   na02f04 U19700 (.o(n23526),
	.a(n19958),
	.b(n19957));
   na04f10 U19701 (.o(n17999),
	.a(n18355),
	.b(n18000),
	.c(n17737),
	.d(n17736));
   na02f08 U19702 (.o(n17736),
	.a(proc_input_NIB_storage_data_f_7__44_),
	.b(FE_OFN20_n17779));
   na02f10 U19703 (.o(n17737),
	.a(proc_input_NIB_storage_data_f_3__44_),
	.b(n21768));
   ao22f06 U19704 (.o(n19557),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__34_),
	.c(n19769),
	.d(proc_input_NIB_storage_data_f_14__34_));
   ao22f04 U19705 (.o(n19636),
	.a(FE_OCPN25963_n18039),
	.b(proc_input_NIB_storage_data_f_10__52_),
	.c(FE_OFN25673_n18033),
	.d(proc_input_NIB_storage_data_f_11__52_));
   no02f04 U19706 (.o(n19783),
	.a(n19775),
	.b(n19774));
   no03f08 U19707 (.o(n20378),
	.a(n24998),
	.b(n23482),
	.c(n25405));
   in01f02 U19708 (.o(n18555),
	.a(n20383));
   na02f10 U19709 (.o(n18070),
	.a(n18072),
	.b(n18071));
   no02f08 U19711 (.o(n17853),
	.a(n19700),
	.b(n19693));
   no03f04 U19712 (.o(n25390),
	.a(n25389),
	.b(n25396),
	.c(n25388));
   ao22f08 U19713 (.o(n19619),
	.a(n18016),
	.b(n18020),
	.c(n17914),
	.d(n18024));
   na02f08 U19714 (.o(n19549),
	.a(myLocY_f_2_),
	.b(n23973));
   na02f06 U19715 (.o(n18738),
	.a(myLocX_f_2_),
	.b(n18744));
   no02f08 U19717 (.o(n19851),
	.a(n19086),
	.b(n18733));
   ao22f06 U19718 (.o(n18739),
	.a(n21365),
	.b(south_input_NIB_storage_data_f_2__42_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__42_));
   in01f03 U19719 (.o(n19325),
	.a(myLocY_f_0_));
   na02f03 U19720 (.o(n25114),
	.a(n20466),
	.b(n20467));
   no02f08 U19721 (.o(n20154),
	.a(myLocY_f_1_),
	.b(n22837));
   na03f06 U19722 (.o(n20224),
	.a(n24998),
	.b(n24997),
	.c(n25405));
   na02f08 U19723 (.o(n18240),
	.a(n18527),
	.b(FE_OFN428_n22902));
   ao22f02 U19724 (.o(n20039),
	.a(n21768),
	.b(proc_input_NIB_storage_data_f_3__25_),
	.c(FE_OFN156_n24129),
	.d(proc_input_NIB_storage_data_f_1__25_));
   ao22f08 U19725 (.o(n18975),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__36_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__36_));
   ao22f04 U19726 (.o(n19534),
	.a(n17779),
	.b(proc_input_NIB_storage_data_f_7__38_),
	.c(FE_OFN188_n24453),
	.d(proc_input_NIB_storage_data_f_2__38_));
   ao22f04 U19727 (.o(n18319),
	.a(proc_input_NIB_storage_data_f_8__41_),
	.b(FE_OFN169_n24343),
	.c(proc_input_NIB_storage_data_f_4__41_),
	.d(n17744));
   ao22f04 U19728 (.o(n19204),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__42_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__42_));
   ao22f04 U19729 (.o(n18370),
	.a(proc_input_NIB_storage_data_f_0__43_),
	.b(FE_OCPN25933_n24342),
	.c(proc_input_NIB_storage_data_f_13__43_),
	.d(FE_OFN191_n24454));
   ao22f04 U19731 (.o(n18162),
	.a(proc_input_NIB_storage_data_f_13__56_),
	.b(FE_OFN25602_n19530),
	.c(proc_input_NIB_storage_data_f_6__56_),
	.d(n19503));
   na02f03 U19732 (.o(n17957),
	.a(proc_input_NIB_storage_data_f_7__59_),
	.b(FE_OFN20_n17779));
   na02f08 U19733 (.o(n19811),
	.a(myLocY_f_6_),
	.b(n23183));
   oa22f04 U19734 (.o(n18292),
	.a(n19057),
	.b(n25132),
	.c(n19056),
	.d(n25128));
   no02f01 U19735 (.o(n18602),
	.a(n18754),
	.b(n18603));
   no02f06 U19736 (.o(n25052),
	.a(proc_output_current_route_connection_1_),
	.b(n25422));
   no02f01 U19737 (.o(n17930),
	.a(FE_OFN24806_n19655),
	.b(n17931));
   no02f06 U19738 (.o(n18148),
	.a(n20506),
	.b(n19375));
   na02f08 U19739 (.o(n20252),
	.a(n19414),
	.b(n20240));
   no02f10 U19740 (.o(n25132),
	.a(n17812),
	.b(n17936));
   ao22f02 U19741 (.o(n19992),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__29_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__29_));
   ao22m02 U19742 (.o(n19974),
	.a(n19973),
	.b(south_input_NIB_storage_data_f_2__22_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__22_));
   in01f08 U19743 (.o(n17800),
	.a(n26020));
   na02f04 U19744 (.o(n19066),
	.a(proc_output_control_planned_f),
	.b(n18803));
   na02f08 U19745 (.o(n22517),
	.a(south_output_current_route_connection_2_),
	.b(n24953));
   ao22f02 U19746 (.o(n20016),
	.a(n21768),
	.b(proc_input_NIB_storage_data_f_3__22_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__22_));
   ao22f02 U19747 (.o(n19962),
	.a(FE_OCPN25941_n24965),
	.b(south_input_NIB_storage_data_f_3__25_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__25_));
   ao22m02 U19748 (.o(n19960),
	.a(FE_OCPN25941_n24965),
	.b(south_input_NIB_storage_data_f_3__27_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__27_));
   no03f20 U19749 (.o(n20424),
	.a(n18802),
	.b(n18801),
	.c(n18800));
   no03f10 U19750 (.o(n23185),
	.a(n19136),
	.b(n19135),
	.c(n19134));
   ao22f06 U19751 (.o(n19275),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__46_),
	.c(n19400),
	.d(east_input_NIB_storage_data_f_3__46_));
   na02f06 U19752 (.o(n18022),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__62_));
   in01f02 U19753 (.o(n18142),
	.a(n17889));
   oa12f04 U19754 (.o(n20618),
	.a(n19099),
	.b(north_input_control_thanks_all_f),
	.c(n19100));
   ao12f04 U19756 (.o(n18082),
	.a(n18083),
	.b(thanksIn_P),
	.c(n18128));
   no02f08 U19758 (.o(n25301),
	.a(n25008),
	.b(n25061));
   no02f08 U19759 (.o(n25152),
	.a(n20538),
	.b(n19445));
   no02m08 U19760 (.o(n25499),
	.a(n20123),
	.b(n19856));
   na03f10 U19761 (.o(n17876),
	.a(n17878),
	.b(n18224),
	.c(n17877));
   na04f20 U19762 (.o(n21508),
	.a(n19581),
	.b(n19580),
	.c(n19582),
	.d(n19583));
   no02f10 U19763 (.o(n19059),
	.a(north_output_current_route_connection_1_),
	.b(n19058));
   ao22s02 U19764 (.o(n21655),
	.a(proc_input_control_count_f_7_),
	.b(n21654),
	.c(n21653),
	.d(n21652));
   na02f04 U19765 (.o(n25421),
	.a(n25312),
	.b(n25037));
   no03f40 U19776 (.o(n24761),
	.a(FE_OFN25600_reset),
	.b(east_input_NIB_tail_ptr_f_1_),
	.c(n24920));
   in01f08 U19778 (.o(n19446),
	.a(n25152));
   ao22f08 U19786 (.o(n19211),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__45_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__45_));
   in01m10 U19793 (.o(n19635),
	.a(myChipID_f_6_));
   na02f03 U19800 (.o(n22902),
	.a(proc_input_valid),
	.b(n20620));
   na02f08 U19801 (.o(n18239),
	.a(n18419),
	.b(n17738));
   ao22f06 U19802 (.o(n17738),
	.a(proc_input_NIB_storage_data_f_4__57_),
	.b(n21749),
	.c(proc_input_NIB_storage_data_f_6__57_),
	.d(n19503));
   ao22f08 U19803 (.o(n18705),
	.a(south_input_NIB_storage_data_f_1__36_),
	.b(FE_OFN24742_n18683),
	.c(south_input_NIB_storage_data_f_0__36_),
	.d(n24472));
   no02f10 U19804 (.o(n20381),
	.a(n19730),
	.b(n19731));
   ao22f06 U19805 (.o(n19578),
	.a(proc_input_NIB_storage_data_f_13__61_),
	.b(n24454),
	.c(proc_input_NIB_storage_data_f_14__61_),
	.d(n19769));
   no02f10 U19806 (.o(n20407),
	.a(n20152),
	.b(n20377));
   no02f10 U19811 (.o(n18059),
	.a(n19719),
	.b(n23304));
   no02f08 U19812 (.o(n17915),
	.a(n19546),
	.b(n19545));
   ao12f08 U19813 (.o(n18826),
	.a(myLocX_f_2_),
	.b(FE_RN_58),
	.c(n18832));
   na02f04 U19814 (.o(n19568),
	.a(n19561),
	.b(n19742));
   no02f20 U19820 (.o(n19012),
	.a(n18469),
	.b(east_output_control_planned_f));
   oa12f06 U19821 (.o(n19312),
	.a(n19310),
	.b(n20506),
	.c(n19311));
   oa12f10 U19822 (.o(n19383),
	.a(n19381),
	.b(n20506),
	.c(n19382));
   oa12f10 U19823 (.o(n19271),
	.a(n19269),
	.b(n20506),
	.c(n19270));
   ao22f08 U19824 (.o(n19179),
	.a(FE_RN_10),
	.b(north_input_NIB_storage_data_f_3__57_),
	.c(FE_OFN24773_n19075),
	.d(north_input_NIB_storage_data_f_0__57_));
   na02f03 U19825 (.o(n20418),
	.a(n20417),
	.b(n20416));
   oa12f08 U19826 (.o(n18814),
	.a(n19066),
	.b(n20417),
	.c(n18409));
   ao22f08 U19827 (.o(n19571),
	.a(FE_OCPN25962_n18039),
	.b(proc_input_NIB_storage_data_f_10__58_),
	.c(FE_OFN168_n24343),
	.d(proc_input_NIB_storage_data_f_8__58_));
   no02f20 U19828 (.o(n18469),
	.a(n20437),
	.b(n18470));
   no04f10 U19830 (.o(n18071),
	.a(n18528),
	.b(n19594),
	.c(n18531),
	.d(n18532));
   na02f20 U19831 (.o(n18068),
	.a(n19594),
	.b(n18064));
   na03f04 U19832 (.o(n18427),
	.a(n18429),
	.b(n25180),
	.c(n18428));
   no02f04 U19833 (.o(n18497),
	.a(n18500),
	.b(n18498));
   no02m02 U19834 (.o(n25012),
	.a(n25414),
	.b(n25011));
   in01m02 U19835 (.o(n25055),
	.a(n25412));
   no02m02 U19836 (.o(n25014),
	.a(n25412),
	.b(n25414));
   na02f02 U19837 (.o(n18498),
	.a(n18499),
	.b(n17757));
   in01f02 U19838 (.o(n18197),
	.a(n18198));
   na03f06 U19839 (.o(n24956),
	.a(n24955),
	.b(n24961),
	.c(n18080));
   na02f02 U19840 (.o(n18193),
	.a(n20524),
	.b(n20505));
   no03f02 U19841 (.o(n25011),
	.a(n25010),
	.b(n25027),
	.c(n25009));
   no02f06 U19842 (.o(n25412),
	.a(n25010),
	.b(n25009));
   in01f02 U19843 (.o(n17757),
	.a(n25417));
   na02f08 U19844 (.o(n18209),
	.a(n17866),
	.b(n18210));
   ao22f08 U19845 (.o(n25128),
	.a(n20410),
	.b(n20179),
	.c(n20180),
	.d(n21893));
   no02f08 U19847 (.o(n20451),
	.a(n24996),
	.b(n24995));
   na02f03 U19848 (.o(n25065),
	.a(FE_OFN412_n21671),
	.b(n25393));
   in01f04 U19849 (.o(n25054),
	.a(n24995));
   in01m01 U19850 (.o(n18215),
	.a(n20262));
   no02f02 U19851 (.o(n19826),
	.a(n21907),
	.b(n20146));
   na03f06 U19852 (.o(n17938),
	.a(n18476),
	.b(n20450),
	.c(n17937));
   in01f02 U19853 (.o(n18535),
	.a(n20467));
   in01f02 U19854 (.o(n18471),
	.a(n18472));
   in01f02 U19855 (.o(n17937),
	.a(n18477));
   na02f02 U19856 (.o(n18214),
	.a(n20265),
	.b(FE_OFN24833_n25232));
   no02f03 U19858 (.o(n20265),
	.a(n20227),
	.b(n17813));
   in01f04 U19859 (.o(n19865),
	.a(n19864));
   in01f02 U19860 (.o(n18409),
	.a(n18410));
   na02f02 U19861 (.o(n17807),
	.a(n20300),
	.b(n17808));
   no02m02 U19862 (.o(n19855),
	.a(n19837),
	.b(n19836));
   in01m01 U19863 (.o(n18478),
	.a(n19885));
   in01f04 U19864 (.o(n19790),
	.a(n19824));
   oa12f02 U19865 (.o(n22934),
	.a(n22900),
	.b(FE_OFN947_n25096),
	.c(n22901));
   in01f03 U19866 (.o(n19703),
	.a(n19722));
   in01m01 U19867 (.o(n18476),
	.a(n20191));
   no02m02 U19868 (.o(n20420),
	.a(n20276),
	.b(n20275));
   na03f02 U19869 (.o(dataOut_P_32_),
	.a(n23491),
	.b(n23490),
	.c(n23489));
   na03f02 U19870 (.o(dataOut_E_32_),
	.a(n21429),
	.b(n21428),
	.c(n21427));
   in01m01 U19871 (.o(n18538),
	.a(n19853));
   in01f01 U19872 (.o(n18557),
	.a(n20382));
   na03f02 U19873 (.o(dataOut_N_32_),
	.a(n21444),
	.b(n21443),
	.c(n21442));
   na03f02 U19874 (.o(dataOut_W_32_),
	.a(n21732),
	.b(n21731),
	.c(n21730));
   in01f01 U19875 (.o(n20331),
	.a(n20330));
   no02f02 U19876 (.o(n18410),
	.a(n18812),
	.b(n18813));
   na03f02 U19877 (.o(dataOut_S_32_),
	.a(n22308),
	.b(n22307),
	.c(n22306));
   in01s01 U19878 (.o(n20440),
	.a(n20429));
   in01m02 U19879 (.o(n20519),
	.a(n20513));
   in01f03 U19880 (.o(n18376),
	.a(n19739));
   na03m02 U19881 (.o(n19835),
	.a(n25247),
	.b(n20423),
	.c(n23481));
   na03f02 U19882 (.o(n19854),
	.a(n19847),
	.b(n19846),
	.c(n19845));
   no03f10 U19883 (.o(n18009),
	.a(n23528),
	.b(n23536),
	.c(n23520));
   na02f01 U19884 (.o(n25006),
	.a(n25005),
	.b(n25029));
   no02f01 U19885 (.o(n20191),
	.a(n19883),
	.b(n19882));
   na02m01 U19886 (.o(n20291),
	.a(n20269),
	.b(n24993));
   oa12f04 U19887 (.o(n20283),
	.a(n20279),
	.b(n20281),
	.c(n20280));
   in01f01 U19888 (.o(n20275),
	.a(n20274));
   no02f01 U19889 (.o(n23594),
	.a(n18101),
	.b(n18029));
   no03f01 U19890 (.o(n23315),
	.a(n23314),
	.b(n23313),
	.c(n23312));
   no02f08 U19891 (.o(n19004),
	.a(n19874),
	.b(n19878));
   in01m02 U19892 (.o(n19955),
	.a(n19911));
   na02f03 U19893 (.o(n20144),
	.a(n19819),
	.b(n19818));
   no02m01 U19894 (.o(n25230),
	.a(FE_OFN24831_n25232),
	.b(n25229));
   na02f08 U19895 (.o(n20229),
	.a(n20185),
	.b(n20183));
   na02f02 U19896 (.o(n20502),
	.a(n20138),
	.b(n19054));
   in01s01 U19897 (.o(n20136),
	.a(n20138));
   in01f03 U19898 (.o(n19045),
	.a(n19044));
   in01f01 U19899 (.o(n20447),
	.a(n20446));
   in01m02 U19900 (.o(n19867),
	.a(n20182));
   no02f02 U19901 (.o(n24719),
	.a(n24320),
	.b(n24319));
   no02f02 U19902 (.o(n24645),
	.a(n24162),
	.b(n24161));
   no02f02 U19903 (.o(n24584),
	.a(n24116),
	.b(n24115));
   no02f06 U19904 (.o(n24749),
	.a(n24207),
	.b(n24206));
   no02f04 U19905 (.o(n23567),
	.a(n21824),
	.b(n21823));
   no02f04 U19906 (.o(n24018),
	.a(n21358),
	.b(n21357));
   no02f06 U19907 (.o(n24683),
	.a(n24254),
	.b(n24253));
   no02f06 U19908 (.o(n24759),
	.a(n24389),
	.b(n24388));
   no02f02 U19909 (.o(n24729),
	.a(n24185),
	.b(n24184));
   no02f04 U19910 (.o(n24627),
	.a(n24231),
	.b(n24230));
   no02f02 U19911 (.o(n23576),
	.a(n21801),
	.b(n21800));
   no02f06 U19912 (.o(n23154),
	.a(n21755),
	.b(n21754));
   in01f01 U19913 (.o(n23481),
	.a(n20424));
   no02f04 U19914 (.o(n24606),
	.a(n24276),
	.b(n24275));
   no02f04 U19915 (.o(n20061),
	.a(n20060),
	.b(n20059));
   no02f06 U19916 (.o(n24593),
	.a(n24298),
	.b(n24297));
   na02f03 U19917 (.o(n20214),
	.a(n19020),
	.b(n20213));
   no02m01 U19918 (.o(n21381),
	.a(FE_OFN24831_n25232),
	.b(n21380));
   no02f08 U19919 (.o(n19876),
	.a(n19001),
	.b(n19883));
   no02f06 U19920 (.o(n20190),
	.a(n19873),
	.b(n18988));
   no02f06 U19921 (.o(n18437),
	.a(n18438),
	.b(n20186));
   in01f08 U19922 (.o(n17822),
	.a(n17823));
   na02f03 U19923 (.o(n20324),
	.a(n19019),
	.b(n20213));
   na02f08 U19924 (.o(n20247),
	.a(n19280),
	.b(n19267));
   no02m01 U19925 (.o(n25730),
	.a(n25728),
	.b(n25727));
   na02f06 U19926 (.o(n20570),
	.a(n23987),
	.b(n21893));
   no02m01 U19927 (.o(n25792),
	.a(n25791),
	.b(n25790));
   na02f08 U19928 (.o(n24992),
	.a(n25247),
	.b(n20424));
   in01f06 U19929 (.o(n17815),
	.a(n18291));
   no02f06 U19930 (.o(n20167),
	.a(n19118),
	.b(n19127));
   no02f06 U19931 (.o(n20168),
	.a(n19119),
	.b(n19094));
   in01f01 U19932 (.o(n19819),
	.a(n19813));
   na02s02 U19933 (.o(n19818),
	.a(n19817),
	.b(n19816));
   no02f02 U19934 (.o(n24027),
	.a(n21856),
	.b(n21855));
   no02f04 U19935 (.o(n23982),
	.a(n21308),
	.b(n21307));
   no02f02 U19936 (.o(n24710),
	.a(n24071),
	.b(n24070));
   no02f04 U19937 (.o(n24692),
	.a(n24047),
	.b(n24046));
   no02f04 U19938 (.o(n24670),
	.a(n24094),
	.b(n24093));
   no02f02 U19939 (.o(n24739),
	.a(n24356),
	.b(n24355));
   no02f04 U19940 (.o(n17864),
	.a(n23524),
	.b(n23957));
   no03f10 U19941 (.o(n19834),
	.a(n18785),
	.b(n18784),
	.c(n18783));
   in01f02 U19942 (.o(n17841),
	.a(n17976));
   in01f10 U19945 (.o(n22877),
	.a(n18708));
   in01f04 U19947 (.o(n17821),
	.a(n19516));
   na02f08 U19948 (.o(n17820),
	.a(n19515),
	.b(n19509));
   in01f02 U19949 (.o(n24996),
	.a(n25051));
   no02f03 U19950 (.o(n17884),
	.a(n19720),
	.b(n23294));
   ao22m01 U19951 (.o(n21159),
	.a(n21565),
	.b(n23623),
	.c(FE_OFN575_n25463),
	.d(n21903));
   in01m02 U19952 (.o(n19472),
	.a(n23710));
   no02f04 U19955 (.o(n22939),
	.a(n18551),
	.b(n18548));
   in01f04 U19956 (.o(n18882),
	.a(n22820));
   na02f04 U19957 (.o(n18440),
	.a(FE_OFN67_n19548),
	.b(n23966));
   no02f04 U19958 (.o(n18988),
	.a(n19132),
	.b(n19003));
   in01f06 U19959 (.o(n19002),
	.a(n20759));
   no03m01 U19960 (.o(n20228),
	.a(n21426),
	.b(n23479),
	.c(n25051));
   na02f08 U19961 (.o(n20243),
	.a(n19328),
	.b(n19327));
   ao12f02 U19962 (.o(n19813),
	.a(n19810),
	.b(n19812),
	.c(n19811));
   no02f04 U19964 (.o(n20007),
	.a(n24970),
	.b(n23984));
   in01f08 U19965 (.o(n19294),
	.a(n23322));
   no02f04 U19966 (.o(n23987),
	.a(n19894),
	.b(n17865));
   na02f01 U19967 (.o(n25511),
	.a(n19152),
	.b(n19151));
   na02f08 U19968 (.o(n18775),
	.a(n18771),
	.b(n18770));
   in01f02 U19969 (.o(n19240),
	.a(n19239));
   in01f08 U19970 (.o(n18761),
	.a(n18755));
   ao22m01 U19971 (.o(n25813),
	.a(ec_cfg_14_),
	.b(n25812),
	.c(n25811),
	.d(n25810));
   na02f06 U19972 (.o(n23488),
	.a(n19102),
	.b(n19101));
   na02f02 U19973 (.o(n23343),
	.a(n21289),
	.b(n21288));
   na02m02 U19974 (.o(n23511),
	.a(n21295),
	.b(n21294));
   no03f10 U19975 (.o(n23035),
	.a(n19109),
	.b(n19108),
	.c(n19107));
   ao22m01 U19976 (.o(n25751),
	.a(ec_cfg_5_),
	.b(n25750),
	.c(n25749),
	.d(n25748));
   na02f08 U19977 (.o(n20912),
	.a(n19316),
	.b(n19315));
   no02m01 U19978 (.o(n21895),
	.a(n21891),
	.b(n21890));
   na02f03 U19979 (.o(n23710),
	.a(n19256),
	.b(n19255));
   no03f08 U19980 (.o(n20408),
	.a(n19116),
	.b(n19115),
	.c(n19114));
   na02f10 U19981 (.o(n23965),
	.a(n19318),
	.b(n19317));
   na02f02 U19982 (.o(n18548),
	.a(n18550),
	.b(n18549));
   na02f10 U19983 (.o(n18716),
	.a(n18710),
	.b(n18709));
   in01f08 U19984 (.o(n18802),
	.a(n18796));
   na02f02 U19985 (.o(n19025),
	.a(n19024),
	.b(n19023));
   in01f01 U19987 (.o(n21638),
	.a(n21678));
   no02f02 U19988 (.o(n19256),
	.a(n19254),
	.b(n19253));
   no02m01 U19989 (.o(n21538),
	.a(FE_OFN24831_n25232),
	.b(n20616));
   oa12m01 U19990 (.o(n25819),
	.a(n20498),
	.b(n20500),
	.c(n20499));
   no02m01 U19991 (.o(n22072),
	.a(n22071),
	.b(n22070));
   in01f03 U19993 (.o(n18784),
	.a(n18780));
   na02f06 U19994 (.o(n20211),
	.a(n20422),
	.b(n20463));
   ao22f01 U19995 (.o(n25815),
	.a(n25359),
	.b(n25358),
	.c(n25357),
	.d(n25356));
   in01f02 U19996 (.o(n19141),
	.a(n19140));
   in01s02 U19997 (.o(n18551),
	.a(n19060));
   no03f10 U19998 (.o(n22843),
	.a(n19273),
	.b(n19272),
	.c(n19271));
   in01f04 U20000 (.o(n21672),
	.a(n19019));
   no02f04 U20001 (.o(n19136),
	.a(FE_OFN24776_n19073),
	.b(n19078));
   no02f04 U20002 (.o(n19135),
	.a(FE_OFN176_n24364),
	.b(n19079));
   oa22m02 U20003 (.o(n19253),
	.a(n19456),
	.b(n22518),
	.c(n19455),
	.d(n21667));
   no02m01 U20004 (.o(n25448),
	.a(n25446),
	.b(n25445));
   no02m01 U20005 (.o(n22073),
	.a(n22066),
	.b(n22069));
   no02m01 U20006 (.o(n25363),
	.a(n25361),
	.b(n25360));
   na02f01 U20007 (.o(n21586),
	.a(n25433),
	.b(FE_OFN100_n21907));
   oa22f02 U20008 (.o(n18789),
	.a(n19453),
	.b(n25027),
	.c(n19455),
	.d(n25411));
   oa22f02 U20009 (.o(n18788),
	.a(n19456),
	.b(n20501),
	.c(n19452),
	.d(n25029));
   no02f10 U20010 (.o(n25521),
	.a(n25130),
	.b(n19058));
   in01f06 U20011 (.o(n21662),
	.a(FE_OFN45_n19054));
   in01m06 U20013 (.o(n19016),
	.a(n19015));
   na02f06 U20014 (.o(n25474),
	.a(n25475),
	.b(n18791));
   in01f02 U20015 (.o(n25008),
	.a(n18790));
   in01m04 U20016 (.o(n18819),
	.a(n18816));
   in01m06 U20017 (.o(n18810),
	.a(n18809));
   in01m06 U20018 (.o(n18811),
	.a(n18808));
   in01m01 U20019 (.o(n25972),
	.a(n25974));
   in01f02 U20020 (.o(n23928),
	.a(dataIn_P_41_));
   in01m03 U20021 (.o(n23808),
	.a(dataIn_P_42_));
   in01m03 U20022 (.o(n23806),
	.a(dataIn_P_43_));
   in01f02 U20023 (.o(n23920),
	.a(dataIn_P_44_));
   in01f02 U20024 (.o(n23942),
	.a(dataIn_P_45_));
   in01m03 U20025 (.o(n23916),
	.a(dataIn_P_46_));
   in01m03 U20026 (.o(n23914),
	.a(dataIn_P_47_));
   in01f03 U20027 (.o(n23912),
	.a(dataIn_P_48_));
   in01m03 U20028 (.o(n23908),
	.a(dataIn_P_49_));
   in01m03 U20029 (.o(n23903),
	.a(dataIn_P_50_));
   in01m03 U20030 (.o(n23947),
	.a(dataIn_P_51_));
   in01m03 U20031 (.o(n23890),
	.a(dataIn_P_52_));
   in01f02 U20032 (.o(n23922),
	.a(dataIn_P_53_));
   in01f03 U20033 (.o(n23910),
	.a(dataIn_P_55_));
   in01f02 U20034 (.o(n23930),
	.a(dataIn_P_56_));
   in01m03 U20035 (.o(n23932),
	.a(dataIn_P_57_));
   in01m03 U20036 (.o(n23936),
	.a(dataIn_P_58_));
   in01m03 U20037 (.o(n23938),
	.a(dataIn_P_59_));
   in01m03 U20038 (.o(n23926),
	.a(dataIn_P_60_));
   in01m03 U20039 (.o(n23918),
	.a(dataIn_P_61_));
   in01f03 U20040 (.o(n23810),
	.a(dataIn_P_62_));
   in01m03 U20041 (.o(n23827),
	.a(dataIn_P_63_));
   in01f02 U20042 (.o(n23820),
	.a(dataIn_P_22_));
   in01f02 U20043 (.o(n23793),
	.a(dataIn_P_23_));
   in01f02 U20044 (.o(n23802),
	.a(dataIn_P_25_));
   in01f02 U20045 (.o(n23818),
	.a(dataIn_P_26_));
   in01f02 U20046 (.o(n23822),
	.a(dataIn_P_27_));
   in01m03 U20047 (.o(n23814),
	.a(dataIn_P_28_));
   in01f02 U20048 (.o(n23804),
	.a(dataIn_P_29_));
   in01f02 U20049 (.o(n23894),
	.a(dataIn_P_30_));
   in01m03 U20050 (.o(n23905),
	.a(dataIn_P_32_));
   in01m03 U20051 (.o(n23816),
	.a(dataIn_P_34_));
   in01m03 U20052 (.o(n23944),
	.a(dataIn_P_35_));
   in01m03 U20053 (.o(n23940),
	.a(dataIn_P_36_));
   in01f02 U20054 (.o(n23796),
	.a(dataIn_P_37_));
   in01m03 U20055 (.o(n23812),
	.a(dataIn_P_38_));
   in01f02 U20056 (.o(n23800),
	.a(dataIn_P_40_));
   na02f04 U20057 (.o(n25291),
	.a(n25432),
	.b(n25290));
   in01f04 U20058 (.o(n25286),
	.a(n25432));
   no02f04 U20059 (.o(n25293),
	.a(n25432),
	.b(n25280));
   no02f02 U20060 (.o(n18189),
	.a(n18191),
	.b(n18190));
   no02f02 U20061 (.o(n18186),
	.a(n18188),
	.b(n18187));
   no02f02 U20062 (.o(n18188),
	.a(n18193),
	.b(n18194));
   na02f02 U20063 (.o(n20525),
	.a(n25316),
	.b(n25147));
   na02f02 U20065 (.o(n18567),
	.a(n24979),
	.b(n18568));
   in01f06 U20066 (.o(n20313),
	.a(n25396));
   na02f08 U20067 (.o(n25147),
	.a(n20505),
	.b(n25329));
   na02f04 U20068 (.o(n20314),
	.a(n25393),
	.b(n20555));
   na03f10 U20069 (.o(n25396),
	.a(n20226),
	.b(n18209),
	.c(n18207));
   no02f02 U20070 (.o(n18276),
	.a(n25130),
	.b(n25128));
   in01f03 U20072 (.o(n18570),
	.a(n20344));
   in01m01 U20073 (.o(n25416),
	.a(n25415));
   no02f02 U20074 (.o(n20556),
	.a(n25393),
	.b(n20550));
   in01f06 U20075 (.o(n18625),
	.a(n20116));
   na02f02 U20076 (.o(n23549),
	.a(validOut_P),
	.b(FE_OFN25599_reset));
   no02m02 U20077 (.o(n18499),
	.a(n25408),
	.b(n25407));
   ao22f04 U20078 (.o(n24995),
	.a(n20450),
	.b(n20449),
	.c(n20448),
	.d(n20447));
   no02f06 U20079 (.o(n20335),
	.a(n19835),
	.b(n25155));
   no03f08 U20080 (.o(n20336),
	.a(n18536),
	.b(n22912),
	.c(n18535));
   ao22f06 U20081 (.o(n17939),
	.a(n20450),
	.b(n18471),
	.c(n19872),
	.d(n20448));
   no03f02 U20082 (.o(n20516),
	.a(n18074),
	.b(n20512),
	.c(n20513));
   na02f02 U20083 (.o(n25159),
	.a(n25158),
	.b(n25157));
   na02f04 U20084 (.o(n18534),
	.a(n20334),
	.b(FE_OFN428_n22902));
   na02f03 U20085 (.o(n18354),
	.a(n25116),
	.b(n25117));
   in01f06 U20086 (.o(n25026),
	.a(n25078));
   na02f06 U20087 (.o(n17829),
	.a(n20442),
	.b(n20463));
   no02f03 U20088 (.o(n25158),
	.a(n20422),
	.b(n20421));
   in01f04 U20089 (.o(n19832),
	.a(n19831));
   na02m02 U20090 (.o(n18168),
	.a(n20117),
	.b(n19956));
   ao12f04 U20091 (.o(n18536),
	.a(n18537),
	.b(n19854),
	.c(n19855));
   no02f03 U20092 (.o(n18477),
	.a(n18479),
	.b(n18478));
   in01f08 U20093 (.o(n18123),
	.a(n19741));
   ao12f04 U20094 (.o(n20421),
	.a(n20418),
	.b(n20420),
	.c(n20419));
   no02f08 U20095 (.o(n20208),
	.a(n19520),
	.b(n19519));
   no04f10 U20096 (.o(n19831),
	.a(n20415),
	.b(n19829),
	.c(n19830),
	.d(n20286));
   oa12f04 U20097 (.o(n20143),
	.a(n19807),
	.b(n19809),
	.c(n19808));
   in01f02 U20098 (.o(n19520),
	.a(n19740));
   na02f10 U20099 (.o(n19741),
	.a(n19543),
	.b(n18374));
   in01m01 U20100 (.o(n18539),
	.a(n19852));
   in01f08 U20101 (.o(n25079),
	.a(FE_RN_16));
   no02f02 U20102 (.o(n18475),
	.a(n19879),
	.b(n20231));
   ao12f04 U20103 (.o(n25028),
	.a(n20006),
	.b(n20007),
	.c(n21539));
   na02f10 U20104 (.o(n20231),
	.a(n19876),
	.b(n19004));
   no04f04 U20105 (.o(n19868),
	.a(n19867),
	.b(n19881),
	.c(n20229),
	.d(n19866));
   in01f08 U20106 (.o(n19789),
	.a(n19785));
   na02f08 U20107 (.o(n19543),
	.a(FE_OFN63_n19518),
	.b(n22931));
   na03f03 U20108 (.o(n18812),
	.a(n17774),
	.b(n23036),
	.c(n20269));
   no02f01 U20110 (.o(n20276),
	.a(n20273),
	.b(n20272));
   in01m02 U20111 (.o(n20306),
	.a(n20404));
   oa12f01 U20112 (.o(n22083),
	.a(n21906),
	.b(n21908),
	.c(FE_OFN100_n21907));
   no02f01 U20113 (.o(n21682),
	.a(n21681),
	.b(n21680));
   na02f01 U20114 (.o(n25500),
	.a(FE_OFN24830_n25499),
	.b(n18093));
   na02f10 U20115 (.o(n23520),
	.a(n20062),
	.b(n20061));
   na02f08 U20116 (.o(n23536),
	.a(n20046),
	.b(n20045));
   na02f10 U20117 (.o(n23528),
	.a(n20032),
	.b(n20031));
   no03m02 U20118 (.o(n20157),
	.a(n20168),
	.b(n20154),
	.c(n20153));
   no02m01 U20119 (.o(n25005),
	.a(n24993),
	.b(n24992));
   ao22f01 U20120 (.o(n21444),
	.a(n19059),
	.b(n24993),
	.c(n19057),
	.d(n23487));
   na02f06 U20121 (.o(n18011),
	.a(n23991),
	.b(FE_OFN428_n22902));
   na03f20 U20122 (.o(n23189),
	.a(n17824),
	.b(n17822),
	.c(n17819));
   no02f01 U20123 (.o(n23593),
	.a(n23592),
	.b(n23591));
   no02m02 U20124 (.o(n20423),
	.a(n23036),
	.b(n24993));
   na04f10 U20125 (.o(n18778),
	.a(n23036),
	.b(n20272),
	.c(n19828),
	.d(n20285));
   in01f06 U20126 (.o(n18713),
	.a(n19036));
   na02f02 U20127 (.o(n20172),
	.a(n20168),
	.b(n20167));
   na02f06 U20128 (.o(n19031),
	.a(n25247),
	.b(n20465));
   no02m01 U20129 (.o(n21383),
	.a(n21382),
	.b(n21381));
   in01f01 U20130 (.o(n20280),
	.a(n20278));
   na02f06 U20131 (.o(n20181),
	.a(n18437),
	.b(n18440));
   no02m02 U20132 (.o(n20414),
	.a(n20277),
	.b(n20285));
   oa22m01 U20133 (.o(n22658),
	.a(n24996),
	.b(n22771),
	.c(n23036),
	.d(n21695));
   oa22f08 U20134 (.o(n19803),
	.a(n19326),
	.b(n20912),
	.c(n19325),
	.d(n19324));
   na02f08 U20135 (.o(n19822),
	.a(n19329),
	.b(n20243));
   in01f02 U20136 (.o(n20409),
	.a(n19245));
   no02f06 U20137 (.o(n20395),
	.a(n17884),
	.b(n20304));
   no02f06 U20138 (.o(n19911),
	.a(n19472),
	.b(n23711));
   na02f10 U20139 (.o(n20433),
	.a(n19729),
	.b(n18882));
   na02f06 U20140 (.o(n19866),
	.a(n18088),
	.b(n18084));
   no02f06 U20141 (.o(n20465),
	.a(n19834),
	.b(n20424));
   no02f06 U20142 (.o(n20138),
	.a(n22939),
	.b(n19063));
   no02f04 U20143 (.o(n20031),
	.a(n20030),
	.b(n20029));
   no02f06 U20144 (.o(n23964),
	.a(n20092),
	.b(n20091));
   oa22m01 U20145 (.o(n21482),
	.a(n23036),
	.b(n25095),
	.c(n24996),
	.d(n21661));
   no02f08 U20146 (.o(n18160),
	.a(n18164),
	.b(n18161));
   oa22m01 U20147 (.o(n21479),
	.a(n24996),
	.b(n21672),
	.c(n23036),
	.d(FE_OFN412_n21671));
   in01f01 U20149 (.o(n18439),
	.a(n18440));
   oa12m02 U20150 (.o(n20305),
	.a(n20400),
	.b(n20304),
	.c(n20390));
   in01f02 U20151 (.o(n20246),
	.a(n20243));
   in01f02 U20152 (.o(n17862),
	.a(n19909));
   in01f02 U20153 (.o(n19977),
	.a(n20564));
   na02f08 U20154 (.o(n19267),
	.a(n19706),
	.b(n23501));
   no02f10 U20155 (.o(n20250),
	.a(n19706),
	.b(n23501));
   ao22f01 U20156 (.o(n24264),
	.a(n19056),
	.b(n24676),
	.c(FE_OFN366_n17753),
	.d(n24675));
   no02f08 U20157 (.o(n20242),
	.a(n19719),
	.b(FE_RN_61));
   no02f08 U20159 (.o(n19278),
	.a(n19701),
	.b(n23322));
   no02f06 U20160 (.o(n19245),
	.a(n20737),
	.b(n23488));
   ao22f01 U20161 (.o(n24437),
	.a(FE_OFN366_n17753),
	.b(n24750),
	.c(n19057),
	.d(FE_OFN546_n24751));
   no02m02 U20162 (.o(n25001),
	.a(n20238),
	.b(n21907));
   no02f06 U20163 (.o(n19279),
	.a(n19720),
	.b(n23292));
   na02f08 U20164 (.o(n17968),
	.a(n17970),
	.b(n17969));
   ao22f01 U20165 (.o(n20742),
	.a(FE_OFN366_n17753),
	.b(n23968),
	.c(n19057),
	.d(n23966));
   na02m02 U20166 (.o(n20029),
	.a(n20028),
	.b(n20027));
   no02f10 U20167 (.o(n20281),
	.a(n18738),
	.b(n18737));
   no02f10 U20168 (.o(n18326),
	.a(n19708),
	.b(n23493));
   in01f08 U20169 (.o(n18749),
	.a(n23493));
   na02f02 U20170 (.o(n20044),
	.a(n20040),
	.b(n20039));
   no02f08 U20171 (.o(n20196),
	.a(n21426),
	.b(n25051));
   no02f06 U20172 (.o(n20213),
	.a(n20319),
	.b(n23398));
   na02f08 U20173 (.o(n18846),
	.a(n19328),
	.b(n20928));
   in01m06 U20174 (.o(n19234),
	.a(n23500));
   ao22f01 U20175 (.o(n24445),
	.a(FE_OFN47_n19056),
	.b(FE_OFN517_n24712),
	.c(FE_OFN366_n17753),
	.d(n24711));
   oa12s01 U20176 (.o(ec_out_2_),
	.a(n25771),
	.b(ec_cfg_8_),
	.c(n25772));
   ao22f01 U20178 (.o(n24194),
	.a(n19056),
	.b(FE_OFN521_n24723),
	.c(FE_OFN366_n17753),
	.d(n24722));
   na02f08 U20179 (.o(n19727),
	.a(n19675),
	.b(n19674));
   na02f02 U20180 (.o(n20053),
	.a(n20048),
	.b(n20047));
   in01f02 U20181 (.o(n18294),
	.a(n18295));
   na04f04 U20182 (.o(n20018),
	.a(n20011),
	.b(n20010),
	.c(n20009),
	.d(n20008));
   no02f08 U20183 (.o(n18717),
	.a(n19132),
	.b(n18716));
   no02f06 U20184 (.o(n20304),
	.a(FE_OFN25614_n19237),
	.b(n19701));
   na04f10 U20185 (.o(n19726),
	.a(n19679),
	.b(n19678),
	.c(n19677),
	.d(n19676));
   ao22f01 U20186 (.o(n21318),
	.a(n19056),
	.b(n23977),
	.c(FE_OFN366_n17753),
	.d(n23976));
   ao22f01 U20187 (.o(n24081),
	.a(n19056),
	.b(FE_OFN515_n24702),
	.c(FE_OFN366_n17753),
	.d(n24703));
   ao22f01 U20188 (.o(n21878),
	.a(FE_OFN366_n17753),
	.b(n23561),
	.c(n19057),
	.d(n23562));
   na02f08 U20189 (.o(n17996),
	.a(n18356),
	.b(n17997));
   ao22f01 U20190 (.o(n21368),
	.a(n19056),
	.b(FE_OFN487_n24013),
	.c(FE_OFN366_n17753),
	.d(n24012));
   na02f08 U20191 (.o(n17896),
	.a(n17898),
	.b(n17897));
   ao22f01 U20192 (.o(n24416),
	.a(FE_OFN47_n19056),
	.b(FE_OFN530_n24733),
	.c(FE_OFN366_n17753),
	.d(n24734));
   in01m01 U20193 (.o(n23397),
	.a(n20319));
   ao22f01 U20194 (.o(n24404),
	.a(FE_OFN47_n19056),
	.b(n24686),
	.c(FE_OFN366_n17753),
	.d(n24687));
   ao12m01 U20195 (.o(n20569),
	.a(n20568),
	.b(FE_OFN24831_n25232),
	.c(n23984));
   ao22f01 U20196 (.o(n24150),
	.a(FE_OFN44_n19054),
	.b(n24693),
	.c(FE_OFN366_n17753),
	.d(n24694));
   ao22f01 U20197 (.o(n21839),
	.a(n19056),
	.b(FE_OFN477_n23578),
	.c(FE_OFN366_n17753),
	.d(n23577));
   ao22f01 U20198 (.o(n24286),
	.a(FE_OFN366_n17753),
	.b(n24598),
	.c(n19057),
	.d(n24599));
   ao22f01 U20199 (.o(n24308),
	.a(n19056),
	.b(FE_OFN497_n24586),
	.c(FE_OFN366_n17753),
	.d(n24585));
   in01f04 U20200 (.o(n20926),
	.a(n18748));
   ao22f01 U20201 (.o(n24126),
	.a(n19056),
	.b(FE_OFN493_n24577),
	.c(FE_OFN366_n17753),
	.d(n24576));
   ao22m02 U20202 (.o(n21811),
	.a(FE_OFN366_n17753),
	.b(n23570),
	.c(n19057),
	.d(n23571));
   in01s01 U20203 (.o(n17869),
	.a(n20211));
   na02f04 U20204 (.o(n23535),
	.a(n19903),
	.b(n19904));
   no02f02 U20205 (.o(n19257),
	.a(n23711),
	.b(FE_OFN25651_n25499));
   na02f02 U20206 (.o(n18803),
	.a(n18793),
	.b(n18792));
   na02f04 U20207 (.o(n23300),
	.a(n19264),
	.b(n19263));
   na02f06 U20208 (.o(n25494),
	.a(n19460),
	.b(n19459));
   in01f06 U20209 (.o(n18769),
	.a(n18763));
   na02f10 U20211 (.o(n23322),
	.a(n19277),
	.b(n19276));
   na02f04 U20213 (.o(n23957),
	.a(n19901),
	.b(n19902));
   na02f08 U20214 (.o(n20928),
	.a(n18845),
	.b(n18844));
   na02f04 U20215 (.o(n25051),
	.a(n18962),
	.b(n18961));
   oa12s01 U20216 (.o(n20728),
	.a(n21379),
	.b(n20727),
	.c(n20726));
   na02f08 U20217 (.o(n19064),
	.a(n18751),
	.b(n18750));
   no03f10 U20219 (.o(n22820),
	.a(n18862),
	.b(n18861),
	.c(n18860));
   na02f02 U20220 (.o(n19894),
	.a(n19893),
	.b(n19892));
   na02f10 U20221 (.o(n18708),
	.a(n18703),
	.b(n18702));
   ao22m01 U20222 (.o(n25818),
	.a(n22381),
	.b(n22383),
	.c(n22380),
	.d(n22379));
   in01f03 U20224 (.o(n18844),
	.a(n18843));
   in01f04 U20225 (.o(n18760),
	.a(n18756));
   in01s01 U20228 (.o(n25141),
	.a(n17935));
   oa22m01 U20229 (.o(n25814),
	.a(n25376),
	.b(n25375),
	.c(n25374),
	.d(n25373));
   no02f02 U20230 (.o(n18793),
	.a(n18789),
	.b(n18788));
   no02f03 U20231 (.o(n19460),
	.a(n19458),
	.b(n19457));
   na02s02 U20232 (.o(n21379),
	.a(n20727),
	.b(n20726));
   no02s01 U20234 (.o(n17935),
	.a(FE_OFN25613_n17934),
	.b(FE_RN_28));
   no02f01 U20235 (.o(n22899),
	.a(n21659),
	.b(n21658));
   na02s02 U20237 (.o(n23553),
	.a(n23308),
	.b(n22500));
   in01f04 U20238 (.o(n21661),
	.a(n19057));
   oa22f02 U20239 (.o(n19457),
	.a(n19456),
	.b(n22773),
	.c(n19455),
	.d(n22772));
   in01s01 U20242 (.o(n20767),
	.a(FE_OFN100_n21907));
   na02f01 U20243 (.o(n20933),
	.a(n25826),
	.b(n20932));
   in01m06 U20244 (.o(n21673),
	.a(n19017));
   na02f02 U20245 (.o(n21910),
	.a(n21943),
	.b(n25976));
   na02s01 U20246 (.o(n19886),
	.a(n25232),
	.b(n24982));
   na02s02 U20247 (.o(n20633),
	.a(n20630),
	.b(n20624));
   no02f08 U20249 (.o(n25232),
	.a(n19453),
	.b(n20589));
   no02f10 U20250 (.o(n20379),
	.a(n18811),
	.b(n18810));
   in01s01 U20251 (.o(n19251),
	.a(n19249));
   in01f08 U20252 (.o(n19018),
	.a(n20266));
   in01f04 U20253 (.o(n18806),
	.a(n18805));
   in01f04 U20255 (.o(n18807),
	.a(n18804));
   na02f02 U20256 (.o(n20970),
	.a(validIn_S),
	.b(FE_OFN575_n25463));
   na02f02 U20257 (.o(n21051),
	.a(validIn_W),
	.b(FE_OFN571_n25463));
   in01s01 U20258 (.o(n21173),
	.a(n21172));
   in01s01 U20259 (.o(n25316),
	.a(validIn_E));
   na02f02 U20260 (.o(n20526),
	.a(n18189),
	.b(n18186));
   no03f02 U20261 (.o(n20347),
	.a(n20346),
	.b(n20345),
	.c(n18567));
   no02f02 U20262 (.o(n18638),
	.a(n18639),
	.b(n18507));
   in01m02 U20263 (.o(n25321),
	.a(n25338));
   na02f02 U20264 (.o(n25413),
	.a(n25412),
	.b(n25411));
   in01f02 U20265 (.o(n20554),
	.a(n20559));
   no03f04 U20266 (.o(n19857),
	.a(n20335),
	.b(n20336),
	.c(n18032));
   in01f02 U20267 (.o(n18199),
	.a(n20522));
   no02m02 U20268 (.o(n25419),
	.a(n25415),
	.b(n25410));
   na02f04 U20269 (.o(n20555),
	.a(FE_OFN565_n25385),
	.b(FE_OFN25642_n25062));
   in01f02 U20270 (.o(n20120),
	.a(n20119));
   na02f04 U20271 (.o(n25417),
	.a(n24996),
	.b(n25054));
   in01f08 U20272 (.o(n20344),
	.a(n24952));
   no02f04 U20274 (.o(n18401),
	.a(n21907),
	.b(n18404));
   no02f06 U20275 (.o(n24973),
	.a(n20336),
	.b(n20335));
   in01m01 U20276 (.o(n25386),
	.a(n25393));
   no02f04 U20277 (.o(n20426),
	.a(n25158),
	.b(n20425));
   no02f03 U20278 (.o(n25414),
	.a(n17760),
	.b(n25004));
   oa22f08 U20279 (.o(n24952),
	.a(n17760),
	.b(n18444),
	.c(n18445),
	.d(n18446));
   na02f06 U20280 (.o(n18139),
	.a(n17939),
	.b(n17938));
   no02f02 U20281 (.o(n20523),
	.a(n20516),
	.b(n20515));
   no02f02 U20282 (.o(n18403),
	.a(n20149),
	.b(n20150));
   in01f04 U20283 (.o(n18446),
	.a(n19826));
   no02f06 U20284 (.o(n20150),
	.a(n20145),
	.b(n20146));
   na02f02 U20285 (.o(n18553),
	.a(n17774),
	.b(n20225));
   no02f06 U20286 (.o(n20443),
	.a(n19869),
	.b(n18473));
   no02f08 U20287 (.o(n19793),
	.a(n19804),
	.b(n19790));
   ao22f04 U20288 (.o(n20308),
	.a(n20305),
	.b(n20306),
	.c(n20307),
	.d(n17807));
   ao12f04 U20289 (.o(n20210),
	.a(n20208),
	.b(n17827),
	.c(n20209));
   in01f04 U20290 (.o(n20268),
	.a(n20267));
   na03m02 U20291 (.o(n25118),
	.a(n19056),
	.b(n25117),
	.c(n25116));
   oa12m02 U20292 (.o(dataOut_S_56_),
	.a(n22625),
	.b(n23619),
	.c(FE_OFN25652_n25499));
   no02f02 U20293 (.o(n18537),
	.a(n18539),
	.b(n18538));
   in01f02 U20294 (.o(n19567),
	.a(n19566));
   oa12m02 U20295 (.o(dataOut_E_56_),
	.a(n21337),
	.b(n23619),
	.c(FE_OFN25895_n25395));
   na02f10 U20296 (.o(n19476),
	.a(n19820),
	.b(n19330));
   oa12f01 U20297 (.o(dataOut_W_56_),
	.a(n22286),
	.b(n23619),
	.c(FE_OFN25883_n19446));
   na04f02 U20298 (.o(n22060),
	.a(n21897),
	.b(n21896),
	.c(n21895),
	.d(n21894));
   oa12f01 U20299 (.o(FE_OFN679_dataOut_S_42),
	.a(n21602),
	.b(n22850),
	.c(FE_OFN266_n25499));
   oa12m02 U20300 (.o(dataOut_P_56_),
	.a(n23618),
	.b(n23619),
	.c(FE_OFN24730_n));
   no02f08 U20301 (.o(n17827),
	.a(n19741),
	.b(n18375));
   na02f02 U20302 (.o(n18141),
	.a(n19824),
	.b(n19825));
   oa12f01 U20303 (.o(FE_OFN755_dataOut_W_42),
	.a(n22628),
	.b(n22850),
	.c(FE_OFN25880_n19446));
   na02f02 U20304 (.o(n20117),
	.a(n20330),
	.b(n22216));
   oa12f01 U20305 (.o(FE_OFN607_dataOut_E_42),
	.a(n20931),
	.b(n22850),
	.c(FE_OFN25891_n25395));
   oa12f01 U20306 (.o(FE_OFN829_dataOut_P_42),
	.a(n22849),
	.b(n22850),
	.c(n24728));
   na02f04 U20307 (.o(n18473),
	.a(n18475),
	.b(n18474));
   oa12f01 U20309 (.o(dataOut_N_56_),
	.a(n21341),
	.b(n23619),
	.c(FE_OFN25981_n21666));
   oa12f01 U20310 (.o(FE_OFN290_dataOut_N_42),
	.a(n21140),
	.b(n22850),
	.c(n21666));
   oa12f02 U20311 (.o(dataOut_S_57_),
	.a(n21614),
	.b(FE_OCPN25821_n19632),
	.c(FE_OFN25652_n25499));
   oa12f01 U20312 (.o(dataOut_N_57_),
	.a(n20647),
	.b(FE_OCPN25821_n19632),
	.c(FE_OFN25978_n21666));
   oa12m01 U20313 (.o(ec_out_0_),
	.a(n25733),
	.b(ec_cfg_2_),
	.c(n25734));
   oa12f01 U20314 (.o(dataOut_E_57_),
	.a(n20733),
	.b(FE_OCPN25821_n19632),
	.c(FE_OFN25895_n25395));
   no02f02 U20315 (.o(n20207),
	.a(n20200),
	.b(n20199));
   oa12f01 U20316 (.o(FE_OFN611_dataOut_E_38),
	.a(n21147),
	.b(n18031),
	.c(FE_OFN25891_n25395));
   oa12f02 U20317 (.o(dataOut_P_57_),
	.a(n22872),
	.b(FE_OCPN25821_n19632),
	.c(FE_OFN524_n24728));
   na02f01 U20318 (.o(n21894),
	.a(n21893),
	.b(n21892));
   oa12f01 U20319 (.o(FE_OFN294_dataOut_N_38),
	.a(n21144),
	.b(n18031),
	.c(n21666));
   in01f02 U20320 (.o(n19869),
	.a(n19868));
   oa12f02 U20321 (.o(dataOut_W_57_),
	.a(n22539),
	.b(FE_OCPN25821_n19632),
	.c(FE_OFN25883_n19446));
   in01f04 U20322 (.o(n18118),
	.a(n18119));
   no03f10 U20323 (.o(n19330),
	.a(n19789),
	.b(n19803),
	.c(n19822));
   ao12m02 U20324 (.o(n19885),
	.a(n20189),
	.b(n19878),
	.c(n19877));
   no02f06 U20325 (.o(n18375),
	.a(n19541),
	.b(n18376));
   oa12f01 U20326 (.o(FE_OFN292_dataOut_N_39),
	.a(n20765),
	.b(n22857),
	.c(n21666));
   oa12f01 U20327 (.o(FE_OFN25723_dataOut_W_31),
	.a(n22659),
	.b(n24998),
	.c(FE_OFN25880_n19446));
   oa12f01 U20328 (.o(FE_OFN25703_dataOut_N_37),
	.a(n20787),
	.b(n18104),
	.c(FE_OFN25869_n21666));
   oa12f02 U20329 (.o(dataOut_W_29_),
	.a(n22232),
	.b(FE_OFN142_n23964),
	.c(FE_OFN25880_n19446));
   oa12f01 U20330 (.o(FE_OFN25715_dataOut_W_37),
	.a(n22770),
	.b(n18104),
	.c(FE_OFN25880_n19446));
   oa12f01 U20331 (.o(dataOut_E_62_),
	.a(n21551),
	.b(n22896),
	.c(FE_OFN25895_n25395));
   oa12f01 U20332 (.o(dataOut_P_60_),
	.a(n23547),
	.b(n18102),
	.c(FE_OFN24730_n));
   oa12f01 U20333 (.o(FE_OFN705_dataOut_S_24),
	.a(n22438),
	.b(FE_OFN155_n24036),
	.c(FE_OFN266_n25499));
   oa12f01 U20334 (.o(FE_OFN763_dataOut_W_36),
	.a(n22236),
	.b(n23973),
	.c(FE_OFN25880_n19446));
   oa12f01 U20335 (.o(FE_OFN707_dataOut_S_23),
	.a(n22508),
	.b(n23628),
	.c(FE_OFN266_n25499));
   oa22f01 U20336 (.o(n21139),
	.a(n22844),
	.b(n25095),
	.c(n22843),
	.d(n21662));
   no02f04 U20337 (.o(n18119),
	.a(n18883),
	.b(n18884));
   oa12f01 U20338 (.o(dataOut_N_60_),
	.a(n20751),
	.b(n18102),
	.c(FE_OFN25980_n21666));
   oa12f01 U20339 (.o(dataOut_P_62_),
	.a(n22895),
	.b(n22896),
	.c(FE_OFN24730_n));
   oa12f01 U20340 (.o(FE_OFN767_dataOut_W_34),
	.a(n22776),
	.b(n22834),
	.c(FE_OFN25880_n19446));
   oa12f01 U20341 (.o(FE_OFN757_dataOut_W_39),
	.a(n22759),
	.b(n22857),
	.c(FE_OFN25880_n19446));
   oa12f01 U20342 (.o(FE_OFN25721_dataOut_N_31),
	.a(n21483),
	.b(n24998),
	.c(FE_OFN25869_n21666));
   oa12f01 U20343 (.o(FE_OFN316_dataOut_N_23),
	.a(n21398),
	.b(n23628),
	.c(n21666));
   oa12f01 U20344 (.o(FE_OFN314_dataOut_N_24),
	.a(n21448),
	.b(FE_OFN155_n24036),
	.c(n21666));
   oa12f01 U20345 (.o(dataOut_N_62_),
	.a(n21411),
	.b(n22896),
	.c(FE_OFN25979_n21666));
   oa12m02 U20346 (.o(FE_OFN308_dataOut_N_29),
	.a(n20964),
	.b(FE_OFN142_n23964),
	.c(n21666));
   oa12f01 U20347 (.o(FE_OFN25713_dataOut_W_48),
	.a(n22662),
	.b(n22865),
	.c(FE_OFN25880_n19446));
   oa12f01 U20348 (.o(FE_OFN781_dataOut_W_24),
	.a(n22442),
	.b(FE_OFN155_n24036),
	.c(FE_OFN25880_n19446));
   oa12f01 U20349 (.o(FE_OFN25709_dataOut_W_49),
	.a(n22491),
	.b(n22826),
	.c(FE_OFN25880_n19446));
   oa12f01 U20350 (.o(FE_OFN310_dataOut_N_28),
	.a(n21137),
	.b(n23956),
	.c(n21666));
   oa12f01 U20351 (.o(FE_OFN783_dataOut_W_23),
	.a(n22228),
	.b(n23628),
	.c(FE_OFN25880_n19446));
   oa12f01 U20352 (.o(FE_OFN298_dataOut_N_36),
	.a(n20744),
	.b(n23973),
	.c(n21666));
   oa12f01 U20353 (.o(FE_OFN773_dataOut_W_28),
	.a(n22224),
	.b(n23956),
	.c(FE_OFN25880_n19446));
   oa12f01 U20354 (.o(dataOut_W_62_),
	.a(n22767),
	.b(n22896),
	.c(FE_OFN25883_n19446));
   oa22f01 U20355 (.o(n22627),
	.a(n22843),
	.b(n24731),
	.c(n22844),
	.d(n21695));
   in01s01 U20356 (.o(n20376),
	.a(n20375));
   oa12f01 U20357 (.o(FE_OFN302_dataOut_N_34),
	.a(n20922),
	.b(n22834),
	.c(n21666));
   oa12f01 U20358 (.o(dataOut_W_60_),
	.a(n22536),
	.b(n18102),
	.c(FE_OFN25883_n19446));
   na02f08 U20359 (.o(n19702),
	.a(n19720),
	.b(n23296));
   oa12f01 U20360 (.o(FE_OFN25711_dataOut_P_49),
	.a(n22825),
	.b(n22826),
	.c(n24728));
   oa12f01 U20361 (.o(FE_OFN25725_dataOut_E_37),
	.a(n20790),
	.b(n18104),
	.c(FE_OFN569_n25395));
   oa12f01 U20362 (.o(FE_OFN831_dataOut_P_39),
	.a(n22856),
	.b(n22857),
	.c(n24728));
   no02f03 U20363 (.o(n20221),
	.a(n20381),
	.b(n20374));
   in01f02 U20364 (.o(n18223),
	.a(n20198));
   oa12f01 U20365 (.o(FE_OFN665_dataOut_S_49),
	.a(n21599),
	.b(n22826),
	.c(FE_OFN25651_n25499));
   oa12f01 U20366 (.o(FE_OFN615_dataOut_E_36),
	.a(n20777),
	.b(n23973),
	.c(FE_OFN25891_n25395));
   oa12f01 U20367 (.o(FE_OFN25886_dataOut_S_48),
	.a(n21611),
	.b(n22865),
	.c(FE_OFN25651_n25499));
   oa12f01 U20368 (.o(FE_OFN847_dataOut_P_28),
	.a(n23955),
	.b(n23956),
	.c(n24728));
   oa12f01 U20369 (.o(FE_OFN25717_dataOut_P_37),
	.a(n22880),
	.b(n18104),
	.c(n24728));
   oa22f01 U20370 (.o(n21601),
	.a(n22843),
	.b(n22518),
	.c(n22844),
	.d(FE_OFN24835_n22517));
   oa12f01 U20371 (.o(FE_OFN619_dataOut_E_34),
	.a(n20925),
	.b(n22834),
	.c(FE_OFN25891_n25395));
   oa12f01 U20372 (.o(FE_OFN837_dataOut_P_36),
	.a(n23972),
	.b(n23973),
	.c(n24728));
   oa12f01 U20373 (.o(FE_OFN681_dataOut_S_39),
	.a(n21622),
	.b(n22857),
	.c(FE_OFN266_n25499));
   oa22f01 U20374 (.o(n20930),
	.a(n22843),
	.b(n21673),
	.c(n22844),
	.d(FE_OFN412_n21671));
   oa22f01 U20375 (.o(n22848),
	.a(n22844),
	.b(n25029),
	.c(n22843),
	.d(FE_OFN902_n18421));
   oa12f01 U20376 (.o(dataOut_S_62_),
	.a(n21608),
	.b(n22896),
	.c(FE_OFN25652_n25499));
   oa12f01 U20377 (.o(dataOut_S_60_),
	.a(n22522),
	.b(n18102),
	.c(FE_OFN25652_n25499));
   oa12f01 U20378 (.o(FE_OFN855_dataOut_P_24),
	.a(n24035),
	.b(FE_OFN155_n24036),
	.c(n24728));
   oa12f02 U20379 (.o(dataOut_E_48_),
	.a(n21458),
	.b(n22865),
	.c(FE_OFN25891_n25395));
   no03f03 U20380 (.o(n20205),
	.a(n20203),
	.b(n20202),
	.c(n20201));
   oa12f02 U20381 (.o(dataOut_E_49_),
	.a(n20780),
	.b(n22826),
	.c(FE_OFN25891_n25395));
   oa12f01 U20382 (.o(FE_OFN25697_dataOut_E_39),
	.a(n20762),
	.b(n22857),
	.c(FE_OFN25891_n25395));
   oa12f01 U20383 (.o(FE_OFN857_dataOut_P_23),
	.a(n23627),
	.b(n23628),
	.c(n24728));
   oa12f01 U20384 (.o(FE_OFN25699_dataOut_P_48),
	.a(n22864),
	.b(n22865),
	.c(n24728));
   oa12f02 U20385 (.o(dataOut_E_31_),
	.a(n21480),
	.b(n24998),
	.c(FE_OFN569_n25395));
   oa12f01 U20386 (.o(FE_OFN697_dataOut_S_28),
	.a(n22504),
	.b(n23956),
	.c(FE_OFN266_n25499));
   oa12f01 U20387 (.o(FE_OFN631_dataOut_E_24),
	.a(n21452),
	.b(FE_OFN155_n24036),
	.c(FE_OFN25891_n25395));
   oa12f01 U20388 (.o(FE_OFN695_dataOut_S_29),
	.a(n22512),
	.b(FE_OFN142_n23964),
	.c(FE_OFN266_n25499));
   na02f01 U20389 (.o(n22324),
	.a(FE_OFN24829_n25499),
	.b(n23520));
   oa12f01 U20390 (.o(FE_OFN25884_dataOut_N_48),
	.a(n21455),
	.b(n22865),
	.c(FE_OFN25975_n21666));
   in01s01 U20391 (.o(n20337),
	.a(n23482));
   oa12f01 U20392 (.o(FE_OFN1006_dataOut_S_31),
	.a(n21605),
	.b(n24998),
	.c(FE_OFN25651_n25499));
   oa12f01 U20393 (.o(FE_OFN633_dataOut_E_23),
	.a(n21402),
	.b(n23628),
	.c(FE_OFN25891_n25395));
   oa12f01 U20394 (.o(dataOut_E_60_),
	.a(n20794),
	.b(n18102),
	.c(FE_OFN25895_n25395));
   oa12f02 U20395 (.o(dataOut_N_49_),
	.a(n20783),
	.b(n22826),
	.c(FE_OFN25975_n21666));
   oa12f01 U20396 (.o(FE_OFN691_dataOut_S_34),
	.a(n21631),
	.b(n22834),
	.c(FE_OFN266_n25499));
   oa12f01 U20397 (.o(FE_OFN841_dataOut_P_34),
	.a(n22833),
	.b(n22834),
	.c(n24728));
   oa12f01 U20398 (.o(FE_OFN687_dataOut_S_36),
	.a(n22529),
	.b(n23973),
	.c(FE_OFN266_n25499));
   oa12f01 U20399 (.o(FE_OFN685_dataOut_S_37),
	.a(n21596),
	.b(n18104),
	.c(FE_OFN25651_n25499));
   oa12f01 U20400 (.o(FE_OFN623_dataOut_E_29),
	.a(n20968),
	.b(FE_OFN142_n23964),
	.c(FE_OFN25891_n25395));
   oa12m02 U20401 (.o(FE_OFN625_dataOut_E_28),
	.a(n21133),
	.b(n23956),
	.c(FE_OFN25891_n25395));
   oa12m02 U20402 (.o(FE_OFN845_dataOut_P_29),
	.a(n23963),
	.b(FE_OFN142_n23964),
	.c(n24728));
   oa12f01 U20403 (.o(FE_OFN25727_dataOut_P_31),
	.a(n23039),
	.b(n24998),
	.c(n24728));
   ao22f01 U20404 (.o(n21339),
	.a(n17753),
	.b(n23614),
	.c(n19057),
	.d(n23612));
   ao22f01 U20405 (.o(n23350),
	.a(n25295),
	.b(n25516),
	.c(FE_OFN79_n20501),
	.d(n25497));
   no02f01 U20406 (.o(n21681),
	.a(n24036),
	.b(FE_OFN947_n25096));
   oa22f01 U20407 (.o(n22929),
	.a(n22928),
	.b(n25029),
	.c(n22927),
	.d(n25411));
   in01m01 U20408 (.o(n20198),
	.a(n20197));
   ao22f01 U20409 (.o(n22291),
	.a(n19493),
	.b(n23502),
	.c(FE_OFN105_n22517),
	.d(n23503));
   ao22m01 U20410 (.o(n22304),
	.a(FE_OFN105_n22517),
	.b(n23303),
	.c(FE_OFN93_n21667),
	.d(n23302));
   ao22f01 U20411 (.o(n22313),
	.a(n19493),
	.b(n23495),
	.c(FE_OFN93_n21667),
	.d(n23494));
   ao22f01 U20412 (.o(n22332),
	.a(FE_OFN105_n22517),
	.b(n23325),
	.c(n25498),
	.d(n23322));
   oa22s01 U20413 (.o(n21531),
	.a(n22927),
	.b(FE_OFN536_n24743),
	.c(n22926),
	.d(n24982));
   ao22f01 U20414 (.o(n23328),
	.a(n17787),
	.b(n23325),
	.c(n25294),
	.d(n23324));
   ao22f01 U20415 (.o(n22623),
	.a(FE_OFN105_n22517),
	.b(n23614),
	.c(FE_OFN577_n25498),
	.d(n23611));
   ao22f01 U20416 (.o(n23615),
	.a(FE_OFN25_n17787),
	.b(n23614),
	.c(n25294),
	.d(n23613));
   ao22m01 U20417 (.o(n23306),
	.a(n17787),
	.b(n23303),
	.c(n25294),
	.d(n23302));
   ao22m01 U20418 (.o(n22308),
	.a(FE_OFN105_n22517),
	.b(n24993),
	.c(n25498),
	.d(n23486));
   ao22f01 U20419 (.o(n23506),
	.a(n17787),
	.b(n23503),
	.c(FE_OFN259_n25295),
	.d(n23502));
   ao22f01 U20420 (.o(n21165),
	.a(n17753),
	.b(n23632),
	.c(n19057),
	.d(n23630));
   ao22f01 U20421 (.o(n22296),
	.a(FE_OFN396_n19493),
	.b(n23508),
	.c(FE_OFN105_n22517),
	.d(n22293));
   ao22f01 U20422 (.o(n23498),
	.a(FE_OFN259_n25295),
	.b(n23495),
	.c(n25294),
	.d(n23494));
   ao22f01 U20423 (.o(n21464),
	.a(n19059),
	.b(n23481),
	.c(n19057),
	.d(n23479));
   ao22f01 U20424 (.o(n21298),
	.a(FE_OFN42_n19022),
	.b(n22293),
	.c(n19019),
	.d(n23508));
   in01f04 U20425 (.o(n19882),
	.a(n19866));
   na02f06 U20427 (.o(n19879),
	.a(n20190),
	.b(n20184));
   ao22f01 U20428 (.o(n21335),
	.a(FE_OFN25872_FE_OFN42_n19022),
	.b(n23614),
	.c(n19019),
	.d(n23612));
   ao22f01 U20429 (.o(n21564),
	.a(n19056),
	.b(n23516),
	.c(n19057),
	.d(n23517));
   ao22f01 U20430 (.o(n21461),
	.a(n19022),
	.b(n23481),
	.c(n19019),
	.d(n23479));
   no02f06 U20431 (.o(n19820),
	.a(n19323),
	.b(n19808));
   na04f10 U20432 (.o(n19804),
	.a(n19439),
	.b(n19814),
	.c(n19812),
	.d(n19811));
   na02f01 U20433 (.o(n19845),
	.a(n19844),
	.b(n19843));
   in01s01 U20434 (.o(n19846),
	.a(n19838));
   ao22f01 U20435 (.o(n21394),
	.a(n19059),
	.b(n23325),
	.c(n19057),
	.d(n23323));
   ao22f01 U20436 (.o(n23490),
	.a(n17787),
	.b(n24993),
	.c(n25294),
	.d(n23488));
   ao22f01 U20437 (.o(n21429),
	.a(n19022),
	.b(n24993),
	.c(n19019),
	.d(n23487));
   oa22s01 U20439 (.o(n21541),
	.a(n22925),
	.b(n21662),
	.c(n22927),
	.d(FE_OFN563_n25120));
   oa12f04 U20440 (.o(n18883),
	.a(n20433),
	.b(n20430),
	.c(n20434));
   ao22f01 U20441 (.o(n21476),
	.a(n19057),
	.b(n23495),
	.c(n19056),
	.d(n23494));
   ao22f01 U20442 (.o(n21378),
	.a(n19022),
	.b(n23325),
	.c(n19019),
	.d(n23323));
   ao22f01 U20443 (.o(n21344),
	.a(n19017),
	.b(n23300),
	.c(n19020),
	.d(n23302));
   ao22f01 U20444 (.o(n21405),
	.a(n19022),
	.b(n23503),
	.c(n19019),
	.d(n23502));
   ao22f01 U20445 (.o(n21473),
	.a(n19019),
	.b(n23495),
	.c(n19020),
	.d(n23494));
   oa22s01 U20446 (.o(n21527),
	.a(n22925),
	.b(n21673),
	.c(n22927),
	.d(FE_OFN565_n25385));
   ao22f01 U20447 (.o(n21413),
	.a(n19059),
	.b(n23503),
	.c(n19057),
	.d(n23502));
   ao22f01 U20448 (.o(n21347),
	.a(n19054),
	.b(n23300),
	.c(n19056),
	.d(n23302));
   ao22f01 U20449 (.o(n21704),
	.a(FE_OFN111_n22773),
	.b(n23300),
	.c(n17755),
	.d(n23302));
   ao22f01 U20450 (.o(n21710),
	.a(FE_OFN94_n21695),
	.b(n23503),
	.c(n17786),
	.d(n23502));
   ao22f01 U20451 (.o(n21720),
	.a(FE_OFN94_n21695),
	.b(n22293),
	.c(FE_OFN389_n17786),
	.d(n23508));
   no02f08 U20452 (.o(n21539),
	.a(n20003),
	.b(n20002));
   ao22f01 U20453 (.o(n21728),
	.a(n17786),
	.b(n23495),
	.c(n17755),
	.d(n23494));
   oa22s01 U20454 (.o(n21523),
	.a(n22925),
	.b(n22773),
	.c(n22927),
	.d(n22772));
   ao22f01 U20455 (.o(n21708),
	.a(FE_OFN94_n21695),
	.b(n23481),
	.c(n17786),
	.d(n23479));
   ao22f01 U20456 (.o(n21328),
	.a(n17753),
	.b(n22293),
	.c(n19057),
	.d(n23508));
   ao22f01 U20457 (.o(n21732),
	.a(FE_OFN94_n21695),
	.b(n24993),
	.c(n17786),
	.d(n23487));
   in01f01 U20458 (.o(n20431),
	.a(n20430));
   na02f02 U20459 (.o(n18092),
	.a(n19621),
	.b(n19620));
   ao22f01 U20460 (.o(n22284),
	.a(FE_OFN94_n21695),
	.b(n23614),
	.c(FE_OFN389_n17786),
	.d(n23612));
   no02f06 U20461 (.o(n17861),
	.a(n17862),
	.b(n23620));
   ao22f01 U20462 (.o(n21702),
	.a(FE_OFN94_n21695),
	.b(n23325),
	.c(n17786),
	.d(n23323));
   ao22f01 U20463 (.o(n22906),
	.a(FE_OFN111_n22773),
	.b(n25497),
	.c(n17755),
	.d(n25518));
   ao22f01 U20464 (.o(n23515),
	.a(FE_OFN25_n17787),
	.b(n22293),
	.c(n25295),
	.d(n23508));
   oa22f01 U20465 (.o(n21600),
	.a(n22845),
	.b(FE_OFN539_n24743),
	.c(n22846),
	.d(FE_OFN247_n24982));
   oa22s01 U20466 (.o(n22871),
	.a(n22867),
	.b(n25029),
	.c(n22866),
	.d(FE_OFN78_n20501));
   oa22f01 U20467 (.o(n21630),
	.a(n22827),
	.b(n22518),
	.c(n22830),
	.d(FE_OFN24834_n22517));
   oa22f01 U20468 (.o(n21603),
	.a(n23035),
	.b(n21667),
	.c(n24996),
	.d(n24982));
   ao22s01 U20469 (.o(n23336),
	.a(n25295),
	.b(FE_RN_25),
	.c(FE_OFN79_n20501),
	.d(n23330));
   ao22f01 U20470 (.o(n22307),
	.a(n19493),
	.b(n23487),
	.c(FE_OFN93_n21667),
	.d(n23488));
   oa22f01 U20471 (.o(n22870),
	.a(n22869),
	.b(n25411),
	.c(n22868),
	.d(n25027));
   oa22f01 U20472 (.o(n23591),
	.a(n23590),
	.b(n25029),
	.c(n23589),
	.d(n25411));
   oa22f01 U20473 (.o(n21591),
	.a(n22883),
	.b(FE_OFN535_n24743),
	.c(n22882),
	.d(FE_OFN247_n24982));
   oa22f01 U20474 (.o(n21623),
	.a(FE_OFN25623_n19123),
	.b(FE_OFN533_n24743),
	.c(n22836),
	.d(FE_OFN247_n24982));
   no02s01 U20475 (.o(n18270),
	.a(n21485),
	.b(n25411));
   oa22f01 U20476 (.o(n21592),
	.a(n22881),
	.b(n22518),
	.c(n22884),
	.d(FE_OFN387_n17783));
   oa22f01 U20477 (.o(n21664),
	.a(n22760),
	.b(n25095),
	.c(n23993),
	.d(n21661));
   oa22f01 U20478 (.o(n23546),
	.a(n23541),
	.b(n25029),
	.c(n23540),
	.d(FE_OFN78_n20501));
   ao22f01 U20479 (.o(n21491),
	.a(n17753),
	.b(n18670),
	.c(n19057),
	.d(n23317));
   oa22f01 U20480 (.o(n21594),
	.a(n22876),
	.b(n24743),
	.c(n22875),
	.d(n24982));
   oa22f01 U20481 (.o(n21595),
	.a(n22874),
	.b(n22518),
	.c(n22877),
	.d(n22517));
   no02s01 U20482 (.o(n18261),
	.a(n21485),
	.b(FE_OFN563_n25120));
   oa22f01 U20483 (.o(n22894),
	.a(n22890),
	.b(n25027),
	.c(n22889),
	.d(FE_OFN902_n18421));
   oa22m01 U20484 (.o(n21532),
	.a(n22925),
	.b(n22518),
	.c(n22928),
	.d(n22517));
   oa22f01 U20485 (.o(n21604),
	.a(n23034),
	.b(n22518),
	.c(n23036),
	.d(n22517));
   oa22f01 U20486 (.o(n21629),
	.a(n22829),
	.b(FE_OFN538_n24743),
	.c(n22828),
	.d(FE_OFN247_n24982));
   oa22m01 U20488 (.o(n21501),
	.a(n23183),
	.b(n22518),
	.c(n23186),
	.d(n17783));
   na02f04 U20489 (.o(n20323),
	.a(n19022),
	.b(n20213));
   oa22f01 U20490 (.o(n21663),
	.a(n23992),
	.b(n21662),
	.c(n22761),
	.d(FE_OFN563_n25120));
   ao22s01 U20491 (.o(n22322),
	.a(n19493),
	.b(n23479),
	.c(FE_OFN93_n21667),
	.d(n23480));
   oa22f01 U20492 (.o(n21620),
	.a(n22853),
	.b(FE_OFN537_n24743),
	.c(n22852),
	.d(FE_OFN247_n24982));
   oa22f01 U20493 (.o(n21621),
	.a(n22851),
	.b(n22518),
	.c(n17751),
	.d(FE_OFN386_n17783));
   oa22f01 U20494 (.o(n24007),
	.a(n24002),
	.b(n25027),
	.c(FE_OFN25696_n19372),
	.d(FE_OFN902_n18421));
   oa22f01 U20495 (.o(n21409),
	.a(n22889),
	.b(n21662),
	.c(n22891),
	.d(FE_OFN563_n25120));
   oa22f01 U20496 (.o(n22626),
	.a(n22845),
	.b(n22772),
	.c(n22846),
	.d(FE_OFN110_n22771));
   oa22f01 U20497 (.o(n21410),
	.a(n22892),
	.b(n25095),
	.c(n22890),
	.d(n21661));
   ao22m01 U20498 (.o(n21725),
	.a(n17786),
	.b(n23295),
	.c(n17755),
	.d(n23294));
   oa22f01 U20499 (.o(n21513),
	.a(FE_OFN25696_n19372),
	.b(n21662),
	.c(n22753),
	.d(FE_OFN563_n25120));
   oa22f01 U20500 (.o(n21514),
	.a(n22752),
	.b(n25095),
	.c(n24002),
	.d(n21661));
   oa22m01 U20501 (.o(n22661),
	.a(n22859),
	.b(n22771),
	.c(n22861),
	.d(n21695));
   oa22m01 U20502 (.o(n22490),
	.a(n22820),
	.b(n22771),
	.c(n22822),
	.d(n21695));
   oa22m01 U20503 (.o(n22489),
	.a(n22819),
	.b(n22773),
	.c(n22821),
	.d(n22772));
   ao22f01 U20504 (.o(n21717),
	.a(FE_OFN94_n21695),
	.b(n23341),
	.c(FE_OFN389_n17786),
	.d(n23340));
   ao22f01 U20505 (.o(n21716),
	.a(FE_OFN111_n22773),
	.b(n23343),
	.c(n17755),
	.d(FE_OFN25630_n19165));
   in01f01 U20506 (.o(n20397),
	.a(n20390));
   oa22f01 U20507 (.o(n20750),
	.a(n23541),
	.b(n25095),
	.c(n23540),
	.d(n21662));
   ao22s01 U20508 (.o(n22909),
	.a(FE_OFN111_n22773),
	.b(n23330),
	.c(n17755),
	.d(n23331));
   no02f06 U20509 (.o(n18072),
	.a(n18529),
	.b(n18530));
   oa22f01 U20510 (.o(n22763),
	.a(n23993),
	.b(FE_OFN110_n22771),
	.c(n22760),
	.d(n21695));
   oa22f01 U20511 (.o(n22762),
	.a(n23992),
	.b(FE_OFN525_n24731),
	.c(n22761),
	.d(n22772));
   oa22f01 U20512 (.o(n22769),
	.a(n22875),
	.b(n22771),
	.c(n22877),
	.d(n21695));
   oa22f01 U20513 (.o(n22768),
	.a(n22874),
	.b(n22773),
	.c(n22876),
	.d(n22772));
   oa22f01 U20514 (.o(n22523),
	.a(n22835),
	.b(n22773),
	.c(FE_OFN25623_n19123),
	.d(n22772));
   oa22f01 U20515 (.o(n22524),
	.a(n22836),
	.b(n22771),
	.c(n22838),
	.d(n21695));
   oa22f01 U20516 (.o(n22531),
	.a(n22882),
	.b(FE_OFN110_n22771),
	.c(n22884),
	.d(n21695));
   oa22f01 U20517 (.o(n22774),
	.a(n22827),
	.b(FE_OFN112_n22773),
	.c(n22829),
	.d(n22772));
   oa22f01 U20518 (.o(n22775),
	.a(n22828),
	.b(FE_OFN110_n22771),
	.c(n22830),
	.d(n21695));
   oa22f01 U20519 (.o(n22530),
	.a(n22881),
	.b(n22773),
	.c(n22883),
	.d(n22772));
   oa22m01 U20520 (.o(n22757),
	.a(n22851),
	.b(n22773),
	.c(n22853),
	.d(n22772));
   oa22f01 U20521 (.o(n22657),
	.a(n23034),
	.b(n22773),
	.c(n23035),
	.d(n22772));
   oa22m01 U20522 (.o(n21493),
	.a(n23184),
	.b(n22771),
	.c(n23186),
	.d(n21695));
   oa22m01 U20523 (.o(n21524),
	.a(n22926),
	.b(n22771),
	.c(n22928),
	.d(n21695));
   na02f06 U20524 (.o(n20002),
	.a(n20001),
	.b(n20000));
   na02f04 U20525 (.o(n20003),
	.a(n21558),
	.b(n19991));
   oa22f01 U20526 (.o(n21421),
	.a(n23590),
	.b(n25095),
	.c(n21616),
	.d(n21661));
   na03f02 U20527 (.o(n19949),
	.a(n20766),
	.b(n21569),
	.c(n21582));
   oa22f01 U20528 (.o(n20645),
	.a(n22869),
	.b(FE_OFN563_n25120),
	.c(n22868),
	.d(n21661));
   oa22f01 U20529 (.o(n20646),
	.a(n22867),
	.b(n25095),
	.c(n22866),
	.d(n21662));
   no03f10 U20530 (.o(n19620),
	.a(n17971),
	.b(n17968),
	.c(n17965));
   ao22f01 U20531 (.o(n21714),
	.a(FE_OFN94_n21695),
	.b(n18670),
	.c(FE_OFN389_n17786),
	.d(n23317));
   no02s01 U20532 (.o(n18264),
	.a(n21485),
	.b(n22772));
   oa22f01 U20534 (.o(n22538),
	.a(n22866),
	.b(FE_OFN525_n24731),
	.c(n22867),
	.d(n21695));
   oa22f01 U20535 (.o(n22537),
	.a(n22869),
	.b(n22772),
	.c(n22868),
	.d(FE_OFN110_n22771));
   oa22f01 U20536 (.o(n21424),
	.a(n21616),
	.b(FE_OFN110_n22771),
	.c(n23590),
	.d(n21695));
   oa22f01 U20537 (.o(n22535),
	.a(n23540),
	.b(FE_OFN525_n24731),
	.c(n23541),
	.d(n21695));
   oa22f01 U20538 (.o(n22755),
	.a(n24002),
	.b(FE_OFN110_n22771),
	.c(n22752),
	.d(n21695));
   oa22f01 U20539 (.o(n22754),
	.a(FE_OFN25696_n19372),
	.b(FE_OFN525_n24731),
	.c(n22753),
	.d(n22772));
   oa22f01 U20540 (.o(n22766),
	.a(n22890),
	.b(FE_OFN110_n22771),
	.c(n22892),
	.d(n21695));
   oa22f01 U20541 (.o(n22765),
	.a(n22889),
	.b(FE_OFN525_n24731),
	.c(n22891),
	.d(n22772));
   oa22m01 U20542 (.o(n23187),
	.a(n23186),
	.b(n25029),
	.c(n23185),
	.d(n25411));
   oa22f01 U20543 (.o(n20731),
	.a(n22869),
	.b(FE_OFN565_n25385),
	.c(n22868),
	.d(n21672));
   oa22f01 U20544 (.o(n21481),
	.a(n23034),
	.b(n21662),
	.c(n23035),
	.d(FE_OFN563_n25120));
   oa22f01 U20545 (.o(n22854),
	.a(n17751),
	.b(n25029),
	.c(n22853),
	.d(n25411));
   oa22f01 U20546 (.o(n22855),
	.a(n22852),
	.b(n25027),
	.c(n22851),
	.d(n20501));
   oa22f01 U20547 (.o(n21505),
	.a(n23186),
	.b(n25095),
	.c(n23184),
	.d(n21661));
   oa22f01 U20548 (.o(n20921),
	.a(n22830),
	.b(n25095),
	.c(n22828),
	.d(n21661));
   oa22f01 U20549 (.o(n21542),
	.a(n22928),
	.b(n25095),
	.c(n22926),
	.d(n21661));
   in01m01 U20550 (.o(n19877),
	.a(n19873));
   oa22f01 U20551 (.o(n20913),
	.a(n22835),
	.b(n21673),
	.c(FE_OFN25623_n19123),
	.d(FE_OFN565_n25385));
   oa22f01 U20552 (.o(n20914),
	.a(n22836),
	.b(n21672),
	.c(n22838),
	.d(FE_OFN412_n21671));
   in01f02 U20553 (.o(n23519),
	.a(n21582));
   no02f10 U20554 (.o(n19795),
	.a(n19279),
	.b(n19278));
   oa22f01 U20555 (.o(n22847),
	.a(n22846),
	.b(n25027),
	.c(n22845),
	.d(n25411));
   in01f06 U20556 (.o(n17802),
	.a(n17803));
   oa22f01 U20557 (.o(n20923),
	.a(n22827),
	.b(n21673),
	.c(n22829),
	.d(FE_OFN565_n25385));
   oa22f01 U20558 (.o(n20924),
	.a(n22828),
	.b(n21672),
	.c(n22830),
	.d(FE_OFN412_n21671));
   ao12f06 U20559 (.o(n19281),
	.a(n20242),
	.b(n20250),
	.c(n19280));
   oa22f01 U20560 (.o(n20732),
	.a(n22866),
	.b(n21673),
	.c(n22867),
	.d(n21671));
   oa22f01 U20561 (.o(n21606),
	.a(n22891),
	.b(FE_OFN540_n24743),
	.c(n22890),
	.d(FE_OFN247_n24982));
   no02f06 U20562 (.o(n19794),
	.a(n19806),
	.b(n19815));
   oa22f01 U20563 (.o(n23038),
	.a(n24996),
	.b(n25027),
	.c(n23034),
	.d(n20501));
   oa22f01 U20564 (.o(n21418),
	.a(n21616),
	.b(n21672),
	.c(n23590),
	.d(n21671));
   in01s01 U20565 (.o(n21640),
	.a(n21651));
   ao22f01 U20566 (.o(n21330),
	.a(FE_OFN44_n19054),
	.b(n23343),
	.c(FE_OFN47_n19056),
	.d(FE_OFN25630_n19165));
   ao22m01 U20567 (.o(n21331),
	.a(n17753),
	.b(n23341),
	.c(n19057),
	.d(n23340));
   in01m01 U20568 (.o(n19844),
	.a(n19839));
   oa22m01 U20569 (.o(n23037),
	.a(n23036),
	.b(n25029),
	.c(n23035),
	.d(n25411));
   oa22f01 U20570 (.o(n22839),
	.a(n22838),
	.b(n25029),
	.c(FE_OFN25623_n19123),
	.d(n25411));
   oa22f01 U20571 (.o(n22840),
	.a(n22836),
	.b(n25027),
	.c(n22835),
	.d(n20501));
   oa22f01 U20572 (.o(n20786),
	.a(n22877),
	.b(n25095),
	.c(n22875),
	.d(n21661));
   oa22f01 U20573 (.o(n20793),
	.a(n23540),
	.b(n21673),
	.c(n23541),
	.d(n21671));
   oa22f01 U20574 (.o(n20785),
	.a(n22874),
	.b(n21662),
	.c(n22876),
	.d(FE_OFN563_n25120));
   oa22f01 U20575 (.o(n20781),
	.a(n22819),
	.b(n21662),
	.c(n22821),
	.d(FE_OFN563_n25120));
   oa22f01 U20576 (.o(n20782),
	.a(n22822),
	.b(n25095),
	.c(n22820),
	.d(n21661));
   oa22f01 U20577 (.o(n21143),
	.a(n22884),
	.b(n25095),
	.c(n22882),
	.d(n21661));
   oa22f01 U20578 (.o(n21142),
	.a(n22881),
	.b(n21662),
	.c(n22883),
	.d(FE_OFN563_n25120));
   oa22f01 U20579 (.o(n22831),
	.a(n22830),
	.b(n25029),
	.c(n22829),
	.d(n25411));
   oa22m01 U20580 (.o(n21454),
	.a(n22861),
	.b(n25095),
	.c(n22859),
	.d(n21661));
   oa22f01 U20581 (.o(n22832),
	.a(n22828),
	.b(n25027),
	.c(n22827),
	.d(n20501));
   no04m02 U20582 (.o(n19802),
	.a(n25003),
	.b(n23034),
	.c(n23486),
	.d(n21907));
   oa22f01 U20583 (.o(n21478),
	.a(n23034),
	.b(n21673),
	.c(n23035),
	.d(FE_OFN565_n25385));
   oa22f01 U20584 (.o(n22885),
	.a(n22884),
	.b(n25029),
	.c(n22883),
	.d(n25411));
   oa22f01 U20585 (.o(n20920),
	.a(n22827),
	.b(n21662),
	.c(n22829),
	.d(FE_OFN563_n25120));
   ao22m01 U20586 (.o(n21440),
	.a(n19057),
	.b(n23295),
	.c(n19056),
	.d(n23294));
   oa22f01 U20587 (.o(n21549),
	.a(n22889),
	.b(n21673),
	.c(n22891),
	.d(FE_OFN565_n25385));
   no03f20 U20588 (.o(n20284),
	.a(n18327),
	.b(n20281),
	.c(n18326));
   oa22f01 U20589 (.o(n22886),
	.a(n22882),
	.b(n25027),
	.c(n22881),
	.d(n20501));
   oa22f01 U20590 (.o(n21550),
	.a(n22890),
	.b(n21672),
	.c(n22892),
	.d(n21671));
   na02f08 U20591 (.o(n18965),
	.a(n19720),
	.b(n23295));
   oa22f01 U20592 (.o(n22878),
	.a(n22877),
	.b(n25029),
	.c(n22876),
	.d(n25411));
   na02f06 U20593 (.o(n19808),
	.a(n19322),
	.b(n19805));
   oa22f01 U20594 (.o(n20763),
	.a(n22851),
	.b(n21662),
	.c(n22853),
	.d(FE_OFN563_n25120));
   oa22f01 U20595 (.o(n20917),
	.a(n22838),
	.b(n25095),
	.c(n22836),
	.d(n21661));
   oa22f01 U20596 (.o(n22879),
	.a(n22875),
	.b(n25027),
	.c(n22874),
	.d(n20501));
   oa22f01 U20597 (.o(n21510),
	.a(FE_OFN25696_n19372),
	.b(n21673),
	.c(n22753),
	.d(FE_OFN565_n25385));
   oa22f01 U20598 (.o(n20916),
	.a(n22835),
	.b(n21662),
	.c(FE_OFN25623_n19123),
	.d(FE_OFN563_n25120));
   oa22f01 U20599 (.o(n21511),
	.a(n24002),
	.b(n21672),
	.c(n22752),
	.d(n21671));
   ao22f01 U20600 (.o(n21291),
	.a(FE_OFN35_n19017),
	.b(n23343),
	.c(n19020),
	.d(FE_OFN25630_n19165));
   oa22m01 U20601 (.o(n22823),
	.a(n22822),
	.b(n25029),
	.c(n22821),
	.d(n25411));
   oa22m01 U20602 (.o(n22862),
	.a(n22861),
	.b(n25029),
	.c(n22860),
	.d(n25411));
   oa22f01 U20603 (.o(n20929),
	.a(n22846),
	.b(n21672),
	.c(n22845),
	.d(FE_OFN565_n25385));
   ao22s01 U20604 (.o(n22311),
	.a(FE_OFN105_n22517),
	.b(n23332),
	.c(FE_OFN577_n25498),
	.d(n23330));
   in01f01 U20605 (.o(n23629),
	.a(n21163));
   oa22f01 U20606 (.o(n21669),
	.a(n23992),
	.b(FE_OFN108_n22518),
	.c(n22760),
	.d(FE_OFN24836_n22517));
   oa22f01 U20607 (.o(n21668),
	.a(n22761),
	.b(FE_OFN540_n24743),
	.c(n23993),
	.d(FE_OFN247_n24982));
   oa22s01 U20608 (.o(n21528),
	.a(n22926),
	.b(n21672),
	.c(n22928),
	.d(FE_OFN412_n21671));
   na02f06 U20609 (.o(n20170),
	.a(n19518),
	.b(n21522));
   ao22s01 U20610 (.o(n22317),
	.a(FE_OFN105_n22517),
	.b(n18670),
	.c(FE_OFN577_n25498),
	.d(n23316));
   oa22f01 U20611 (.o(n21497),
	.a(n23184),
	.b(n21672),
	.c(n23186),
	.d(FE_OFN412_n21671));
   no02s01 U20612 (.o(n18267),
	.a(n21485),
	.b(FE_OFN540_n24743));
   no02f08 U20613 (.o(n23991),
	.a(n20018),
	.b(n20017));
   oa22f01 U20614 (.o(n21138),
	.a(n22846),
	.b(n21661),
	.c(n22845),
	.d(FE_OFN563_n25120));
   oa22m01 U20615 (.o(n20760),
	.a(n22851),
	.b(n21673),
	.c(n22853),
	.d(FE_OFN565_n25385));
   ao22m01 U20616 (.o(n22319),
	.a(n19493),
	.b(n23295),
	.c(FE_OFN93_n21667),
	.d(n23294));
   oa22m01 U20617 (.o(n21457),
	.a(n22859),
	.b(n21672),
	.c(n22861),
	.d(FE_OFN412_n21671));
   oa22m01 U20618 (.o(n20779),
	.a(n22820),
	.b(n21672),
	.c(n22822),
	.d(FE_OFN412_n21671));
   ao22m01 U20619 (.o(n21149),
	.a(n19019),
	.b(n23295),
	.c(n19020),
	.d(n23294));
   oa22m01 U20620 (.o(n21610),
	.a(n22858),
	.b(n22518),
	.c(n22861),
	.d(FE_OFN106_n22517));
   oa22m01 U20621 (.o(n21598),
	.a(n22819),
	.b(n22518),
	.c(n22822),
	.d(FE_OFN106_n22517));
   oa22m01 U20622 (.o(n20778),
	.a(n22819),
	.b(n21673),
	.c(n22821),
	.d(FE_OFN565_n25385));
   ao22s01 U20623 (.o(n21467),
	.a(FE_OFN44_n19054),
	.b(n23330),
	.c(FE_OFN47_n19056),
	.d(n23331));
   ao22f01 U20624 (.o(n23346),
	.a(FE_OFN79_n20501),
	.b(n23343),
	.c(n25294),
	.d(FE_OFN25630_n19165));
   oa22m01 U20625 (.o(n21597),
	.a(n22821),
	.b(FE_OFN536_n24743),
	.c(n22820),
	.d(n24982));
   ao22m01 U20626 (.o(n23347),
	.a(FE_OFN25_n17787),
	.b(n23341),
	.c(n25295),
	.d(n23340));
   ao22s01 U20627 (.o(n22289),
	.a(FE_OFN396_n19493),
	.b(n23340),
	.c(FE_OFN105_n22517),
	.d(n23341));
   ao22f01 U20628 (.o(n22288),
	.a(FE_OFN577_n25498),
	.b(n23343),
	.c(FE_OFN93_n21667),
	.d(FE_OFN25630_n19165));
   ao22s01 U20629 (.o(n21292),
	.a(FE_OFN42_n19022),
	.b(n23341),
	.c(n19019),
	.d(n23340));
   oa22f01 U20630 (.o(n21145),
	.a(n22881),
	.b(n21673),
	.c(n22883),
	.d(FE_OFN565_n25385));
   oa22f01 U20631 (.o(n21618),
	.a(n21615),
	.b(FE_OFN108_n22518),
	.c(n23590),
	.d(FE_OFN24836_n22517));
   oa22f01 U20632 (.o(n21675),
	.a(n23993),
	.b(n21672),
	.c(n22760),
	.d(n21671));
   in01f01 U20633 (.o(n23534),
	.a(n21569));
   no02f04 U20634 (.o(n19120),
	.a(n19119),
	.b(n19118));
   oa22f01 U20635 (.o(n21674),
	.a(n23992),
	.b(n21673),
	.c(n22761),
	.d(FE_OFN565_n25385));
   oa22f01 U20636 (.o(n21146),
	.a(n22882),
	.b(n21672),
	.c(n22884),
	.d(FE_OFN412_n21671));
   no02f04 U20637 (.o(n20046),
	.a(n20038),
	.b(n20037));
   ao22s01 U20638 (.o(n21488),
	.a(FE_OFN42_n19022),
	.b(n18670),
	.c(n19019),
	.d(n23317));
   in01f06 U20639 (.o(n20434),
	.a(n18873));
   no02f02 U20640 (.o(n20045),
	.a(n20044),
	.b(n20043));
   no02s01 U20641 (.o(n18258),
	.a(n21485),
	.b(FE_OFN565_n25385));
   oa22f01 U20642 (.o(n22521),
	.a(n23540),
	.b(FE_OFN108_n22518),
	.c(n23541),
	.d(FE_OFN24836_n22517));
   oa22f01 U20643 (.o(n20788),
	.a(n22874),
	.b(n21673),
	.c(n22876),
	.d(FE_OFN565_n25385));
   oa22f01 U20644 (.o(n21627),
	.a(FE_OFN25696_n19372),
	.b(FE_OFN108_n22518),
	.c(n22752),
	.d(FE_OFN24836_n22517));
   in01f02 U20645 (.o(n22927),
	.a(n21522));
   oa22f01 U20646 (.o(n21626),
	.a(n22753),
	.b(FE_OFN540_n24743),
	.c(n24002),
	.d(FE_OFN247_n24982));
   oa22f01 U20647 (.o(n21607),
	.a(n22889),
	.b(FE_OFN108_n22518),
	.c(n22892),
	.d(FE_OFN24836_n22517));
   oa22f01 U20648 (.o(n21613),
	.a(n22866),
	.b(FE_OFN108_n22518),
	.c(n22867),
	.d(FE_OFN24836_n22517));
   oa22f01 U20649 (.o(n20789),
	.a(n22875),
	.b(n21672),
	.c(n22877),
	.d(FE_OFN412_n21671));
   ao22m01 U20650 (.o(n22493),
	.a(FE_OFN35_n19017),
	.b(n23330),
	.c(n19020),
	.d(n23331));
   oa22f01 U20651 (.o(n21612),
	.a(n22869),
	.b(FE_OFN540_n24743),
	.c(n22868),
	.d(FE_OFN247_n24982));
   ao22m01 U20652 (.o(n23298),
	.a(FE_OFN259_n25295),
	.b(n23295),
	.c(n25294),
	.d(n23294));
   no02f01 U20653 (.o(n21382),
	.a(n21558),
	.b(n24970));
   in01f06 U20654 (.o(n18308),
	.a(n19662));
   na02f02 U20655 (.o(n20037),
	.a(n20036),
	.b(n20035));
   in01f04 U20656 (.o(n17998),
	.a(n18357));
   no02f06 U20657 (.o(n20444),
	.a(n24970),
	.b(n23479));
   ao22f01 U20658 (.o(n21348),
	.a(n19059),
	.b(n23303),
	.c(n19057),
	.d(n23301));
   no02f08 U20659 (.o(n22821),
	.a(n19241),
	.b(n19240));
   na02f08 U20660 (.o(n17837),
	.a(n17975),
	.b(n17838));
   na02m02 U20661 (.o(n20038),
	.a(n20034),
	.b(n20033));
   ao22f01 U20662 (.o(n24104),
	.a(FE_OFN47_n19056),
	.b(n24663),
	.c(FE_OFN44_n19054),
	.d(FE_OFN221_n24662));
   no02f06 U20663 (.o(n18735),
	.a(n19325),
	.b(n20919));
   no02f06 U20664 (.o(n18296),
	.a(n18298),
	.b(n18297));
   ao22f01 U20665 (.o(n21414),
	.a(n19054),
	.b(n23501),
	.c(n19056),
	.d(n23500));
   no02f08 U20666 (.o(n19837),
	.a(n19321),
	.b(n18708));
   ao22f01 U20667 (.o(n21297),
	.a(FE_OFN35_n19017),
	.b(n23511),
	.c(n19020),
	.d(n23510));
   ao22f01 U20668 (.o(n20791),
	.a(n19019),
	.b(n23543),
	.c(n19020),
	.d(n23542));
   ao22m01 U20669 (.o(n25509),
	.a(FE_OFN25872_FE_OFN42_n19022),
	.b(n18028),
	.c(n19019),
	.d(n25516));
   na02f08 U20670 (.o(n17900),
	.a(n17902),
	.b(n17901));
   na02f02 U20671 (.o(n20043),
	.a(n20042),
	.b(n20041));
   ao22f01 U20673 (.o(n24436),
	.a(n19056),
	.b(n24754),
	.c(FE_OFN44_n19054),
	.d(n24752));
   ao22f01 U20674 (.o(n24149),
	.a(n19056),
	.b(FE_OFN513_n24695),
	.c(n19057),
	.d(n24696));
   ao22m01 U20675 (.o(n21521),
	.a(n19056),
	.b(n23524),
	.c(n19057),
	.d(n23525));
   ao22f01 U20676 (.o(n24217),
	.a(n19056),
	.b(n24742),
	.c(FE_OFN44_n19054),
	.d(FE_OFN242_n24744));
   oa12s01 U20677 (.o(n20738),
	.a(FE_OFN575_n25463),
	.b(n20737),
	.c(n23516));
   ao22f01 U20678 (.o(n24444),
	.a(FE_OFN44_n19054),
	.b(n24713),
	.c(n19057),
	.d(n24714));
   na02f06 U20679 (.o(n19700),
	.a(n19696),
	.b(n19695));
   no02f08 U20680 (.o(n19089),
	.a(n21141),
	.b(n19132));
   na03f06 U20681 (.o(n19479),
	.a(n25003),
	.b(n25002),
	.c(n20238));
   ao22m01 U20682 (.o(n21446),
	.a(n19057),
	.b(n24029),
	.c(n19059),
	.d(n24028));
   ao22m01 U20683 (.o(n21445),
	.a(n19056),
	.b(n24031),
	.c(n19054),
	.d(n24030));
   in01f10 U20684 (.o(n19150),
	.a(n23331));
   ao22f01 U20685 (.o(n21393),
	.a(n19054),
	.b(n23322),
	.c(n19056),
	.d(n23324));
   ao22f01 U20686 (.o(n25515),
	.a(n17753),
	.b(n25510),
	.c(n19057),
	.d(n21696));
   ao22m01 U20687 (.o(n21395),
	.a(n19054),
	.b(FE_OFN136_n23623),
	.c(n19059),
	.d(n23622));
   no02f08 U20688 (.o(n17803),
	.a(n19411),
	.b(n17804));
   ao22f01 U20689 (.o(n21396),
	.a(n19056),
	.b(n23620),
	.c(n19057),
	.d(n23621));
   na02f04 U20690 (.o(n19693),
	.a(n19692),
	.b(n19691));
   no02f04 U20691 (.o(n19094),
	.a(n19325),
	.b(n19122));
   ao22m01 U20692 (.o(n21557),
	.a(n19057),
	.b(n23533),
	.c(n19059),
	.d(n23532));
   ao22f01 U20693 (.o(n21468),
	.a(n17753),
	.b(n23332),
	.c(n19057),
	.d(FE_RN_25));
   ao22f01 U20694 (.o(n24285),
	.a(n19056),
	.b(FE_OFN499_n24601),
	.c(FE_OFN44_n19054),
	.d(FE_OFN203_n24600));
   ao22m01 U20695 (.o(n21435),
	.a(n19057),
	.b(n23984),
	.c(n19059),
	.d(n23983));
   in01f02 U20696 (.o(n23986),
	.a(n21431));
   no02f06 U20697 (.o(n20394),
	.a(n23500),
	.b(n19706));
   ao22f01 U20698 (.o(n24307),
	.a(n19054),
	.b(n24587),
	.c(n19057),
	.d(n24588));
   ao22m01 U20699 (.o(n21441),
	.a(n19059),
	.b(n23293),
	.c(n19054),
	.d(n23292));
   ao22f01 U20700 (.o(n21879),
	.a(FE_OFN47_n19056),
	.b(FE_OFN473_n23560),
	.c(FE_OFN44_n19054),
	.d(FE_OFN130_n23559));
   na04f04 U20701 (.o(n20091),
	.a(n20090),
	.b(n20089),
	.c(n20088),
	.d(n20087));
   ao22f01 U20702 (.o(n22622),
	.a(FE_OFN396_n19493),
	.b(n23612),
	.c(FE_OFN93_n21667),
	.d(n23613));
   ao22f01 U20703 (.o(n22310),
	.a(FE_OFN396_n19493),
	.b(FE_RN_25),
	.c(FE_OFN93_n21667),
	.d(n23331));
   ao22f01 U20704 (.o(n22328),
	.a(FE_OFN396_n19493),
	.b(n21696),
	.c(FE_OFN93_n21667),
	.d(FE_OFN579_n25511));
   ao22m01 U20705 (.o(n22329),
	.a(FE_OFN105_n22517),
	.b(n25510),
	.c(FE_OFN577_n25498),
	.d(n25512));
   oa22m01 U20706 (.o(n21609),
	.a(n22860),
	.b(FE_OFN536_n24743),
	.c(n22859),
	.d(n24982));
   na02f06 U20707 (.o(n17823),
	.a(n19517),
	.b(n19512));
   ao22s01 U20708 (.o(n22331),
	.a(n19493),
	.b(n23323),
	.c(FE_OFN93_n21667),
	.d(n23324));
   ao22m01 U20709 (.o(n22320),
	.a(FE_OFN105_n22517),
	.b(n23293),
	.c(n25498),
	.d(n23292));
   ao22f01 U20710 (.o(n22305),
	.a(n19493),
	.b(n23301),
	.c(n25498),
	.d(n23300));
   in01f02 U20711 (.o(n23480),
	.a(n20408));
   no02f01 U20712 (.o(n22496),
	.a(n22912),
	.b(n23518));
   ao22f01 U20713 (.o(n22292),
	.a(n25498),
	.b(n23501),
	.c(FE_OFN93_n21667),
	.d(n23500));
   ao22f01 U20714 (.o(n22314),
	.a(FE_OFN105_n22517),
	.b(n23493),
	.c(n25498),
	.d(n23492));
   ao22f01 U20715 (.o(n21545),
	.a(n17786),
	.b(n23984),
	.c(FE_OFN94_n21695),
	.d(n23983));
   oa22f01 U20716 (.o(n21504),
	.a(n23183),
	.b(n21662),
	.c(n23185),
	.d(FE_OFN563_n25120));
   ao12f01 U20717 (.o(n21391),
	.a(n21390),
	.b(n25247),
	.c(n23532));
   ao22f01 U20718 (.o(n22226),
	.a(n17786),
	.b(n23621),
	.c(n17755),
	.d(n23620));
   oa22m01 U20719 (.o(n21500),
	.a(n23185),
	.b(FE_OFN534_n24743),
	.c(n23184),
	.d(FE_OFN247_n24982));
   ao22f01 U20720 (.o(n22440),
	.a(n17786),
	.b(n24029),
	.c(FE_OFN94_n21695),
	.d(n24028));
   ao22f01 U20721 (.o(n23307),
	.a(FE_OFN259_n25295),
	.b(n23301),
	.c(FE_OFN79_n20501),
	.d(n23300));
   ao22m01 U20722 (.o(n23299),
	.a(n17787),
	.b(n23293),
	.c(FE_OFN79_n20501),
	.d(n23292));
   ao22s01 U20723 (.o(n23329),
	.a(FE_OFN259_n25295),
	.b(n23323),
	.c(FE_OFN79_n20501),
	.d(n23322));
   oa22m01 U20724 (.o(n22863),
	.a(n22859),
	.b(n25027),
	.c(n22858),
	.d(n20501));
   ao12s01 U20725 (.o(n21680),
	.a(FE_OFN428_n22902),
	.b(n21679),
	.c(n21678));
   oa22m01 U20726 (.o(n22824),
	.a(n22820),
	.b(n25027),
	.c(n22819),
	.d(n20501));
   ao22m01 U20727 (.o(n23339),
	.a(n25295),
	.b(n21696),
	.c(FE_OFN79_n20501),
	.d(n25512));
   ao22f01 U20728 (.o(n23338),
	.a(FE_OFN25_n17787),
	.b(n25510),
	.c(n25294),
	.d(FE_OFN579_n25511));
   na02f06 U20729 (.o(n18289),
	.a(n18315),
	.b(n18316));
   ao22s01 U20730 (.o(n23335),
	.a(FE_OFN25_n17787),
	.b(n23332),
	.c(n25294),
	.d(n23331));
   oa22m01 U20731 (.o(n23998),
	.a(n23993),
	.b(n25027),
	.c(n23992),
	.d(FE_OFN78_n20501));
   ao22s01 U20732 (.o(n23996),
	.a(n17787),
	.b(n23995),
	.c(n25294),
	.d(n23994));
   ao22f01 U20733 (.o(n20962),
	.a(n19056),
	.b(n23957),
	.c(n19057),
	.d(n25231));
   ao22f01 U20734 (.o(n20748),
	.a(n19057),
	.b(n23543),
	.c(FE_OFN47_n19056),
	.d(n23542));
   ao22s01 U20735 (.o(n23321),
	.a(n25295),
	.b(n23317),
	.c(FE_OFN79_n20501),
	.d(n23316));
   ao22f01 U20736 (.o(n23616),
	.a(n25295),
	.b(n23612),
	.c(FE_OFN79_n20501),
	.d(n23611));
   na02s01 U20737 (.o(n20772),
	.a(n20771),
	.b(FE_OFN100_n21907));
   ao22f01 U20738 (.o(n23588),
	.a(n25295),
	.b(n23587),
	.c(FE_OFN79_n20501),
	.d(n23586));
   ao22m01 U20739 (.o(n20961),
	.a(n19054),
	.b(FE_OFN140_n23959),
	.c(n19059),
	.d(n23958));
   ao22m01 U20740 (.o(n23349),
	.a(FE_OFN25_n17787),
	.b(n18028),
	.c(n25294),
	.d(n25518));
   ao22f01 U20741 (.o(n23544),
	.a(n25295),
	.b(n23543),
	.c(n25294),
	.d(n23542));
   ao22f01 U20742 (.o(n24005),
	.a(n17787),
	.b(n24004),
	.c(n25294),
	.d(n24003));
   ao22f01 U20744 (.o(n23514),
	.a(FE_OFN79_n20501),
	.b(n23511),
	.c(n25294),
	.d(n23510));
   ao22f01 U20745 (.o(n22295),
	.a(FE_OFN577_n25498),
	.b(n23511),
	.c(FE_OFN93_n21667),
	.d(n23510));
   ao22f01 U20746 (.o(n22519),
	.a(n19493),
	.b(n23543),
	.c(FE_OFN93_n21667),
	.d(n23542));
   ao22f01 U20747 (.o(n21871),
	.a(FE_OFN44_n19054),
	.b(FE_OFN151_n24019),
	.c(n19057),
	.d(n24020));
   ao22f01 U20748 (.o(n21699),
	.a(FE_OFN94_n21695),
	.b(n25510),
	.c(FE_OFN389_n17786),
	.d(n21696));
   ao22f01 U20749 (.o(n21698),
	.a(FE_OFN111_n22773),
	.b(n25512),
	.c(n17755),
	.d(FE_OFN579_n25511));
   ao22f01 U20750 (.o(n22910),
	.a(FE_OFN94_n21695),
	.b(n23332),
	.c(FE_OFN389_n17786),
	.d(FE_RN_25));
   na02m01 U20751 (.o(n18263),
	.a(n23316),
	.b(FE_OFN111_n22773));
   ao22f01 U20752 (.o(n22283),
	.a(FE_OFN111_n22773),
	.b(n23611),
	.c(n17755),
	.d(n23613));
   in01f01 U20753 (.o(n22838),
	.a(n20911));
   in01f01 U20754 (.o(n22835),
	.a(n20912));
   ao22f01 U20755 (.o(n22907),
	.a(FE_OFN94_n21695),
	.b(n18028),
	.c(FE_OFN389_n17786),
	.d(n25516));
   ao22f01 U20756 (.o(n22533),
	.a(FE_OFN389_n17786),
	.b(n23543),
	.c(n17755),
	.d(n23542));
   ao22m01 U20757 (.o(n20741),
	.a(n19054),
	.b(n23965),
	.c(n19056),
	.d(n23967));
   ao22f01 U20758 (.o(n21719),
	.a(FE_OFN111_n22773),
	.b(n23511),
	.c(n17755),
	.d(n23510));
   na02f01 U20759 (.o(n20574),
	.a(n21565),
	.b(n21431));
   ao22f01 U20760 (.o(n21723),
	.a(n17786),
	.b(n23533),
	.c(FE_OFN94_n21695),
	.d(n23532));
   ao22m01 U20761 (.o(n21738),
	.a(n17786),
	.b(n23525),
	.c(n17755),
	.d(n23524));
   ao22f01 U20762 (.o(n22526),
	.a(n19493),
	.b(n23966),
	.c(FE_OFN93_n21667),
	.d(n23967));
   ao22m01 U20763 (.o(n22527),
	.a(FE_OFN105_n22517),
	.b(n23968),
	.c(n25498),
	.d(n23965));
   ao22f01 U20764 (.o(n22221),
	.a(n17786),
	.b(n23951),
	.c(FE_OFN94_n21695),
	.d(n23950));
   ao22f01 U20765 (.o(n22230),
	.a(n17786),
	.b(n25231),
	.c(n17755),
	.d(n23957));
   ao22m01 U20766 (.o(n21731),
	.a(FE_OFN526_n24731),
	.b(n23486),
	.c(n17755),
	.d(n23488));
   ao22f01 U20767 (.o(n22510),
	.a(n19493),
	.b(n25231),
	.c(FE_OFN93_n21667),
	.d(n23957));
   ao22f01 U20768 (.o(n22501),
	.a(n19493),
	.b(n23951),
	.c(FE_OFN105_n22517),
	.d(n23950));
   ao22f01 U20769 (.o(n22234),
	.a(FE_OFN94_n21695),
	.b(n23968),
	.c(n17786),
	.d(n23966));
   ao22f01 U20770 (.o(n22233),
	.a(FE_OFN526_n24731),
	.b(n23965),
	.c(n17755),
	.d(n23967));
   ao22m01 U20771 (.o(n22302),
	.a(n19493),
	.b(n23525),
	.c(FE_OFN93_n21667),
	.d(n23524));
   ao22m01 U20772 (.o(n22299),
	.a(n19493),
	.b(n23533),
	.c(FE_OFN105_n22517),
	.d(n23532));
   ao22m01 U20773 (.o(n22436),
	.a(n19493),
	.b(n24029),
	.c(FE_OFN105_n22517),
	.d(n24028));
   ao22f01 U20774 (.o(n22506),
	.a(n19493),
	.b(n23621),
	.c(FE_OFN93_n21667),
	.d(n23620));
   oa22m01 U20775 (.o(n21492),
	.a(n23183),
	.b(n22773),
	.c(n23185),
	.d(n22772));
   ao22f01 U20776 (.o(n21729),
	.a(FE_OFN94_n21695),
	.b(n23493),
	.c(FE_OFN111_n22773),
	.d(n23492));
   ao22f01 U20777 (.o(n21711),
	.a(FE_OFN111_n22773),
	.b(n23501),
	.c(n17755),
	.d(n23500));
   no02f01 U20778 (.o(n25053),
	.a(n25052),
	.b(n25051));
   ao22f01 U20779 (.o(n21705),
	.a(FE_OFN94_n21695),
	.b(n23303),
	.c(n17786),
	.d(n23301));
   ao22m01 U20780 (.o(n21726),
	.a(n17773),
	.b(n23293),
	.c(FE_OFN526_n24731),
	.d(n23292));
   ao22f01 U20781 (.o(n21327),
	.a(FE_OFN44_n19054),
	.b(n23511),
	.c(FE_OFN47_n19056),
	.d(n23510));
   ao22m01 U20782 (.o(n21443),
	.a(n19054),
	.b(n23486),
	.c(n19056),
	.d(n23488));
   ao22f01 U20783 (.o(n21701),
	.a(FE_OFN526_n24731),
	.b(n23322),
	.c(n17755),
	.d(n23324));
   ao22f01 U20784 (.o(n20775),
	.a(n19022),
	.b(n23968),
	.c(n19019),
	.d(n23966));
   ao22s01 U20785 (.o(n21406),
	.a(n19017),
	.b(n23501),
	.c(n19020),
	.d(n23500));
   ao22f01 U20786 (.o(n23625),
	.a(FE_OFN259_n25295),
	.b(n23621),
	.c(n25294),
	.d(n23620));
   na02f06 U20787 (.o(n18389),
	.a(n19715),
	.b(n19716));
   ao12f01 U20788 (.o(n20635),
	.a(n20634),
	.b(FE_OFN24831_n25232),
	.c(n24029));
   ao22m01 U20789 (.o(n23969),
	.a(n17787),
	.b(n23968),
	.c(n25294),
	.d(n23967));
   ao22f01 U20790 (.o(n21400),
	.a(n19019),
	.b(n23621),
	.c(n19020),
	.d(n23620));
   ao22f01 U20791 (.o(n23970),
	.a(FE_OFN259_n25295),
	.b(n23966),
	.c(FE_OFN79_n20501),
	.d(n23965));
   ao22m01 U20792 (.o(n21450),
	.a(n19019),
	.b(n24029),
	.c(n19022),
	.d(n24028));
   ao22f01 U20793 (.o(n21345),
	.a(n19022),
	.b(n23303),
	.c(n19019),
	.d(n23301));
   ao22m01 U20795 (.o(n24033),
	.a(FE_OFN260_n25295),
	.b(n24029),
	.c(n17787),
	.d(n24028));
   ao22m01 U20796 (.o(n21554),
	.a(n19019),
	.b(n23533),
	.c(n19022),
	.d(n23532));
   ao22m01 U20797 (.o(n23539),
	.a(FE_OFN259_n25295),
	.b(n23533),
	.c(n17787),
	.d(n23532));
   ao22m01 U20798 (.o(n21518),
	.a(n19019),
	.b(n23525),
	.c(n19020),
	.d(n23524));
   no02s01 U20799 (.o(n20617),
	.a(n24970),
	.b(n23621));
   ao22m01 U20800 (.o(n21150),
	.a(n19022),
	.b(n23293),
	.c(n19017),
	.d(n23292));
   na02f02 U20801 (.o(n20059),
	.a(n20058),
	.b(n20057));
   ao22m01 U20802 (.o(n21130),
	.a(n19019),
	.b(n23951),
	.c(n19022),
	.d(n23950));
   ao22m01 U20803 (.o(n21428),
	.a(n19017),
	.b(n23486),
	.c(n19020),
	.d(n23488));
   ao22f01 U20804 (.o(n23485),
	.a(FE_OFN259_n25295),
	.b(n23479),
	.c(FE_OFN79_n20501),
	.d(n23478));
   ao22f01 U20805 (.o(n20966),
	.a(n19019),
	.b(n25231),
	.c(n19020),
	.d(n23957));
   ao22m01 U20806 (.o(n23531),
	.a(FE_OFN259_n25295),
	.b(n23525),
	.c(n25294),
	.d(n23524));
   in01f01 U20807 (.o(n23589),
	.a(n18459));
   ao22f01 U20808 (.o(n21377),
	.a(n19017),
	.b(n23322),
	.c(n19020),
	.d(n23324));
   ao22f01 U20809 (.o(n23961),
	.a(FE_OFN259_n25295),
	.b(n25231),
	.c(n25294),
	.d(n23957));
   ao22m01 U20810 (.o(n23952),
	.a(FE_OFN260_n25295),
	.b(n23951),
	.c(n17787),
	.d(n23950));
   na02f02 U20811 (.o(n20030),
	.a(n20026),
	.b(n20025));
   ao22m01 U20812 (.o(n22494),
	.a(FE_OFN42_n19022),
	.b(n23332),
	.c(n19019),
	.d(FE_RN_25));
   ao22f01 U20813 (.o(n21477),
	.a(n19059),
	.b(n23493),
	.c(n19054),
	.d(n23492));
   ao22f01 U20814 (.o(n23499),
	.a(n17787),
	.b(n23493),
	.c(FE_OFN79_n20501),
	.d(n23492));
   ao22f01 U20815 (.o(n21338),
	.a(FE_OFN44_n19054),
	.b(n23611),
	.c(FE_OFN47_n19056),
	.d(n23613));
   oa22m01 U20816 (.o(n22930),
	.a(n22926),
	.b(n25027),
	.c(n22925),
	.d(n20501));
   ao22f01 U20817 (.o(n21134),
	.a(n19057),
	.b(n23951),
	.c(n19059),
	.d(n23950));
   oa22f01 U20818 (.o(n21496),
	.a(n23183),
	.b(n21673),
	.c(n23185),
	.d(FE_OFN565_n25385));
   ao22m01 U20819 (.o(n25505),
	.a(FE_OFN42_n19022),
	.b(n25510),
	.c(n19019),
	.d(n21696));
   ao22f01 U20820 (.o(n21474),
	.a(n19022),
	.b(n23493),
	.c(n19017),
	.d(n23492));
   ao22f01 U20821 (.o(n23507),
	.a(FE_OFN79_n20501),
	.b(n23501),
	.c(n25294),
	.d(n23500));
   oa22m01 U20822 (.o(n23188),
	.a(n23184),
	.b(n25027),
	.c(n23183),
	.d(n20501));
   ao22f01 U20823 (.o(n21334),
	.a(FE_OFN35_n19017),
	.b(n23611),
	.c(n19020),
	.d(n23613));
   ao22m01 U20824 (.o(n20774),
	.a(n19017),
	.b(n23965),
	.c(n19020),
	.d(n23967));
   na02f10 U20825 (.o(n23500),
	.a(n19210),
	.b(n19209));
   na02f04 U20826 (.o(n23524),
	.a(n19905),
	.b(n19906));
   ao12m01 U20827 (.o(n25820),
	.a(n20487),
	.b(n20489),
	.c(n20488));
   na02f02 U20828 (.o(n23045),
	.a(n23100),
	.b(n25980));
   na03f10 U20829 (.o(n23294),
	.a(n17887),
	.b(n17886),
	.c(n17885));
   na02f06 U20830 (.o(n24031),
	.a(n19896),
	.b(n19895));
   in01f04 U20831 (.o(n18879),
	.a(n18874));
   oa22m01 U20832 (.o(n22660),
	.a(n22858),
	.b(n22773),
	.c(n22860),
	.d(n22772));
   na02f04 U20833 (.o(n23984),
	.a(n19979),
	.b(n19978));
   na02f04 U20834 (.o(n23532),
	.a(n19962),
	.b(n19961));
   na02f04 U20836 (.o(n23622),
	.a(n19966),
	.b(n19965));
   oa22s01 U20837 (.o(n21453),
	.a(n22858),
	.b(n21662),
	.c(n22860),
	.d(FE_OFN563_n25120));
   oa12s01 U20838 (.o(n20627),
	.a(n24970),
	.b(n20727),
	.c(n20626));
   ao22m01 U20839 (.o(n25822),
	.a(n25444),
	.b(n25443),
	.c(n25442),
	.d(n25441));
   oa22f01 U20840 (.o(n21456),
	.a(n22858),
	.b(n21673),
	.c(n22860),
	.d(FE_OFN565_n25385));
   na02f06 U20843 (.o(n19122),
	.a(n19093),
	.b(n19092));
   na02f04 U20844 (.o(n23518),
	.a(n19960),
	.b(n19959));
   na02f08 U20845 (.o(n23516),
	.a(n19898),
	.b(n19897));
   na02f10 U20846 (.o(n23966),
	.a(n18976),
	.b(n18975));
   na02f04 U20847 (.o(n23950),
	.a(n19968),
	.b(n19967));
   na02m02 U20848 (.o(n19985),
	.a(n19984),
	.b(n19983));
   no04f20 U20849 (.o(n22926),
	.a(n18087),
	.b(n18086),
	.c(n19000),
	.d(n18085));
   na02f10 U20850 (.o(n19003),
	.a(n18987),
	.b(n18986));
   na02s01 U20851 (.o(n25156),
	.a(n25247),
	.b(n25153));
   ao12s01 U20852 (.o(n20634),
	.a(FE_OFN24831_n25232),
	.b(n20633),
	.c(n20632));
   na02f08 U20853 (.o(n18774),
	.a(n18773),
	.b(n18772));
   in01f08 U20855 (.o(n18768),
	.a(n18764));
   oa22m01 U20856 (.o(n25821),
	.a(n25461),
	.b(n25460),
	.c(n25459),
	.d(n25458));
   no02f01 U20857 (.o(n18563),
	.a(FE_OFN24806_n19655),
	.b(n18564));
   no02f08 U20858 (.o(n18752),
	.a(n18349),
	.b(n18347));
   no02f01 U20859 (.o(n18559),
	.a(FE_OFN24806_n19655),
	.b(n18560));
   no02f02 U20860 (.o(n17848),
	.a(FE_OFN24806_n19655),
	.b(n17849));
   no02s01 U20861 (.o(n18561),
	.a(FE_OFN24806_n19655),
	.b(n18562));
   ao22f04 U20863 (.o(n19461),
	.a(n19451),
	.b(n19450),
	.c(n20514),
	.d(n21907));
   na02f02 U20864 (.o(n20971),
	.a(n20994),
	.b(n25896));
   na02f02 U20865 (.o(n21914),
	.a(n21943),
	.b(n23760));
   in01f03 U20866 (.o(n21671),
	.a(n19022));
   na02f02 U20867 (.o(n21944),
	.a(n21943),
	.b(n23736));
   na03f01 U20868 (.o(n25431),
	.a(n17888),
	.b(n19225),
	.c(n25427));
   na02f02 U20870 (.o(n23735),
	.a(n23734),
	.b(n23733));
   no02s01 U20871 (.o(n18345),
	.a(n18715),
	.b(n18346));
   na02f10 U20872 (.o(n19871),
	.a(n20422),
	.b(n20379));
   na02f10 U20873 (.o(n25027),
	.a(n25052),
	.b(n25061));
   no02s01 U20874 (.o(n25041),
	.a(n25475),
	.b(n25040));
   no02m01 U20875 (.o(n22376),
	.a(n22385),
	.b(n22392));
   in01s01 U20876 (.o(n23760),
	.a(n21913));
   no02f02 U20877 (.o(n21584),
	.a(n21151),
	.b(n20768));
   no02f10 U20878 (.o(n19056),
	.a(n25129),
	.b(n20462));
   na02f06 U20879 (.o(n24982),
	.a(n19252),
	.b(n20123));
   oa12m01 U20880 (.o(n25476),
	.a(n25474),
	.b(n25475),
	.c(n25482));
   in01f10 U20881 (.o(n18715),
	.a(FE_RN_41));
   no02f10 U20882 (.o(n20422),
	.a(n18807),
	.b(n18806));
   in01s01 U20883 (.o(n23736),
	.a(n21942));
   no02m01 U20884 (.o(n22071),
	.a(n22067),
	.b(n22082));
   in01f02 U20885 (.o(n18644),
	.a(n20970));
   no02f01 U20887 (.o(n18337),
	.a(FE_OFN24745_n18648),
	.b(n18338));
   no02f01 U20888 (.o(n18335),
	.a(FE_OFN24745_n18648),
	.b(n18336));
   na02f10 U20889 (.o(n25029),
	.a(n18790),
	.b(n25061));
   no02s01 U20890 (.o(n25131),
	.a(n25130),
	.b(n25129));
   in01m06 U20891 (.o(n19058),
	.a(n25123));
   in01f01 U20894 (.o(n22956),
	.a(n22955));
   no02f04 U20896 (.o(n25292),
	.a(n25286),
	.b(n25285));
   no02f04 U20897 (.o(n18496),
	.a(n18497),
	.b(n25420));
   no03f04 U20898 (.o(n20544),
	.a(n25184),
	.b(n25183),
	.c(n20533));
   oa22f02 U20899 (.o(n25165),
	.a(n18430),
	.b(n18427),
	.c(n25170),
	.d(n25164));
   na02f02 U20900 (.o(n18190),
	.a(n18196),
	.b(n18195));
   na02f02 U20901 (.o(n25073),
	.a(n25463),
	.b(n25149));
   na02f02 U20902 (.o(n25400),
	.a(n25399),
	.b(n25398));
   no02f04 U20903 (.o(n18280),
	.a(n18282),
	.b(n18281));
   no02f02 U20904 (.o(n18612),
	.a(n18613),
	.b(n18399));
   no02f02 U20905 (.o(n18608),
	.a(n18609),
	.b(n18399));
   in01f02 U20906 (.o(n18494),
	.a(n25034));
   oa22f02 U20907 (.o(n25341),
	.a(n25340),
	.b(n25339),
	.c(n25338),
	.d(n25337));
   na02f02 U20908 (.o(n20546),
	.a(n20554),
	.b(n25506));
   no02f04 U20909 (.o(n18636),
	.a(n18637),
	.b(n18507));
   na02f04 U20910 (.o(n25478),
	.a(n25485),
	.b(n25482));
   no02f04 U20911 (.o(n18593),
	.a(n24967),
	.b(n18399));
   no02f02 U20912 (.o(n18634),
	.a(n18635),
	.b(n18507));
   no02f06 U20913 (.o(n25034),
	.a(n18112),
	.b(n25032));
   no02f02 U20914 (.o(n24963),
	.a(n25499),
	.b(n18057));
   no03f06 U20915 (.o(n25098),
	.a(n18293),
	.b(n25094),
	.c(n18292));
   in01f02 U20916 (.o(n18282),
	.a(n20479));
   na02f04 U20917 (.o(n25338),
	.a(n25318),
	.b(n25317));
   na02f02 U20918 (.o(n18195),
	.a(n18458),
	.b(n18601));
   no02f04 U20919 (.o(n18568),
	.a(n18570),
	.b(n18569));
   na02f04 U20920 (.o(n24957),
	.a(FE_OFN25651_n25499),
	.b(n24956));
   na02f02 U20921 (.o(n25013),
	.a(n25415),
	.b(n25417));
   na02m02 U20922 (.o(n18079),
	.a(n20339),
	.b(n18080));
   na03f08 U20923 (.o(n18627),
	.a(n20344),
	.b(n24973),
	.c(n18443));
   na02f06 U20924 (.o(n20540),
	.a(n20539),
	.b(n20538));
   no02f06 U20925 (.o(n25102),
	.a(n18526),
	.b(n25090));
   in01m02 U20926 (.o(n18525),
	.a(n25389));
   na02f02 U20927 (.o(n20558),
	.a(n25065),
	.b(n20555));
   na02f02 U20928 (.o(n25337),
	.a(n25336),
	.b(n25335));
   na02f04 U20929 (.o(n19887),
	.a(FE_OFN428_n22902),
	.b(n18080));
   na02m02 U20930 (.o(n20339),
	.a(n21667),
	.b(n24968));
   in01f02 U20931 (.o(n17758),
	.a(n24974));
   no02f03 U20932 (.o(n25397),
	.a(n19019),
	.b(n20312));
   na02f04 U20933 (.o(n25082),
	.a(n25081),
	.b(n25080));
   na02f02 U20934 (.o(n25434),
	.a(validOut_W),
	.b(FE_OFN25596_reset));
   na02f08 U20935 (.o(n25124),
	.a(n18401),
	.b(n18400));
   na02f08 U20936 (.o(n18205),
	.a(n21673),
	.b(n20545));
   na02f06 U20937 (.o(n18400),
	.a(n18402),
	.b(n18403));
   in01f06 U20938 (.o(n20545),
	.a(n25387));
   in01f04 U20939 (.o(n18432),
	.a(n20384));
   na02f02 U20940 (.o(n24760),
	.a(validOut_E),
	.b(FE_OFN25599_reset));
   na02f08 U20941 (.o(n24955),
	.a(FE_OFN428_n22902),
	.b(n24954));
   no02f03 U20942 (.o(n20312),
	.a(n18215),
	.b(n18213));
   na02f02 U20943 (.o(n23558),
	.a(validOut_N),
	.b(FE_OFN25599_reset));
   no02f03 U20944 (.o(n25415),
	.a(n25300),
	.b(n25008));
   no02f04 U20945 (.o(n18404),
	.a(n20150),
	.b(n18492));
   in01f06 U20946 (.o(n18211),
	.a(n18212));
   no02f04 U20947 (.o(n20449),
	.a(n20445),
	.b(n20446));
   no02f06 U20948 (.o(n25007),
	.a(n25018),
	.b(n20268));
   oa12f02 U20949 (.o(n18213),
	.a(n18214),
	.b(n20264),
	.c(n20263));
   na02f02 U20950 (.o(n25160),
	.a(n25162),
	.b(n25159));
   in01m02 U20951 (.o(n25024),
	.a(n18542));
   ao12m02 U20952 (.o(n20262),
	.a(n21673),
	.b(n20450),
	.c(n20261));
   in01f08 U20953 (.o(n25018),
	.a(n18622));
   no02f02 U20954 (.o(n20402),
	.a(n20399),
	.b(n20398));
   no03f04 U20955 (.o(n20452),
	.a(n20442),
	.b(n20441),
	.c(n24970));
   na02f10 U20956 (.o(n20294),
	.a(n20379),
	.b(n20407));
   no02f02 U20957 (.o(n20261),
	.a(n20260),
	.b(n20263));
   na02f04 U20958 (.o(n20209),
	.a(n20207),
	.b(n20206));
   na02f06 U20959 (.o(n18379),
	.a(n20381),
	.b(n20369));
   no02f02 U20960 (.o(n19561),
	.a(n20200),
	.b(n19740));
   oa12f04 U20961 (.o(n20419),
	.a(n20282),
	.b(n20284),
	.c(n20283));
   in01s02 U20962 (.o(n20393),
	.a(n20391));
   na02f04 U20964 (.o(n24977),
	.a(n24999),
	.b(FE_OFN945_n24998));
   na02f02 U20965 (.o(n20206),
	.a(n20205),
	.b(n20204));
   no02m02 U20966 (.o(n20163),
	.a(n20162),
	.b(n20161));
   na02f01 U20967 (.o(n22321),
	.a(n25499),
	.b(FE_OFN120_n23482));
   na02f01 U20968 (.o(n21718),
	.a(FE_OFN251_n25152),
	.b(n23512));
   na02f01 U20969 (.o(n21715),
	.a(FE_OFN251_n25152),
	.b(n23344));
   na02f01 U20970 (.o(n22306),
	.a(n25499),
	.b(n25405));
   na02f01 U20971 (.o(n25522),
	.a(n25521),
	.b(n18092));
   na02f01 U20972 (.o(n22908),
	.a(FE_OFN251_n25152),
	.b(FE_RN_36));
   na02f01 U20973 (.o(n21502),
	.a(FE_OFN557_n24969),
	.b(n23189));
   na02f01 U20974 (.o(n21724),
	.a(n25152),
	.b(n23296));
   na03f10 U20975 (.o(n21892),
	.a(n17864),
	.b(n17863),
	.c(n17861));
   na02f01 U20976 (.o(n21733),
	.a(n25152),
	.b(n23520));
   na02f01 U20977 (.o(n21697),
	.a(FE_OFN251_n25152),
	.b(n18064));
   na02f01 U20978 (.o(n21703),
	.a(n25152),
	.b(n23304));
   na02f01 U20979 (.o(n21727),
	.a(n25152),
	.b(n23496));
   na02f01 U20980 (.o(n21706),
	.a(n25152),
	.b(FE_OFN120_n23482));
   in01f08 U20981 (.o(n19734),
	.a(n23304));
   na02f01 U20982 (.o(n21709),
	.a(n25152),
	.b(n23504));
   in01f10 U20983 (.o(n19648),
	.a(n23318));
   na02f01 U20984 (.o(n21700),
	.a(n25152),
	.b(n23326));
   na02f01 U20985 (.o(n21721),
	.a(n25152),
	.b(FE_OFN128_n23536));
   na02f01 U20986 (.o(n21494),
	.a(n25152),
	.b(n23189));
   na02f01 U20987 (.o(n21730),
	.a(n25152),
	.b(n25405));
   na02f01 U20988 (.o(n21712),
	.a(FE_OFN251_n25152),
	.b(n23318));
   na02f01 U20989 (.o(n22300),
	.a(FE_OFN24826_n25499),
	.b(n23528));
   na02f02 U20990 (.o(n22297),
	.a(FE_OFN24826_n25499),
	.b(FE_OFN128_n23536));
   na02f01 U20991 (.o(n21736),
	.a(n25152),
	.b(n23528));
   na02f01 U20992 (.o(n21525),
	.a(n25152),
	.b(n22931));
   na02f01 U20993 (.o(n21392),
	.a(n25521),
	.b(n23326));
   na02f01 U20994 (.o(n23529),
	.a(n25301),
	.b(n23528));
   na02f01 U20995 (.o(n21442),
	.a(n25521),
	.b(n25405));
   ao22f01 U20996 (.o(n21590),
	.a(FE_OFN24831_n25232),
	.b(n21539),
	.c(n21538),
	.d(n21537));
   na02f01 U20998 (.o(n23537),
	.a(n25301),
	.b(FE_OFN128_n23536));
   oa12m02 U20999 (.o(n20161),
	.a(n20170),
	.b(n20160),
	.c(n20159));
   na02f01 U21000 (.o(n21346),
	.a(n25521),
	.b(n23304));
   na02f01 U21001 (.o(n23513),
	.a(FE_OFN262_n25301),
	.b(n23512));
   no03m02 U21002 (.o(n20162),
	.a(n20157),
	.b(n20156),
	.c(n20166));
   na02f01 U21003 (.o(n21412),
	.a(n25521),
	.b(n23504));
   na02f01 U21004 (.o(n21498),
	.a(n25506),
	.b(n23189));
   na02f01 U21005 (.o(n21555),
	.a(n25521),
	.b(FE_OFN128_n23536));
   na02f01 U21006 (.o(n21529),
	.a(n25506),
	.b(n22931));
   na02f01 U21007 (.o(n21475),
	.a(n25521),
	.b(n23496));
   na02f01 U21008 (.o(n25513),
	.a(n25521),
	.b(n18064));
   na02f01 U21009 (.o(n21296),
	.a(FE_OFN269_n25506),
	.b(n23512));
   no02f02 U21010 (.o(n20307),
	.a(n20392),
	.b(n20298));
   na02f01 U21011 (.o(n22294),
	.a(FE_OFN24830_n25499),
	.b(n23512));
   na02f01 U21012 (.o(n22932),
	.a(n25301),
	.b(n22931));
   na02f01 U21013 (.o(n23190),
	.a(n25301),
	.b(n23189));
   na02f01 U21014 (.o(n23497),
	.a(n25301),
	.b(n23496));
   na02f01 U21015 (.o(n23505),
	.a(n25301),
	.b(n23504));
   na02f01 U21016 (.o(n23305),
	.a(n25301),
	.b(n23304));
   na02f01 U21017 (.o(n21552),
	.a(FE_OFN269_n25506),
	.b(FE_OFN128_n23536));
   na02f01 U21018 (.o(n23297),
	.a(n25301),
	.b(n23296));
   na02f01 U21019 (.o(n23327),
	.a(n25301),
	.b(n23326));
   na02f01 U21020 (.o(n21516),
	.a(FE_OFN269_n25506),
	.b(n23528));
   na02f01 U21021 (.o(n21466),
	.a(n25521),
	.b(FE_RN_36));
   na02f01 U21022 (.o(n21559),
	.a(FE_OFN269_n25506),
	.b(n23520));
   na02f01 U21023 (.o(n23345),
	.a(FE_OFN262_n25301),
	.b(n23344));
   na02f01 U21024 (.o(n23337),
	.a(FE_OFN262_n25301),
	.b(n18064));
   na02f01 U21025 (.o(n21439),
	.a(n25521),
	.b(n23296));
   na02f01 U21026 (.o(n23334),
	.a(FE_OFN262_n25301),
	.b(FE_RN_36));
   in01f01 U21028 (.o(n21649),
	.a(n23528));
   na02f01 U21029 (.o(n23489),
	.a(n25301),
	.b(n25405));
   na02f01 U21030 (.o(n23319),
	.a(FE_OFN262_n25301),
	.b(n23318));
   na02f01 U21031 (.o(n21459),
	.a(n25506),
	.b(FE_OFN120_n23482));
   na02f01 U21033 (.o(n23483),
	.a(n25301),
	.b(FE_OFN120_n23482));
   na02f01 U21034 (.o(n21427),
	.a(n25506),
	.b(n25405));
   na02f01 U21035 (.o(n21462),
	.a(n25521),
	.b(FE_OFN120_n23482));
   na02f01 U21036 (.o(n23521),
	.a(n25301),
	.b(n23520));
   no02m02 U21037 (.o(n20435),
	.a(n20432),
	.b(n20431));
   no02f02 U21038 (.o(n20330),
	.a(n21667),
	.b(n19955));
   no02f10 U21039 (.o(n19048),
	.a(n19040),
	.b(n19039));
   na02f01 U21040 (.o(n22287),
	.a(FE_OFN24830_n25499),
	.b(n23344));
   na02f01 U21041 (.o(n21148),
	.a(n25506),
	.b(n23296));
   na02f01 U21042 (.o(n21376),
	.a(n25506),
	.b(n23326));
   na02f01 U21043 (.o(n21486),
	.a(FE_OFN269_n25506),
	.b(n23318));
   na02f01 U21044 (.o(n22327),
	.a(FE_OFN24830_n25499),
	.b(n18064));
   na02f01 U21045 (.o(n21343),
	.a(n25506),
	.b(n23304));
   na02f01 U21046 (.o(n21519),
	.a(n25521),
	.b(n23528));
   na02f01 U21047 (.o(n22309),
	.a(FE_OFN24830_n25499),
	.b(FE_RN_36));
   na02f01 U21048 (.o(n21404),
	.a(n25506),
	.b(n23504));
   na02f01 U21049 (.o(n22330),
	.a(FE_OFN559_n24969),
	.b(n23326));
   na02f01 U21050 (.o(n21489),
	.a(n25521),
	.b(n23318));
   na02f01 U21051 (.o(n21562),
	.a(n25521),
	.b(n23520));
   na02f01 U21052 (.o(n22318),
	.a(FE_OFN558_n24969),
	.b(n23296));
   na02f01 U21053 (.o(n25507),
	.a(FE_OFN269_n25506),
	.b(n18093));
   na02f01 U21054 (.o(n21329),
	.a(n25521),
	.b(n23344));
   na02f01 U21055 (.o(n22303),
	.a(FE_OFN24827_n25499),
	.b(n23304));
   na02f01 U21056 (.o(n21543),
	.a(n25521),
	.b(n22931));
   na02f01 U21057 (.o(n22315),
	.a(FE_OFN24830_n25499),
	.b(n23318));
   na02f01 U21058 (.o(n22492),
	.a(FE_OFN269_n25506),
	.b(FE_RN_36));
   na02f01 U21059 (.o(n21290),
	.a(FE_OFN269_n25506),
	.b(n23344));
   na02f01 U21060 (.o(n22290),
	.a(FE_OFN24828_n25499),
	.b(n23504));
   na02f01 U21061 (.o(n25503),
	.a(FE_OFN269_n25506),
	.b(n18064));
   na02f01 U21062 (.o(n22312),
	.a(FE_OFN24825_n25499),
	.b(n23496));
   na02f01 U21063 (.o(n21506),
	.a(n25521),
	.b(n23189));
   na02f01 U21064 (.o(n21472),
	.a(n25506),
	.b(n23496));
   na02f01 U21065 (.o(n21326),
	.a(n25521),
	.b(n23512));
   na02f01 U21066 (.o(n21533),
	.a(FE_RN_18_0),
	.b(n22931));
   in01f01 U21067 (.o(n18030),
	.a(FE_RN_21));
   no02f08 U21068 (.o(n19131),
	.a(n19120),
	.b(n20153));
   na03f10 U21069 (.o(n20429),
	.a(n20430),
	.b(n18965),
	.c(n20433));
   na02f10 U21070 (.o(n25405),
	.a(n19757),
	.b(n19756));
   na02f08 U21071 (.o(n25520),
	.a(n19620),
	.b(n19621));
   in01f04 U21072 (.o(n18463),
	.a(n18464));
   in01m01 U21073 (.o(n19850),
	.a(n19848));
   ao22f01 U21074 (.o(n25248),
	.a(n25247),
	.b(n25246),
	.c(n25245),
	.d(n25244));
   na03f02 U21075 (.o(n20295),
	.a(n23035),
	.b(n20408),
	.c(n20293));
   no02f02 U21076 (.o(n20404),
	.a(n20303),
	.b(n20302));
   na02f06 U21077 (.o(n20104),
	.a(n23964),
	.b(n24036));
   no02f04 U21078 (.o(n21908),
	.a(n19949),
	.b(n19948));
   oa12f08 U21079 (.o(n20352),
	.a(n19976),
	.b(n25246),
	.c(n19977));
   no02f08 U21080 (.o(n23628),
	.a(n20082),
	.b(n20081));
   in01f06 U21081 (.o(n19125),
	.a(n19124));
   no02f06 U21082 (.o(n19757),
	.a(n19749),
	.b(n19748));
   in01f06 U21083 (.o(n17855),
	.a(n18508));
   in01f06 U21084 (.o(n17854),
	.a(n18515));
   no02f08 U21085 (.o(n17852),
	.a(n19699),
	.b(n19694));
   oa12f04 U21086 (.o(n19463),
	.a(n20350),
	.b(n19871),
	.c(n19479));
   in01s01 U21087 (.o(n18596),
	.a(n22939));
   no02f03 U21089 (.o(n24009),
	.a(n21509),
	.b(n21508));
   no02f08 U21090 (.o(n18367),
	.a(n18371),
	.b(n18368));
   in01f01 U21091 (.o(n20927),
	.a(n20926));
   na02f06 U21092 (.o(n25246),
	.a(n19972),
	.b(n19971));
   na02f02 U21093 (.o(n19948),
	.a(n19947),
	.b(n19946));
   in01f01 U21094 (.o(n19786),
	.a(n20242));
   no02f06 U21095 (.o(n18020),
	.a(n19347),
	.b(n18226));
   in01f01 U21096 (.o(n25497),
	.a(n22904));
   in01f04 U21097 (.o(n19629),
	.a(n18029));
   no02f06 U21098 (.o(n19756),
	.a(n19755),
	.b(n19754));
   no03f10 U21099 (.o(n17995),
	.a(n17999),
	.b(n17998),
	.c(n17996));
   in01s01 U21100 (.o(n20401),
	.a(n20400));
   in01f01 U21101 (.o(n23502),
	.a(n21403));
   in01f01 U21102 (.o(n22760),
	.a(n23995));
   na02s01 U21103 (.o(n21644),
	.a(n21647),
	.b(n21643));
   in01f06 U21104 (.o(n22829),
	.a(n19122));
   in01f01 U21105 (.o(n22761),
	.a(n23994));
   na02s01 U21107 (.o(n18457),
	.a(FE_OFN428_n22902),
	.b(n25130));
   in01f06 U21108 (.o(n18094),
	.a(n19660));
   in01f01 U21109 (.o(n22753),
	.a(n24003));
   in01f01 U21110 (.o(n22867),
	.a(FE_RN_44));
   na02f08 U21111 (.o(n17817),
	.a(n18321),
	.b(n18318));
   ao22m01 U21112 (.o(n22222),
	.a(n17755),
	.b(n23949),
	.c(FE_OFN111_n22773),
	.d(FE_OFN138_n23948));
   no03f06 U21113 (.o(n19909),
	.a(n24031),
	.b(n23516),
	.c(n23949));
   no02f04 U21114 (.o(n20564),
	.a(n22912),
	.b(n23983));
   no04f08 U21115 (.o(n19971),
	.a(n23958),
	.b(n23622),
	.c(n23950),
	.d(n24028));
   no03f06 U21116 (.o(n19972),
	.a(n23526),
	.b(n23518),
	.c(n23532));
   in01f01 U21117 (.o(n22892),
	.a(n21407));
   no02f04 U21118 (.o(n20001),
	.a(n25231),
	.b(n24029));
   no02f04 U21119 (.o(n19991),
	.a(n23533),
	.b(n23525));
   ao22m01 U21120 (.o(n22502),
	.a(n25498),
	.b(FE_OFN138_n23948),
	.c(FE_OFN93_n21667),
	.d(n23949));
   no02m02 U21121 (.o(n19946),
	.a(n23959),
	.b(n23623));
   in01f01 U21122 (.o(n22852),
	.a(n20759));
   na04f10 U21123 (.o(n19540),
	.a(n19534),
	.b(n19533),
	.c(n19532),
	.d(n19531));
   in01f01 U21124 (.o(n22883),
	.a(n21141));
   ao22m01 U21125 (.o(n25524),
	.a(n17753),
	.b(n18028),
	.c(n19057),
	.d(n25516));
   in01f02 U21126 (.o(n22876),
	.a(n20784));
   in01f01 U21127 (.o(n21615),
	.a(n23586));
   in01f01 U21128 (.o(n23541),
	.a(n20745));
   na04f20 U21130 (.o(n18235),
	.a(n18413),
	.b(n18414),
	.c(n18412),
	.d(n18415));
   in01f01 U21131 (.o(n22752),
	.a(n24004));
   no02f02 U21132 (.o(n22868),
	.a(n20644),
	.b(n20643));
   na02f08 U21133 (.o(n17942),
	.a(n17944),
	.b(n17943));
   in01f01 U21134 (.o(n21471),
	.a(n21470));
   in01s01 U21135 (.o(n21293),
	.a(n23509));
   in01f01 U21136 (.o(n21333),
	.a(FE_RN_68));
   no02f04 U21137 (.o(n19953),
	.a(FE_OFN100_n21907),
	.b(n21431));
   na03f10 U21139 (.o(n17892),
	.a(n17895),
	.b(n17894),
	.c(n17893));
   in01f02 U21140 (.o(n22891),
	.a(n21408));
   na04s02 U21141 (.o(n25239),
	.a(n25238),
	.b(FE_OFN253_n25241),
	.c(n25240),
	.d(n25237));
   na02f01 U21142 (.o(n20753),
	.a(n25247),
	.b(n23622));
   no02m02 U21143 (.o(n19947),
	.a(n23948),
	.b(n24030));
   na02f01 U21144 (.o(n20640),
	.a(n25247),
	.b(n24028));
   na02f01 U21145 (.o(n23311),
	.a(n25247),
	.b(n23526));
   na02s01 U21146 (.o(n18266),
	.a(n23317),
	.b(n19493));
   na02f01 U21147 (.o(n20730),
	.a(FE_OFN24831_n25232),
	.b(n23525));
   in01f04 U21148 (.o(n19231),
	.a(n23494));
   no03f20 U21149 (.o(n22861),
	.a(n18769),
	.b(n18768),
	.c(n18767));
   no03f10 U21150 (.o(n20400),
	.a(n19229),
	.b(n19228),
	.c(n20302));
   na02s01 U21151 (.o(n20654),
	.a(n21893),
	.b(n23535));
   na02f01 U21152 (.o(n23043),
	.a(FE_OFN24831_n25232),
	.b(n23951));
   no03f10 U21153 (.o(n19817),
	.a(n19441),
	.b(n19810),
	.c(n19440));
   na02m02 U21154 (.o(n20292),
	.a(n21893),
	.b(n23488));
   na02f08 U21155 (.o(n17834),
	.a(n17836),
	.b(n17835));
   in01s01 U21156 (.o(n21161),
	.a(n21160));
   na02s06 U21157 (.o(n20107),
	.a(n19257),
	.b(n23710));
   na02f01 U21158 (.o(n20628),
	.a(FE_OFN24831_n25232),
	.b(n23533));
   na03f10 U21159 (.o(n23295),
	.a(n18879),
	.b(n18878),
	.c(n18877));
   in01f04 U21160 (.o(n19133),
	.a(n18171));
   na02f10 U21161 (.o(n20528),
	.a(n19461),
	.b(n25494));
   no02f08 U21162 (.o(n19118),
	.a(FE_OFN67_n19548),
	.b(n23967));
   no02f03 U21163 (.o(n21558),
	.a(n19986),
	.b(n19985));
   na02f04 U21164 (.o(n19699),
	.a(n19698),
	.b(n19697));
   ao22f08 U21165 (.o(n19181),
	.a(n19347),
	.b(n21408),
	.c(FE_OFN73_n19631),
	.d(n19188));
   ao22m01 U21166 (.o(n21155),
	.a(n21565),
	.b(n23948),
	.c(FE_OFN575_n25463),
	.d(n21904));
   na02f04 U21167 (.o(n19694),
	.a(n19690),
	.b(n19689));
   na02f06 U21168 (.o(n17981),
	.a(n17983),
	.b(n17982));
   no03f20 U21169 (.o(n22822),
	.a(n18761),
	.b(n18760),
	.c(n18759));
   ao22m01 U21170 (.o(n21449),
	.a(n19017),
	.b(n24030),
	.c(n19020),
	.d(n24031));
   in01f08 U21171 (.o(n18881),
	.a(n22859));
   in01f01 U21173 (.o(n23487),
	.a(n21426));
   ao22f01 U21174 (.o(n21131),
	.a(n19017),
	.b(FE_OFN138_n23948),
	.c(n19020),
	.d(n23949));
   na02f08 U21175 (.o(n18829),
	.a(n19708),
	.b(n21470));
   na02f02 U21176 (.o(n19748),
	.a(n19747),
	.b(n19746));
   na02s01 U21177 (.o(n23712),
	.a(n23711),
	.b(n23710));
   ao22f01 U21178 (.o(n20965),
	.a(n19017),
	.b(FE_OFN140_n23959),
	.c(n19022),
	.d(n23958));
   na04f04 U21179 (.o(n20082),
	.a(n20076),
	.b(n20075),
	.c(n20074),
	.d(n20073));
   ao22m01 U21180 (.o(n21430),
	.a(n19019),
	.b(n23984),
	.c(n19022),
	.d(n23983));
   na02f04 U21181 (.o(n18515),
	.a(n18517),
	.b(n18516));
   ao22m01 U21182 (.o(n23953),
	.a(n25294),
	.b(n23949),
	.c(FE_OFN79_n20501),
	.d(FE_OFN138_n23948));
   na04f06 U21183 (.o(n20081),
	.a(n20080),
	.b(n20079),
	.c(n20078),
	.d(n20077));
   in01f02 U21184 (.o(n23034),
	.a(n20238));
   no04f08 U21185 (.o(n19082),
	.a(n19136),
	.b(n19135),
	.c(FE_OFN65_n19542),
	.d(n19134));
   no04f08 U21186 (.o(n19083),
	.a(n19140),
	.b(n19139),
	.c(n19138),
	.d(n19518));
   na02f10 U21187 (.o(n20759),
	.a(n18985),
	.b(n18984));
   na02f20 U21188 (.o(n23316),
	.a(n19396),
	.b(n19395));
   na02f10 U21189 (.o(n23303),
	.a(n18747),
	.b(n18746));
   na02f10 U21190 (.o(n19421),
	.a(n19320),
	.b(n19319));
   na02f20 U21191 (.o(n23509),
	.a(n18650),
	.b(n18649));
   na02f02 U21192 (.o(n23737),
	.a(n23736),
	.b(n23788));
   na02f04 U21194 (.o(n23761),
	.a(n23760),
	.b(n23788));
   na02f02 U21195 (.o(n23543),
	.a(n20747),
	.b(n20746));
   na02m01 U21196 (.o(n23631),
	.a(n19154),
	.b(n19153));
   in01f01 U21197 (.o(n20644),
	.a(n20642));
   in01f01 U21198 (.o(n23492),
	.a(n21469));
   na02f04 U21199 (.o(n23089),
	.a(n23100),
	.b(n25976));
   na02f04 U21200 (.o(n21470),
	.a(n18835),
	.b(n18842));
   na02f20 U21201 (.o(n19394),
	.a(n19393),
	.b(n19392));
   na02f04 U21202 (.o(n23959),
	.a(n19943),
	.b(n19942));
   na02f10 U21203 (.o(n23494),
	.a(n19207),
	.b(n19206));
   na02f04 U21204 (.o(n23739),
	.a(n25980),
	.b(n23788));
   na02f04 U21205 (.o(n20238),
	.a(n19308),
	.b(n19307));
   no02m01 U21207 (.o(n25825),
	.a(n22073),
	.b(n22072));
   no02s01 U21208 (.o(n18610),
	.a(FE_OFN5_reset),
	.b(n18611));
   na02f10 U21209 (.o(n23967),
	.a(n19096),
	.b(n19095));
   na02f04 U21210 (.o(n23948),
	.a(n19939),
	.b(n19938));
   no03f20 U21211 (.o(n22875),
	.a(n18983),
	.b(n18982),
	.c(n18981));
   na02f10 U21212 (.o(n23293),
	.a(n18753),
	.b(n18752));
   na02f10 U21213 (.o(n18927),
	.a(n18916),
	.b(n18915));
   na02f06 U21214 (.o(n23983),
	.a(n19975),
	.b(n19974));
   no02f10 U21216 (.o(n22851),
	.a(n19426),
	.b(n19425));
   no02f10 U21217 (.o(n22836),
	.a(n18973),
	.b(n18972));
   no02f10 U21218 (.o(n22860),
	.a(n19227),
	.b(n19226));
   no02s01 U21219 (.o(n20487),
	.a(n20494),
	.b(n20486));
   no02f10 U21220 (.o(n23183),
	.a(n19438),
	.b(n19437));
   no02f10 U21221 (.o(n22858),
	.a(n19293),
	.b(n19292));
   na02s01 U21222 (.o(n18129),
	.a(n18406),
	.b(n25978));
   no03f20 U21225 (.o(n23540),
	.a(n19385),
	.b(n19384),
	.c(n19383));
   oa12f06 U21226 (.o(n18874),
	.a(n18865),
	.b(n18866),
	.c(FE_OCPN25809_n18959));
   no02f08 U21227 (.o(n19237),
	.a(n19218),
	.b(n19217));
   no02f04 U21228 (.o(n25002),
	.a(n19305),
	.b(n19304));
   in01f01 U21231 (.o(n23301),
	.a(n21342));
   na02m01 U21232 (.o(n21900),
	.a(n21151),
	.b(FE_OFN100_n21907));
   no02f10 U21234 (.o(n19017),
	.a(n20318),
	.b(n19016));
   in01s01 U21235 (.o(n25133),
	.a(n25127));
   na02f02 U21237 (.o(n25481),
	.a(n25979),
	.b(n25473));
   na02f10 U21238 (.o(n22772),
	.a(n25163),
	.b(n20531));
   in01s01 U21239 (.o(n22272),
	.a(n22270));
   in01f20 U21240 (.o(n17782),
	.a(n18715));
   in01s01 U21242 (.o(n17784),
	.a(n25235));
   na02m01 U21245 (.o(n21687),
	.a(n21683),
	.b(n22898));
   in01f10 U21246 (.o(n17789),
	.a(n25072));
   ao22f20 U21249 (.o(n18673),
	.a(n21806),
	.b(south_input_NIB_storage_data_f_2__51_),
	.c(FE_RN_63),
	.d(south_input_NIB_storage_data_f_1__51_));
   no02f04 U21250 (.o(n18278),
	.a(n18218),
	.b(n17889));
   ao22f20 U21251 (.o(n18671),
	.a(n21806),
	.b(south_input_NIB_storage_data_f_2__53_),
	.c(n17756),
	.d(south_input_NIB_storage_data_f_1__53_));
   no02f08 U21252 (.o(n17792),
	.a(n17794),
	.b(n17793));
   na02f10 U21253 (.o(n17793),
	.a(n20118),
	.b(n20114));
   na03f40 U21254 (.o(n18377),
	.a(n17796),
	.b(n19671),
	.c(n17795));
   no04f40 U21255 (.o(n17795),
	.a(n19625),
	.b(n19624),
	.c(n19651),
	.d(n19650));
   no04f40 U21256 (.o(n17796),
	.a(n19652),
	.b(n19649),
	.c(n19627),
	.d(n19626));
   na02f08 U21257 (.o(n18288),
	.a(n18314),
	.b(n18317));
   na02f08 U21258 (.o(n18290),
	.a(n18319),
	.b(n18323));
   ao22f10 U21259 (.o(n19166),
	.a(FE_RN_10),
	.b(north_input_NIB_storage_data_f_3__56_),
	.c(FE_OFN24773_n19075),
	.d(north_input_NIB_storage_data_f_0__56_));
   ao22f04 U21260 (.o(n19640),
	.a(FE_OFN25681_n17814),
	.b(proc_input_NIB_storage_data_f_9__52_),
	.c(FE_OFN170_n24343),
	.d(proc_input_NIB_storage_data_f_8__52_));
   na02f10 U21261 (.o(n25517),
	.a(n18653),
	.b(n18652));
   no02f02 U21263 (.o(n20473),
	.a(n22902),
	.b(n20472));
   na02f06 U21264 (.o(n18210),
	.a(n18466),
	.b(n18211));
   ao22f08 U21266 (.o(n19189),
	.a(FE_RN_10),
	.b(north_input_NIB_storage_data_f_3__63_),
	.c(FE_OFN24773_n19075),
	.d(north_input_NIB_storage_data_f_0__63_));
   ao22f10 U21267 (.o(n18255),
	.a(FE_OFN24773_n19075),
	.b(north_input_NIB_storage_data_f_0__59_),
	.c(FE_RN_10),
	.d(north_input_NIB_storage_data_f_3__59_));
   na02f20 U21269 (.o(n18664),
	.a(n18060),
	.b(south_input_NIB_storage_data_f_1__55_));
   ao22f20 U21270 (.o(n18941),
	.a(n23612),
	.b(n19635),
	.c(myChipID_f_6_),
	.d(n17797));
   ao22f20 U21271 (.o(n18585),
	.a(FE_RN_63),
	.b(south_input_NIB_storage_data_f_1__54_),
	.c(n24473),
	.d(south_input_NIB_storage_data_f_3__54_));
   oa12f40 U21272 (.o(n18932),
	.a(n18930),
	.b(n18931),
	.c(FE_OCPN25807_n18959));
   oa22f02 U21274 (.o(n25420),
	.a(n25419),
	.b(n25418),
	.c(n25417),
	.d(n25416));
   na02f04 U21275 (.o(n19470),
	.a(n19467),
	.b(n18113));
   ao22f20 U21276 (.o(n18887),
	.a(FE_RN_66),
	.b(west_input_NIB_storage_data_f_0__53_),
	.c(n18828),
	.d(west_input_NIB_storage_data_f_1__53_));
   no03f20 U21277 (.o(n26019),
	.a(n17799),
	.b(n19464),
	.c(n17798));
   no03f10 U21278 (.o(n17798),
	.a(n19444),
	.b(n19475),
	.c(n19477));
   no03f10 U21279 (.o(n17799),
	.a(n19415),
	.b(n19444),
	.c(n19475));
   na02f10 U21281 (.o(n19338),
	.a(FE_OFN24780_n19932),
	.b(east_input_NIB_storage_data_f_0__62_));
   ao22f03 U21282 (.o(n19552),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__34_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__34_));
   ao22f08 U21283 (.o(n19577),
	.a(proc_input_NIB_storage_data_f_11__61_),
	.b(FE_OFN25673_n18033),
	.c(n17754),
	.d(proc_input_NIB_storage_data_f_3__61_));
   ao22f08 U21284 (.o(n19180),
	.a(FE_OFN96_n21865),
	.b(north_input_NIB_storage_data_f_2__57_),
	.c(FE_OFN25610_n19071),
	.d(north_input_NIB_storage_data_f_1__57_));
   na02f08 U21285 (.o(n20230),
	.a(n19882),
	.b(n19008));
   na02f10 U21286 (.o(n19007),
	.a(n19006),
	.b(n19005));
   na03f20 U21289 (.o(n18399),
	.a(n18544),
	.b(n17801),
	.c(n17800));
   no02f08 U21290 (.o(n17801),
	.a(n26015),
	.b(n26024));
   na02f04 U21291 (.o(n20134),
	.a(n25381),
	.b(n18507));
   no02f04 U21292 (.o(n19484),
	.a(n18615),
	.b(n19483));
   ao22f10 U21293 (.o(n18672),
	.a(south_input_NIB_storage_data_f_3__53_),
	.b(n24473),
	.c(south_input_NIB_storage_data_f_0__53_),
	.d(FE_RN_62));
   in01f10 U21295 (.o(n21660),
	.a(n18120));
   no02f20 U21296 (.o(n20529),
	.a(n20427),
	.b(n18394));
   no02f20 U21297 (.o(n20427),
	.a(n18074),
	.b(n20512));
   ao22f06 U21298 (.o(n18363),
	.a(proc_input_NIB_storage_data_f_15__43_),
	.b(FE_RN_50),
	.c(proc_input_NIB_storage_data_f_5__43_),
	.d(FE_RN_49));
   na04f10 U21299 (.o(n18359),
	.a(n18363),
	.b(n18362),
	.c(n18361),
	.d(n18360));
   no04f06 U21301 (.o(n25187),
	.a(n25184),
	.b(n25183),
	.c(n25182),
	.d(n25181));
   in01f06 U21302 (.o(n19732),
	.a(n23496));
   in01f02 U21304 (.o(n19492),
	.a(n19484));
   no02f06 U21305 (.o(n20432),
	.a(n18869),
	.b(n18880));
   no03f20 U21306 (.o(n19051),
	.a(n19035),
	.b(n19034),
	.c(north_output_control_planned_f));
   na02f20 U21307 (.o(n18531),
	.a(n19591),
	.b(n19592));
   no02f20 U21308 (.o(n18384),
	.a(n18531),
	.b(n18530));
   ao22f06 U21310 (.o(n19663),
	.a(FE_OFN25602_n19530),
	.b(proc_input_NIB_storage_data_f_13__53_),
	.c(FE_RN_19),
	.d(proc_input_NIB_storage_data_f_8__53_));
   na02f10 U21311 (.o(n18312),
	.a(n19659),
	.b(n19663));
   no02f10 U21312 (.o(n19785),
	.a(n17805),
	.b(n17802));
   ao22f10 U21314 (.o(n19602),
	.a(FE_OCPN25960_n18039),
	.b(proc_input_NIB_storage_data_f_10__63_),
	.c(FE_RN_49),
	.d(proc_input_NIB_storage_data_f_5__63_));
   no02f20 U21315 (.o(n18039),
	.a(n25140),
	.b(FE_RN_37));
   in01f08 U21316 (.o(n19466),
	.a(n17806));
   na02f10 U21317 (.o(n17806),
	.a(FE_OFN959_n25972),
	.b(n19465));
   ao22f20 U21318 (.o(n18175),
	.a(n18828),
	.b(west_input_NIB_storage_data_f_1__58_),
	.c(FE_OFN26_n18974),
	.d(west_input_NIB_storage_data_f_0__58_));
   oa12m02 U21319 (.o(n2688),
	.a(n18504),
	.b(n25076),
	.c(n18507));
   in01f04 U21320 (.o(n24979),
	.a(n20342));
   na02f08 U21321 (.o(n18514),
	.a(proc_input_NIB_storage_data_f_10__45_),
	.b(FE_OCPN25954_n18039));
   no03f10 U21322 (.o(n20127),
	.a(n26014),
	.b(n26021),
	.c(n25994));
   na02f10 U21323 (.o(n20387),
	.a(n20300),
	.b(n20390));
   no03f40 U21324 (.o(n23992),
	.a(n19353),
	.b(n19352),
	.c(n19351));
   na02f20 U21326 (.o(n18015),
	.a(n18558),
	.b(FE_OFN25609_n18377));
   na03f20 U21327 (.o(n17940),
	.a(n18378),
	.b(n20222),
	.c(n17811));
   no02f04 U21328 (.o(n18554),
	.a(n18555),
	.b(FE_OFN25609_n18377));
   no02f04 U21329 (.o(n18552),
	.a(n18553),
	.b(FE_OFN25609_n18377));
   no03m02 U21331 (.o(n20470),
	.a(n17812),
	.b(n17936),
	.c(n20462));
   no03f08 U21332 (.o(n17812),
	.a(n17831),
	.b(n17830),
	.c(n18223));
   no02f10 U21333 (.o(n20450),
	.a(n19865),
	.b(n17813));
   no02f20 U21335 (.o(n17814),
	.a(n17934),
	.b(FE_RN_37));
   na03f20 U21336 (.o(n22931),
	.a(n17818),
	.b(n17816),
	.c(n17815));
   no02f10 U21337 (.o(n17816),
	.a(n18289),
	.b(n17817));
   no02f10 U21338 (.o(n17818),
	.a(n18290),
	.b(n18288));
   no02f10 U21339 (.o(n17824),
	.a(n17826),
	.b(n17825));
   na02f10 U21340 (.o(n17825),
	.a(n19511),
	.b(n19510));
   no02f04 U21341 (.o(n20113),
	.a(n20112),
	.b(n24990));
   oa12f20 U21342 (.o(n19162),
	.a(n19160),
	.b(n19161),
	.c(n19225));
   no03f40 U21343 (.o(n19165),
	.a(n19164),
	.b(n19163),
	.c(n19162));
   na02f10 U21344 (.o(n19562),
	.a(myLocY_f_5_),
	.b(n22857));
   na02f06 U21345 (.o(n17828),
	.a(n20450),
	.b(n20195));
   na02f02 U21346 (.o(n18455),
	.a(n18456),
	.b(n17832));
   na02f08 U21347 (.o(n18274),
	.a(n25097),
	.b(n17832));
   ao12f04 U21348 (.o(n18218),
	.a(n25106),
	.b(FE_OFN428_n22902),
	.c(n17832));
   na03f10 U21349 (.o(n17832),
	.a(n18220),
	.b(n18219),
	.c(n18221));
   na03f20 U21350 (.o(n23326),
	.a(n17842),
	.b(n17839),
	.c(n17833));
   no02f10 U21351 (.o(n17833),
	.a(n17837),
	.b(n17834));
   no02f10 U21352 (.o(n17842),
	.a(n17846),
	.b(n17843));
   ao12f06 U21354 (.o(n19678),
	.a(n17848),
	.b(FE_OFN156_n24129),
	.c(proc_input_NIB_storage_data_f_1__49_));
   ao12f01 U21356 (.o(n24456),
	.a(n17850),
	.b(FE_OFN25680_n17814),
	.c(proc_input_NIB_storage_data_f_9__16_));
   no02f01 U21357 (.o(n17850),
	.a(FE_OFN24806_n19655),
	.b(n17851));
   in01s01 U21358 (.o(n17851),
	.a(proc_input_NIB_storage_data_f_3__16_));
   ao22f02 U21359 (.o(n19772),
	.a(proc_input_NIB_storage_data_f_9__30_),
	.b(n20012),
	.c(proc_input_NIB_storage_data_f_3__30_),
	.d(n19709));
   no02f10 U21360 (.o(n18025),
	.a(n18059),
	.b(n19721));
   no02f10 U21361 (.o(n19721),
	.a(n19720),
	.b(n23296));
   na02f10 U21362 (.o(n23296),
	.a(n17853),
	.b(n17852));
   na03f20 U21363 (.o(n23304),
	.a(n17856),
	.b(n17855),
	.c(n17854));
   no02f10 U21364 (.o(n17856),
	.a(n18511),
	.b(n18518));
   oa12f02 U21365 (.o(n2583),
	.a(n17857),
	.b(n20333),
	.c(n25429));
   na02f06 U21366 (.o(n17857),
	.a(n20333),
	.b(n26010));
   no02f10 U21367 (.o(n26010),
	.a(n25432),
	.b(FE_OFN25600_reset));
   na02f08 U21368 (.o(n25429),
	.a(FE_OFN25596_reset),
	.b(n25432));
   no02f20 U21369 (.o(n25432),
	.a(n17860),
	.b(n17858));
   no02f08 U21370 (.o(n17859),
	.a(n26028),
	.b(n26018));
   no03f10 U21371 (.o(n26018),
	.a(n20529),
	.b(n22772),
	.c(n20528));
   oa12f10 U21372 (.o(n22216),
	.a(n18109),
	.b(n20570),
	.c(n21892));
   in01f06 U21373 (.o(n20474),
	.a(n17867));
   na02f08 U21374 (.o(n17867),
	.a(n18377),
	.b(n17774));
   na02f08 U21375 (.o(n17868),
	.a(n18377),
	.b(n17869));
   na02f10 U21376 (.o(n24968),
	.a(n18305),
	.b(n17870));
   no02f10 U21377 (.o(n20202),
	.a(n23973),
	.b(myLocY_f_2_));
   no03f20 U21378 (.o(n23973),
	.a(n17879),
	.b(n17876),
	.c(n17873));
   na02f10 U21379 (.o(n17873),
	.a(n17875),
	.b(n17874));
   ao22f04 U21380 (.o(n17874),
	.a(n21768),
	.b(proc_input_NIB_storage_data_f_3__36_),
	.c(FE_OCPN25952_n18039),
	.d(proc_input_NIB_storage_data_f_10__36_));
   ao22f06 U21381 (.o(n17878),
	.a(FE_OCPN25933_n24342),
	.b(proc_input_NIB_storage_data_f_0__36_),
	.c(n19705),
	.d(proc_input_NIB_storage_data_f_9__36_));
   na04f10 U21382 (.o(n17879),
	.a(n17883),
	.b(n17882),
	.c(n17881),
	.d(n17880));
   ao22f08 U21383 (.o(n17880),
	.a(n21739),
	.b(proc_input_NIB_storage_data_f_12__36_),
	.c(n17744),
	.d(proc_input_NIB_storage_data_f_4__36_));
   ao22f08 U21384 (.o(n17881),
	.a(FE_OFN191_n24454),
	.b(proc_input_NIB_storage_data_f_13__36_),
	.c(n17780),
	.d(proc_input_NIB_storage_data_f_15__36_));
   ao22f04 U21385 (.o(n17882),
	.a(proc_input_NIB_storage_data_f_14__36_),
	.b(n19769),
	.c(FE_OCPN25822_n21745),
	.d(proc_input_NIB_storage_data_f_2__36_));
   ao22f06 U21386 (.o(n17883),
	.a(FE_OFN169_n24343),
	.b(proc_input_NIB_storage_data_f_8__36_),
	.c(FE_RN_49),
	.d(proc_input_NIB_storage_data_f_5__36_));
   no03f08 U21387 (.o(n20332),
	.a(n26011),
	.b(n26022),
	.c(n25999));
   no02f08 U21388 (.o(n26022),
	.a(FE_RN_67),
	.b(FE_OFN25972_n20135));
   na02f20 U21389 (.o(thanksIn_P),
	.a(n17890),
	.b(n19465));
   ao12f10 U21390 (.o(n25470),
	.a(reset),
	.b(n19466),
	.c(n17890));
   no03f20 U21391 (.o(n17890),
	.a(n26025),
	.b(n26023),
	.c(n26006));
   na02f20 U21392 (.o(n23318),
	.a(n17899),
	.b(n17891));
   no02f10 U21393 (.o(n17891),
	.a(n17896),
	.b(n17892));
   ao22f08 U21394 (.o(n17893),
	.a(proc_input_NIB_storage_data_f_15__55_),
	.b(FE_OCPN25947_n19595),
	.c(proc_input_NIB_storage_data_f_8__55_),
	.d(FE_RN_19));
   ao22f08 U21395 (.o(n17894),
	.a(proc_input_NIB_storage_data_f_1__55_),
	.b(FE_OFN161_n24129),
	.c(n18077),
	.d(proc_input_NIB_storage_data_f_5__55_));
   ao22f08 U21396 (.o(n17895),
	.a(proc_input_NIB_storage_data_f_11__55_),
	.b(FE_OCPN25922_n19547),
	.c(FE_OFN20_n17779),
	.d(proc_input_NIB_storage_data_f_7__55_));
   na02f06 U21397 (.o(n17897),
	.a(proc_input_NIB_storage_data_f_10__55_),
	.b(FE_OCPN25961_n18039));
   na02f08 U21398 (.o(n17903),
	.a(n17905),
	.b(n17904));
   ao22f08 U21399 (.o(n17905),
	.a(proc_input_NIB_storage_data_f_2__55_),
	.b(FE_RN_38),
	.c(proc_input_NIB_storage_data_f_9__55_),
	.d(FE_OFN25682_n17814));
   in01f10 U21400 (.o(n19588),
	.a(n17906));
   no02f10 U21401 (.o(n17906),
	.a(FE_OFN24806_n19655),
	.b(n17907));
   ao12f02 U21403 (.o(n20079),
	.a(n17908),
	.b(proc_input_NIB_storage_data_f_1__23_),
	.c(FE_OFN156_n24129));
   ao12f01 U21406 (.o(n24132),
	.a(n17912),
	.b(proc_input_NIB_storage_data_f_6__2_),
	.c(n19503));
   no02f01 U21407 (.o(n17912),
	.a(FE_OFN24806_n19655),
	.b(n17913));
   in01s01 U21408 (.o(n17913),
	.a(proc_input_NIB_storage_data_f_3__2_));
   na02f20 U21409 (.o(n23512),
	.a(n17914),
	.b(n18225));
   no02f20 U21410 (.o(n17914),
	.a(n19606),
	.b(n19605));
   no02f10 U21411 (.o(n20203),
	.a(myLocY_f_3_),
	.b(n17915));
   na04f10 U21412 (.o(n19545),
	.a(n17919),
	.b(n17918),
	.c(n17917),
	.d(n17916));
   ao22f03 U21413 (.o(n17916),
	.a(proc_input_NIB_storage_data_f_6__37_),
	.b(n19503),
	.c(proc_input_NIB_storage_data_f_3__37_),
	.d(n19709));
   ao22f08 U21414 (.o(n17917),
	.a(n17742),
	.b(proc_input_NIB_storage_data_f_4__37_),
	.c(proc_input_NIB_storage_data_f_13__37_),
	.d(FE_OFN25604_n19530));
   ao22f08 U21415 (.o(n17918),
	.a(proc_input_NIB_storage_data_f_8__37_),
	.b(n24343),
	.c(n20012),
	.d(proc_input_NIB_storage_data_f_9__37_));
   na04f10 U21417 (.o(n19546),
	.a(n17923),
	.b(n17922),
	.c(n17921),
	.d(n17920));
   ao22f08 U21418 (.o(n17920),
	.a(proc_input_NIB_storage_data_f_10__37_),
	.b(n18038),
	.c(n17779),
	.d(proc_input_NIB_storage_data_f_7__37_));
   ao22f08 U21419 (.o(n17921),
	.a(proc_input_NIB_storage_data_f_11__37_),
	.b(n18033),
	.c(proc_input_NIB_storage_data_f_0__37_),
	.d(FE_OCPN25933_n24342));
   ao22f06 U21420 (.o(n17923),
	.a(proc_input_NIB_storage_data_f_2__37_),
	.b(FE_OFN188_n24453),
	.c(FE_RN_49),
	.d(proc_input_NIB_storage_data_f_5__37_));
   no02f20 U21421 (.o(n19591),
	.a(n17926),
	.b(n17924));
   in01f10 U21422 (.o(n17924),
	.a(n17925));
   na02f20 U21423 (.o(n17925),
	.a(proc_input_NIB_storage_data_f_6__51_),
	.b(n19503));
   no02f10 U21424 (.o(n17926),
	.a(n18036),
	.b(n17927));
   ao12m02 U21426 (.o(n24067),
	.a(n17930),
	.b(FE_OCPN25837_n24342),
	.c(proc_input_NIB_storage_data_f_0__4_));
   in01s01 U21427 (.o(n17931),
	.a(proc_input_NIB_storage_data_f_3__4_));
   no02f04 U21429 (.o(n17932),
	.a(FE_OFN24806_n19655),
	.b(n17933));
   na02f80 U21432 (.o(n17934),
	.a(n19495),
	.b(proc_input_NIB_head_ptr_f_0_));
   no02f10 U21433 (.o(n18527),
	.a(n20210),
	.b(n17940));
   no02f10 U21434 (.o(n24954),
	.a(n19736),
	.b(n17940));
   oa22f06 U21435 (.o(n20342),
	.a(n18534),
	.b(n17940),
	.c(n24971),
	.d(n24970));
   in01f08 U21437 (.o(n17941),
	.a(n17942));
   ao22f06 U21438 (.o(n17947),
	.a(proc_input_NIB_storage_data_f_11__54_),
	.b(FE_OCPN25919_n19547),
	.c(proc_input_NIB_storage_data_f_6__54_),
	.d(n19503));
   no02f10 U21439 (.o(n17949),
	.a(n17953),
	.b(n17950));
   na02f10 U21440 (.o(n17950),
	.a(n17952),
	.b(n17951));
   ao22f20 U21441 (.o(n17951),
	.a(proc_input_NIB_storage_data_f_4__54_),
	.b(n21749),
	.c(proc_input_NIB_storage_data_f_12__54_),
	.d(FE_OFN24803_n19500));
   ao22f10 U21442 (.o(n17952),
	.a(proc_input_NIB_storage_data_f_15__54_),
	.b(FE_OCPN25947_n19595),
	.c(proc_input_NIB_storage_data_f_5__54_),
	.d(n18077));
   na02f10 U21443 (.o(n17953),
	.a(n17955),
	.b(n17954));
   ao22f10 U21444 (.o(n17954),
	.a(proc_input_NIB_storage_data_f_14__54_),
	.b(n19769),
	.c(proc_input_NIB_storage_data_f_2__54_),
	.d(FE_OCPN25829_n21745));
   ao22f10 U21445 (.o(n17955),
	.a(proc_input_NIB_storage_data_f_8__54_),
	.b(FE_RN_19),
	.c(proc_input_NIB_storage_data_f_1__54_),
	.d(FE_OFN161_n24129));
   no03f10 U21446 (.o(n19621),
	.a(n17962),
	.b(n17959),
	.c(n17956));
   na02f08 U21447 (.o(n17956),
	.a(n17958),
	.b(n17957));
   na02f08 U21448 (.o(n17959),
	.a(n17961),
	.b(n17960));
   ao22f08 U21449 (.o(n17963),
	.a(proc_input_NIB_storage_data_f_2__59_),
	.b(FE_OCPN25814_FE_OFN186_n24453),
	.c(proc_input_NIB_storage_data_f_14__59_),
	.d(n19769));
   ao22f08 U21450 (.o(n17964),
	.a(proc_input_NIB_storage_data_f_1__59_),
	.b(FE_OFN165_n24129),
	.c(proc_input_NIB_storage_data_f_4__59_),
	.d(FE_RN_59));
   na02f10 U21451 (.o(n17965),
	.a(n17967),
	.b(n17966));
   ao22f10 U21452 (.o(n17967),
	.a(proc_input_NIB_storage_data_f_8__59_),
	.b(FE_OFN168_n24343),
	.c(proc_input_NIB_storage_data_f_15__59_),
	.d(FE_OCPN25947_n19595));
   na02f08 U21453 (.o(n17971),
	.a(n17973),
	.b(n17972));
   ao22f10 U21454 (.o(n17973),
	.a(proc_input_NIB_storage_data_f_12__59_),
	.b(FE_OCPN25968_n19500),
	.c(FE_RN_49),
	.d(proc_input_NIB_storage_data_f_5__59_));
   na02f03 U21455 (.o(n17977),
	.a(proc_input_NIB_storage_data_f_7__47_),
	.b(n17779));
   na03f20 U21456 (.o(n23344),
	.a(n17988),
	.b(n17984),
	.c(n17978));
   no02f10 U21457 (.o(n17978),
	.a(n17981),
	.b(n17979));
   na02f08 U21458 (.o(n17979),
	.a(n18081),
	.b(n17980));
   na02f04 U21459 (.o(n17982),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__50_));
   in01f08 U21460 (.o(n17984),
	.a(n17985));
   na02f06 U21461 (.o(n17985),
	.a(n17987),
	.b(n17986));
   ao22f04 U21462 (.o(n17987),
	.a(FE_OFN25681_n17814),
	.b(proc_input_NIB_storage_data_f_9__50_),
	.c(proc_input_NIB_storage_data_f_11__50_),
	.d(FE_OCPN25923_n19547));
   no02f10 U21463 (.o(n17988),
	.a(n17992),
	.b(n17989));
   na02f08 U21464 (.o(n17989),
	.a(n17991),
	.b(n17990));
   ao22f08 U21465 (.o(n17990),
	.a(n24454),
	.b(proc_input_NIB_storage_data_f_13__50_),
	.c(FE_OCPN25830_n),
	.d(proc_input_NIB_storage_data_f_0__50_));
   ao22f08 U21466 (.o(n17991),
	.a(n18077),
	.b(proc_input_NIB_storage_data_f_5__50_),
	.c(n19769),
	.d(proc_input_NIB_storage_data_f_14__50_));
   na02f08 U21467 (.o(n17992),
	.a(n17994),
	.b(n17993));
   ao22f06 U21468 (.o(n17993),
	.a(FE_OCPN25947_n19595),
	.b(proc_input_NIB_storage_data_f_15__50_),
	.c(FE_OFN170_n24343),
	.d(proc_input_NIB_storage_data_f_8__50_));
   ao22f06 U21469 (.o(n17994),
	.a(FE_OFN161_n24129),
	.b(proc_input_NIB_storage_data_f_1__50_),
	.c(n17742),
	.d(proc_input_NIB_storage_data_f_4__50_));
   na02f10 U21470 (.o(n23504),
	.a(n18002),
	.b(n17995));
   no02f10 U21471 (.o(n18002),
	.a(n18005),
	.b(n18003));
   na02f08 U21472 (.o(n18003),
	.a(n19704),
	.b(n18004));
   na02f08 U21473 (.o(n18005),
	.a(n18007),
	.b(n18006));
   na02f10 U21474 (.o(n22901),
	.a(n18009),
	.b(n18008));
   oa22f04 U21475 (.o(n18010),
	.a(n25028),
	.b(n20139),
	.c(n25017),
	.d(n20502));
   oa12f10 U21476 (.o(n25078),
	.a(n20106),
	.b(n22901),
	.c(n18011));
   na02f04 U21477 (.o(n19784),
	.a(n18014),
	.b(n23482));
   no02f04 U21478 (.o(n24983),
	.a(n18014),
	.b(n24954));
   no02f06 U21479 (.o(n18208),
	.a(n20224),
	.b(n18015));
   no02f20 U21480 (.o(n20475),
	.a(n19743),
	.b(n18015));
   oa22f08 U21481 (.o(n18431),
	.a(n20386),
	.b(n20385),
	.c(n20363),
	.d(n18015));
   no02f06 U21482 (.o(n18016),
	.a(n18228),
	.b(n18230));
   na04f10 U21483 (.o(n18230),
	.a(n18231),
	.b(n18232),
	.c(n18233),
	.d(n18017));
   ao22f10 U21484 (.o(n18017),
	.a(FE_OCPN25968_n19500),
	.b(proc_input_NIB_storage_data_f_12__62_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__62_));
   na03f10 U21485 (.o(n18228),
	.a(n18229),
	.b(n18019),
	.c(n18018));
   na04f10 U21486 (.o(n18226),
	.a(n18227),
	.b(n18023),
	.c(n18022),
	.d(n18021));
   na02f04 U21487 (.o(n18021),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__62_));
   ao22f08 U21488 (.o(n18023),
	.a(FE_RN_59),
	.b(proc_input_NIB_storage_data_f_4__62_),
	.c(FE_OCPN25947_n19595),
	.d(proc_input_NIB_storage_data_f_15__62_));
   na04f20 U21489 (.o(n18433),
	.a(n18027),
	.b(n18026),
	.c(n20381),
	.d(n18025));
   no02f10 U21490 (.o(n18026),
	.a(n18629),
	.b(n19722));
   no02f10 U21491 (.o(n18027),
	.a(n18628),
	.b(n20365));
   ao22f06 U21492 (.o(n19537),
	.a(FE_OFN25636_n19595),
	.b(proc_input_NIB_storage_data_f_15__38_),
	.c(FE_OCPN25910_n19547),
	.d(proc_input_NIB_storage_data_f_11__38_));
   na02f20 U21493 (.o(n18028),
	.a(n18653),
	.b(n18652));
   na02s01 U21494 (.o(n18605),
	.a(FE_OFN575_n25463),
	.b(south_input_NIB_head_ptr_f_0_));
   ao22f06 U21495 (.o(n19599),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__63_),
	.c(FE_OFN170_n24343),
	.d(proc_input_NIB_storage_data_f_8__63_));
   oa22f10 U21497 (.o(n19625),
	.a(myChipID_f_12_),
	.b(n22896),
	.c(n19622),
	.d(n18093));
   in01f10 U21498 (.o(n22869),
	.a(n19188));
   ao22f04 U21499 (.o(n18485),
	.a(proc_input_NIB_storage_data_f_15__35_),
	.b(n17780),
	.c(proc_input_NIB_storage_data_f_4__35_),
	.d(n17744));
   na02f04 U21500 (.o(n18291),
	.a(n18322),
	.b(n18320));
   na02f02 U21501 (.o(n18320),
	.a(proc_input_NIB_storage_data_f_10__41_),
	.b(n18038));
   na02f06 U21502 (.o(n23621),
	.a(n19999),
	.b(n19998));
   na04f08 U21503 (.o(n18029),
	.a(n19571),
	.b(n19574),
	.c(n19572),
	.d(n19573));
   in01f02 U21504 (.o(n18031),
	.a(n18030));
   ao22f08 U21505 (.o(n18419),
	.a(proc_input_NIB_storage_data_f_11__57_),
	.b(FE_OCPN25919_n19547),
	.c(proc_input_NIB_storage_data_f_0__57_),
	.d(FE_OCPN25933_n24342));
   in01f10 U21506 (.o(n23619),
	.a(n19634));
   na02f10 U21508 (.o(n20115),
	.a(n20352),
	.b(n26015));
   na02f08 U21509 (.o(n20919),
	.a(n18712),
	.b(n18711));
   in01f10 U21510 (.o(n21365),
	.a(n18754));
   in01f06 U21511 (.o(n19235),
	.a(n23302));
   no02f06 U21512 (.o(n20392),
	.a(n23302),
	.b(n19719));
   oa12f10 U21513 (.o(n18069),
	.a(n19584),
	.b(n21509),
	.c(n21508));
   no02f20 U21514 (.o(n26016),
	.a(n20504),
	.b(n20107));
   na02f02 U21515 (.o(n2418),
	.a(n18572),
	.b(n18576));
   ao22f04 U21516 (.o(n18321),
	.a(proc_input_NIB_storage_data_f_11__41_),
	.b(FE_OFN25674_n18033),
	.c(proc_input_NIB_storage_data_f_15__41_),
	.d(FE_OFN25637_n19595));
   no02f08 U21517 (.o(n25175),
	.a(n20534),
	.b(n22771));
   ao22f20 U21518 (.o(n19332),
	.a(n24359),
	.b(east_input_NIB_storage_data_f_2__59_),
	.c(FE_OCPN25813_FE_OFN24735_n19306),
	.d(east_input_NIB_storage_data_f_1__59_));
   na04f40 U21519 (.o(n19410),
	.a(n19361),
	.b(n19360),
	.c(n19359),
	.d(n19358));
   no02f20 U21520 (.o(n19358),
	.a(n19357),
	.b(n19356));
   na04f04 U21521 (.o(n2838),
	.a(n25480),
	.b(n25479),
	.c(n25478),
	.d(n25477));
   na03f10 U21522 (.o(n18480),
	.a(n18483),
	.b(n18482),
	.c(n18481));
   ao22f02 U21523 (.o(n18517),
	.a(proc_input_NIB_storage_data_f_13__45_),
	.b(FE_OFN191_n24454),
	.c(proc_input_NIB_storage_data_f_0__45_),
	.d(FE_OCPN25835_n24342));
   na02f08 U21524 (.o(n18465),
	.a(n20115),
	.b(n20114));
   na02f20 U21525 (.o(n20114),
	.a(n26014),
	.b(n25079));
   in01f40 U21534 (.o(n18754),
	.a(FE_RN_41));
   no02f10 U21535 (.o(n18925),
	.a(FE_RN_7),
	.b(n18922));
   na02f08 U21536 (.o(n18422),
	.a(n22834),
	.b(myLocY_f_0_));
   na04f08 U21537 (.o(n19560),
	.a(n19554),
	.b(n19553),
	.c(n19552),
	.d(n19551));
   na02f06 U21538 (.o(n25151),
	.a(n17779),
	.b(n25995));
   na02f06 U21539 (.o(n21907),
	.a(east_input_valid),
	.b(n20622));
   no02f02 U21540 (.o(n18058),
	.a(n25086),
	.b(n25085));
   no02f06 U21541 (.o(n25101),
	.a(n25086),
	.b(n25085));
   na04f10 U21542 (.o(n19539),
	.a(n19538),
	.b(n19537),
	.c(n19536),
	.d(n19535));
   oa22f08 U21543 (.o(n19739),
	.a(myLocY_f_4_),
	.b(FE_RN_21),
	.c(myLocY_f_5_),
	.d(n22857));
   no02f10 U21544 (.o(n22888),
	.a(n19540),
	.b(n19539));
   ao22f10 U21545 (.o(n19563),
	.a(myLocY_f_4_),
	.b(n22888),
	.c(myLocY_f_3_),
	.d(n18104));
   no02f04 U21546 (.o(n20369),
	.a(n19722),
	.b(n19721));
   na04f20 U21547 (.o(n21416),
	.a(n19570),
	.b(n18067),
	.c(n19569),
	.d(n18066));
   ao22f08 U21548 (.o(n19569),
	.a(n20056),
	.b(proc_input_NIB_storage_data_f_9__58_),
	.c(FE_RN_59),
	.d(proc_input_NIB_storage_data_f_4__58_));
   oa12f02 U21549 (.o(n19469),
	.a(n18082),
	.b(n18405),
	.c(n25470));
   na03f06 U21550 (.o(n25479),
	.a(n25470),
	.b(proc_input_NIB_elements_in_array_f_3_),
	.c(n25469));
   ao22f04 U21551 (.o(n19538),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__38_),
	.c(FE_OFN156_n24129),
	.d(proc_input_NIB_storage_data_f_1__38_));
   oa12f02 U21552 (.o(n20119),
	.a(n20117),
	.b(n20504),
	.c(n20118));
   na02f03 U21553 (.o(n25423),
	.a(FE_OFN25599_reset),
	.b(n18493));
   in01f08 U21554 (.o(n18146),
	.a(n23344));
   no02f10 U21555 (.o(n19564),
	.a(n20203),
	.b(n20202));
   na02f08 U21556 (.o(n18484),
	.a(n18486),
	.b(n18485));
   ao22f20 U21557 (.o(n19592),
	.a(FE_OFN161_n24129),
	.b(proc_input_NIB_storage_data_f_1__51_),
	.c(FE_OFN170_n24343),
	.d(proc_input_NIB_storage_data_f_8__51_));
   na02f08 U21558 (.o(n18216),
	.a(n20352),
	.b(n26024));
   na03f04 U21559 (.o(n25116),
	.a(n20465),
	.b(n23036),
	.c(n20464));
   ao22f06 U21560 (.o(n25155),
	.a(n20467),
	.b(n19833),
	.c(n20464),
	.d(n20379));
   oa22f08 U21561 (.o(n19670),
	.a(myChipID_f_2_),
	.b(n23637),
	.c(n23344),
	.d(n19657));
   no02f08 U21562 (.o(n26021),
	.a(FE_RN_67),
	.b(n20139));
   no02f06 U21563 (.o(validOut_N),
	.a(FE_RN_67),
	.b(n20136));
   no04f40 U21564 (.o(n20417),
	.a(n18701),
	.b(n18699),
	.c(n18700),
	.d(n18698));
   na04f40 U21565 (.o(n18699),
	.a(n18691),
	.b(n18690),
	.c(n18689),
	.d(n18688));
   in01f04 U21566 (.o(n25086),
	.a(n25084));
   oa12f02 U21567 (.o(n24986),
	.a(n24979),
	.b(n25406),
	.c(n24980));
   in01f02 U21568 (.o(n24984),
	.a(n24983));
   na04f10 U21569 (.o(n21509),
	.a(n19579),
	.b(n19578),
	.c(n19577),
	.d(n19576));
   no03f04 U21570 (.o(n18495),
	.a(n25033),
	.b(n25309),
	.c(n25035));
   ao12f08 U21571 (.o(n25387),
	.a(n20257),
	.b(n20258),
	.c(n25000));
   ao22f08 U21572 (.o(n18154),
	.a(proc_input_NIB_storage_data_f_1__56_),
	.b(FE_OFN161_n24129),
	.c(proc_input_NIB_storage_data_f_7__56_),
	.d(FE_OFN20_n17779));
   ao22f06 U21573 (.o(n19521),
	.a(FE_OCPN25913_n19547),
	.b(proc_input_NIB_storage_data_f_11__39_),
	.c(FE_OFN169_n24343),
	.d(proc_input_NIB_storage_data_f_8__39_));
   ao22f10 U21574 (.o(n18886),
	.a(FE_RN_5),
	.b(west_input_NIB_storage_data_f_3__53_),
	.c(n18960),
	.d(west_input_NIB_storage_data_f_2__53_));
   in01f10 U21575 (.o(n19646),
	.a(n23637));
   no02f10 U21577 (.o(n23637),
	.a(n19645),
	.b(n19644));
   ao12m02 U21578 (.o(n20035),
	.a(n18425),
	.b(proc_input_NIB_storage_data_f_6__25_),
	.c(n19503));
   na04f10 U21579 (.o(n19645),
	.a(n19639),
	.b(n19638),
	.c(n19637),
	.d(n19636));
   na02f08 U21580 (.o(n18402),
	.a(n25000),
	.b(n23034));
   no02f04 U21581 (.o(n20133),
	.a(n18640),
	.b(n20132));
   no02f06 U21582 (.o(n18640),
	.a(n18641),
	.b(n18507));
   ao22f20 U21583 (.o(n19359),
	.a(n19594),
	.b(n25512),
	.c(n19347),
	.d(n19346));
   no02f04 U21584 (.o(n20112),
	.a(n19889),
	.b(n19888));
   no02f08 U21585 (.o(n25329),
	.a(n25998),
	.b(n26008));
   no02f10 U21586 (.o(n26008),
	.a(FE_OFN902_n18421),
	.b(n17759));
   no02f08 U21587 (.o(n25985),
	.a(FE_RN_67),
	.b(n20502));
   no02f20 U21588 (.o(n26023),
	.a(n18185),
	.b(n20137));
   oa12f10 U21589 (.o(n18065),
	.a(n19575),
	.b(n21416),
	.c(n21415));
   no02f08 U21590 (.o(n18358),
	.a(n18364),
	.b(n18359));
   na02f10 U21591 (.o(n19606),
	.a(n19602),
	.b(n19601));
   na04f10 U21592 (.o(n21415),
	.a(n19571),
	.b(n19574),
	.c(n19572),
	.d(n19573));
   no02f10 U21593 (.o(n22857),
	.a(n19529),
	.b(n18130));
   na04f10 U21594 (.o(n19644),
	.a(n19643),
	.b(n19642),
	.c(n19641),
	.d(n19640));
   no04f40 U21595 (.o(n19361),
	.a(n19336),
	.b(n19335),
	.c(n19334),
	.d(n19333));
   na02f20 U21596 (.o(n23611),
	.a(n19343),
	.b(n19342));
   ao22f20 U21597 (.o(n19343),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__56_),
	.c(FE_OCPN25813_FE_OFN24735_n19306),
	.d(east_input_NIB_storage_data_f_1__56_));
   na04f10 U21598 (.o(n19529),
	.a(n19528),
	.b(n19527),
	.c(n19526),
	.d(n19525));
   no02f06 U21600 (.o(n18351),
	.a(n18715),
	.b(n18352));
   ao22f08 U21601 (.o(n18745),
	.a(n24472),
	.b(south_input_NIB_storage_data_f_0__44_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__44_));
   na03f08 U21602 (.o(n18622),
	.a(n20417),
	.b(n19027),
	.c(n19833));
   no02f06 U21605 (.o(n21582),
	.a(n19937),
	.b(n19936));
   no02f06 U21606 (.o(n21569),
	.a(n19928),
	.b(n19927));
   na04f10 U21607 (.o(n18130),
	.a(n19523),
	.b(n19524),
	.c(n19521),
	.d(n19522));
   no02f10 U21608 (.o(n20273),
	.a(n19701),
	.b(n23325));
   na04f10 U21609 (.o(n18511),
	.a(n19718),
	.b(n18514),
	.c(n18513),
	.d(n18512));
   no02f04 U21610 (.o(n20425),
	.a(n25155),
	.b(n25154));
   no02f02 U21611 (.o(n25312),
	.a(n25034),
	.b(n25033));
   ao12f04 U21612 (.o(n18297),
	.a(myLocY_f_2_),
	.b(n18705),
	.c(n18704));
   in01f02 U21613 (.o(n20131),
	.a(n18631));
   no02f10 U21614 (.o(n20391),
	.a(n19235),
	.b(myLocX_f_3_));
   na02f04 U21615 (.o(n18084),
	.a(n22926),
	.b(myLocY_f_7_));
   no02f10 U21616 (.o(n18880),
	.a(n19701),
	.b(n23323));
   na02f10 U21617 (.o(n25083),
	.a(n18217),
	.b(n18216));
   no03f10 U21618 (.o(n18378),
	.a(n20372),
	.b(n18380),
	.c(n18379));
   no03f08 U21619 (.o(n20505),
	.a(n25984),
	.b(n25997),
	.c(n25985));
   ao12s01 U21620 (.o(n25368),
	.a(n25370),
	.b(n25374),
	.c(n25367));
   oa22f20 U21621 (.o(n19649),
	.a(myChipID_f_5_),
	.b(n19648),
	.c(n19647),
	.d(n19646));
   na02f10 U21622 (.o(n18415),
	.a(proc_input_NIB_storage_data_f_7__57_),
	.b(FE_OFN20_n17779));
   no04f04 U21623 (.o(n18869),
	.a(n18875),
	.b(n18876),
	.c(n19720),
	.d(n18874));
   no02f06 U21624 (.o(n24997),
	.a(n22902),
	.b(n23482));
   no03f10 U21625 (.o(n19248),
	.a(n20409),
	.b(n19247),
	.c(n19871));
   na02f03 U21626 (.o(n19841),
	.a(n19325),
	.b(n20919));
   na03f06 U21627 (.o(n19796),
	.a(n19795),
	.b(n19794),
	.c(n19817));
   ao22f01 U21628 (.o(n24227),
	.a(proc_input_NIB_storage_data_f_11__15_),
	.b(FE_OCPN25909_n19547),
	.c(proc_input_NIB_storage_data_f_15__15_),
	.d(FE_OFN25635_n19595));
   ao22f02 U21629 (.o(n19773),
	.a(FE_OFN25604_n19530),
	.b(proc_input_NIB_storage_data_f_13__30_),
	.c(n17742),
	.d(proc_input_NIB_storage_data_f_4__30_));
   na02f02 U21630 (.o(n19775),
	.a(n19771),
	.b(n19770));
   ao22f02 U21631 (.o(n19770),
	.a(n17747),
	.b(proc_input_NIB_storage_data_f_12__30_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__30_));
   na02f02 U21632 (.o(n19781),
	.a(n19777),
	.b(n19776));
   ao22f02 U21633 (.o(n19776),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__30_),
	.c(FE_OFN25637_n19595),
	.d(proc_input_NIB_storage_data_f_15__30_));
   ao22f04 U21634 (.o(n19758),
	.a(FE_OFN25678_n17814),
	.b(proc_input_NIB_storage_data_f_9__31_),
	.c(FE_OCPN25933_n24342),
	.d(proc_input_NIB_storage_data_f_0__31_));
   na02f02 U21635 (.o(n19755),
	.a(n19751),
	.b(n19750));
   ao22f02 U21636 (.o(n19751),
	.a(FE_OFN25604_n19530),
	.b(proc_input_NIB_storage_data_f_13__32_),
	.c(n17744),
	.d(proc_input_NIB_storage_data_f_4__32_));
   na02f02 U21637 (.o(n19749),
	.a(n19745),
	.b(n19744));
   ao22f06 U21638 (.o(n19523),
	.a(proc_input_NIB_storage_data_f_0__39_),
	.b(n18131),
	.c(proc_input_NIB_storage_data_f_5__39_),
	.d(FE_RN_49));
   ao22f04 U21639 (.o(n19522),
	.a(n21768),
	.b(proc_input_NIB_storage_data_f_3__39_),
	.c(n19769),
	.d(proc_input_NIB_storage_data_f_14__39_));
   na02f04 U21640 (.o(n18360),
	.a(proc_input_NIB_storage_data_f_1__43_),
	.b(FE_OFN161_n24129));
   na02f06 U21641 (.o(n18513),
	.a(proc_input_NIB_storage_data_f_8__45_),
	.b(FE_OFN167_n24343));
   no02f04 U21642 (.o(n18206),
	.a(n20265),
	.b(n20236));
   na02f02 U21643 (.o(n20236),
	.a(n20235),
	.b(n20264));
   no02f10 U21644 (.o(n19825),
	.a(n20244),
	.b(n20247));
   no03f02 U21645 (.o(n20406),
	.a(n20405),
	.b(n20404),
	.c(n20403));
   no02f04 U21646 (.o(n20384),
	.a(n18556),
	.b(n18554));
   no02f01 U21647 (.o(n21156),
	.a(east_input_control_count_f_0_),
	.b(east_input_control_count_f_1_));
   no04f02 U21648 (.o(n21902),
	.a(east_input_control_count_f_4_),
	.b(east_input_control_count_f_5_),
	.c(east_input_control_count_f_3_),
	.d(east_input_control_count_f_2_));
   no02f08 U21649 (.o(n19147),
	.a(n20166),
	.b(n19117));
   oa22f08 U21650 (.o(n19145),
	.a(n20160),
	.b(n19144),
	.c(n20737),
	.d(n20170));
   no02s01 U21651 (.o(n20703),
	.a(north_input_control_count_f_0_),
	.b(north_input_control_count_f_1_));
   oa22f02 U21652 (.o(n20288),
	.a(n20420),
	.b(n20414),
	.c(n20419),
	.d(n20287));
   ao22f02 U21653 (.o(n20057),
	.a(n19705),
	.b(proc_input_NIB_storage_data_f_9__27_),
	.c(FE_OCPN25953_n18039),
	.d(proc_input_NIB_storage_data_f_10__27_));
   ao22f02 U21654 (.o(n20100),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__24_),
	.c(FE_OFN25637_n19595),
	.d(proc_input_NIB_storage_data_f_15__24_));
   ao22f02 U21655 (.o(n20098),
	.a(n24060),
	.b(proc_input_NIB_storage_data_f_9__24_),
	.c(n18051),
	.d(proc_input_NIB_storage_data_f_10__24_));
   no02s01 U21656 (.o(n25355),
	.a(n25370),
	.b(n25354));
   no02f20 U21657 (.o(n20464),
	.a(n20417),
	.b(n20377));
   ao22f01 U21658 (.o(n24659),
	.a(n25295),
	.b(FE_OFN528_n24732),
	.c(FE_OFN79_n20501),
	.d(FE_OFN237_n24730));
   ao22f01 U21659 (.o(n24651),
	.a(n25295),
	.b(n24685),
	.c(FE_OFN79_n20501),
	.d(FE_OFN229_n24684));
   ao22f01 U21660 (.o(n24654),
	.a(n25295),
	.b(n24705),
	.c(FE_OFN79_n20501),
	.d(FE_OFN231_n24704));
   ao22f01 U21661 (.o(n24580),
	.a(n25295),
	.b(FE_OFN495_n24579),
	.c(FE_OFN79_n20501),
	.d(n24578));
   ao22f01 U21662 (.o(n24589),
	.a(n25295),
	.b(n24588),
	.c(FE_OFN79_n20501),
	.d(n24587));
   ao22f01 U21663 (.o(n24679),
	.a(n25295),
	.b(n24678),
	.c(FE_OFN79_n20501),
	.d(FE_OFN227_n24677));
   ao22f01 U21664 (.o(n24594),
	.a(n25294),
	.b(n24742),
	.c(FE_OFN79_n20501),
	.d(FE_OFN242_n24744));
   ao22f01 U21665 (.o(n24725),
	.a(n25295),
	.b(n24721),
	.c(FE_OFN79_n20501),
	.d(n24720));
   ao22f01 U21666 (.o(n24715),
	.a(n25295),
	.b(n24714),
	.c(FE_OFN79_n20501),
	.d(n24713));
   na02f04 U21667 (.o(n22771),
	.a(west_output_current_route_connection_2_),
	.b(n25153));
   ao22f01 U21668 (.o(n24369),
	.a(n19019),
	.b(FE_OFN528_n24732),
	.c(n19017),
	.d(FE_OFN237_n24730));
   ao22f01 U21669 (.o(n24339),
	.a(n19017),
	.b(FE_OFN221_n24662),
	.c(n19020),
	.d(n24663));
   ao22f01 U21670 (.o(n24440),
	.a(n19019),
	.b(n24705),
	.c(n19017),
	.d(FE_OFN231_n24704));
   ao22f01 U21671 (.o(n24432),
	.a(n19019),
	.b(FE_OFN495_n24579),
	.c(n19017),
	.d(n24578));
   ao22f01 U21672 (.o(n21399),
	.a(n19017),
	.b(FE_OFN136_n23623),
	.c(n19022),
	.d(n23622));
   in01m06 U21673 (.o(n20531),
	.a(west_output_current_route_connection_2_));
   in01f02 U21674 (.o(n18286),
	.a(n18287));
   ao12s01 U21675 (.o(n20705),
	.a(n20704),
	.b(north_input_control_count_f_6_),
	.c(n20707));
   no02s01 U21676 (.o(n20704),
	.a(n20707),
	.b(north_input_control_count_f_6_));
   ao22s01 U21677 (.o(n21897),
	.a(n20723),
	.b(north_input_control_count_f_1_),
	.c(n20722),
	.d(n20721));
   no02f20 U21678 (.o(n18185),
	.a(n19053),
	.b(n19052));
   na02f20 U21679 (.o(n19052),
	.a(n19051),
	.b(n19050));
   no02f10 U21680 (.o(n20388),
	.a(myLocX_f_1_),
	.b(n19231));
   no02f10 U21681 (.o(n20365),
	.a(n19706),
	.b(FE_RN_39));
   oa12f01 U21682 (.o(n20187),
	.a(n20184),
	.b(n20186),
	.c(n20185));
   no02f10 U21683 (.o(n20186),
	.a(myLocY_f_3_),
	.b(n22875));
   oa12f02 U21684 (.o(n19827),
	.a(n20144),
	.b(n19820),
	.c(n20143));
   na02f04 U21685 (.o(n20169),
	.a(n19132),
	.b(n21141));
   na03f06 U21686 (.o(n18171),
	.a(n19085),
	.b(n19084),
	.c(myLocY_f_5_));
   na02f06 U21687 (.o(n20153),
	.a(n19121),
	.b(n19124));
   no02f06 U21688 (.o(n19040),
	.a(n19037),
	.b(n19036));
   na02f06 U21689 (.o(n18779),
	.a(n24165),
	.b(south_input_NIB_storage_data_f_2__32_));
   ao22f06 U21690 (.o(n18482),
	.a(proc_input_NIB_storage_data_f_14__35_),
	.b(FE_OFN25644_n19504),
	.c(proc_input_NIB_storage_data_f_5__35_),
	.d(FE_RN_49));
   na03f10 U21691 (.o(n18156),
	.a(n18154),
	.b(n18153),
	.c(n18152));
   ao22f08 U21692 (.o(n18153),
	.a(proc_input_NIB_storage_data_f_14__56_),
	.b(n19769),
	.c(proc_input_NIB_storage_data_f_5__56_),
	.d(n18077));
   ao22f40 U21693 (.o(n20747),
	.a(FE_OFN24763_n18960),
	.b(west_input_NIB_storage_data_f_2__60_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__60_));
   no02f08 U21694 (.o(n18468),
	.a(myLocY_f_0_),
	.b(n22834));
   no03f08 U21695 (.o(n18884),
	.a(n18880),
	.b(n20434),
	.c(n18965));
   no02f20 U21696 (.o(n19043),
	.a(n19838),
	.b(n19848));
   no02f04 U21697 (.o(n20356),
	.a(west_output_current_route_connection_2_),
	.b(west_output_current_route_connection_0_));
   ao22f08 U21698 (.o(n19005),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__34_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__34_));
   ao22f08 U21699 (.o(n19006),
	.a(FE_OFN28_n18974),
	.b(west_input_NIB_storage_data_f_0__34_),
	.c(FE_OFN24764_n18960),
	.d(west_input_NIB_storage_data_f_2__34_));
   ao22f06 U21700 (.o(n19536),
	.a(n21768),
	.b(proc_input_NIB_storage_data_f_3__38_),
	.c(n17744),
	.d(proc_input_NIB_storage_data_f_4__38_));
   ao22f08 U21701 (.o(n18984),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__39_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__39_));
   ao22f06 U21702 (.o(n19514),
	.a(FE_RN_38),
	.b(proc_input_NIB_storage_data_f_2__40_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__40_));
   ao22f02 U21703 (.o(n19692),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__46_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__46_));
   ao22f02 U21704 (.o(n19697),
	.a(n20012),
	.b(proc_input_NIB_storage_data_f_9__46_),
	.c(FE_OCPN25949_n18039),
	.d(proc_input_NIB_storage_data_f_10__46_));
   ao22f02 U21705 (.o(n19683),
	.a(n17779),
	.b(proc_input_NIB_storage_data_f_7__48_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__48_));
   ao22f02 U21706 (.o(n19682),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__48_),
	.c(FE_OFN25637_n19595),
	.d(proc_input_NIB_storage_data_f_15__48_));
   ao22f02 U21707 (.o(n19680),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__48_),
	.c(FE_OFN25604_n19530),
	.d(proc_input_NIB_storage_data_f_13__48_));
   ao22f02 U21708 (.o(n19681),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__48_),
	.c(n17747),
	.d(proc_input_NIB_storage_data_f_12__48_));
   ao22f04 U21709 (.o(n19672),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__49_),
	.c(FE_OFN25604_n19530),
	.d(proc_input_NIB_storage_data_f_13__49_));
   ao22f02 U21710 (.o(n19673),
	.a(n17747),
	.b(proc_input_NIB_storage_data_f_12__49_),
	.c(proc_input_NIB_storage_data_f_5__49_),
	.d(FE_RN_49));
   na02f08 U21712 (.o(n18236),
	.a(n18416),
	.b(n18418));
   ao22f06 U21713 (.o(n19574),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__58_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__58_));
   in01f06 U21714 (.o(n18100),
	.a(n21416));
   ao22f08 U21715 (.o(n19609),
	.a(FE_OCPN25968_n19500),
	.b(proc_input_NIB_storage_data_f_12__60_),
	.c(FE_OCPN25933_n24342),
	.d(proc_input_NIB_storage_data_f_0__60_));
   ao22f08 U21716 (.o(n19608),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__60_),
	.c(n17741),
	.d(proc_input_NIB_storage_data_f_4__60_));
   ao22f06 U21717 (.o(n19613),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__60_),
	.c(FE_OCPN25814_FE_OFN186_n24453),
	.d(proc_input_NIB_storage_data_f_2__60_));
   ao22f08 U21718 (.o(n19611),
	.a(FE_OFN165_n24129),
	.b(proc_input_NIB_storage_data_f_1__60_),
	.c(FE_OFN170_n24343),
	.d(proc_input_NIB_storage_data_f_8__60_));
   in01f10 U21719 (.o(n18149),
	.a(n19338));
   no02s01 U21720 (.o(n25457),
	.a(west_output_space_count_f_1_),
	.b(west_output_space_count_f_0_));
   no02f06 U21721 (.o(n25094),
	.a(n19054),
	.b(n25124));
   no02f06 U21722 (.o(n19252),
	.a(south_output_current_route_connection_2_),
	.b(n24989));
   no02f03 U21723 (.o(n25300),
	.a(n25007),
	.b(n25006));
   no02f02 U21724 (.o(n18198),
	.a(n26008),
	.b(n18600));
   no02f02 U21725 (.o(n20518),
	.a(n23400),
	.b(n20517));
   no03s02 U21726 (.o(n20707),
	.a(north_input_control_count_f_5_),
	.b(north_input_control_count_f_4_),
	.c(n20734));
   in01s20 U21727 (.o(n20318),
	.a(east_output_current_route_connection_2_));
   no02f03 U21728 (.o(n20547),
	.a(n25028),
	.b(n20324));
   no02f02 U21729 (.o(n18201),
	.a(n20237),
	.b(n24970));
   ao22f02 U21730 (.o(n19023),
	.a(n19020),
	.b(north_input_valid),
	.c(n19022),
	.d(south_input_valid));
   ao22f02 U21731 (.o(n20042),
	.a(FE_OFN169_n24343),
	.b(proc_input_NIB_storage_data_f_8__25_),
	.c(n17744),
	.d(proc_input_NIB_storage_data_f_4__25_));
   ao22m02 U21732 (.o(n20041),
	.a(n19705),
	.b(proc_input_NIB_storage_data_f_9__25_),
	.c(n18034),
	.d(proc_input_NIB_storage_data_f_10__25_));
   no02s01 U21733 (.o(n25352),
	.a(n25374),
	.b(north_output_space_count_f_1_));
   no02s01 U21734 (.o(n25372),
	.a(north_output_space_count_f_0_),
	.b(north_output_space_count_f_1_));
   ao12m02 U21735 (.o(n19975),
	.a(n18339),
	.b(FE_OCPN25941_n24965),
	.c(south_input_NIB_storage_data_f_3__22_));
   no04f01 U21736 (.o(n25241),
	.a(south_input_control_count_f_5_),
	.b(south_input_control_count_f_3_),
	.c(south_input_control_count_f_2_),
	.d(south_input_control_count_f_7_));
   no04f08 U21737 (.o(n19792),
	.a(n20240),
	.b(n19803),
	.c(n19822),
	.d(n19821));
   in01f02 U21738 (.o(n23100),
	.a(n23044));
   na02f02 U21739 (.o(n23044),
	.a(proc_input_NIB_tail_ptr_f_2_),
	.b(n23734));
   no02s01 U21740 (.o(n25791),
	.a(n25789),
	.b(n25788));
   na02f02 U21741 (.o(n24693),
	.a(n24141),
	.b(n24140));
   ao22f01 U21742 (.o(n23979),
	.a(n25295),
	.b(n23975),
	.c(FE_OFN79_n20501),
	.d(n23974));
   ao22f01 U21743 (.o(n23581),
	.a(n25295),
	.b(n23580),
	.c(FE_OFN79_n20501),
	.d(n23579));
   na02f02 U21744 (.o(n24619),
	.a(n24233),
	.b(n24232));
   na02f02 U21745 (.o(n24630),
	.a(n24471),
	.b(n24470));
   na02f02 U21746 (.o(n24637),
	.a(n24164),
	.b(n24163));
   ao22m02 U21747 (.o(n19965),
	.a(FE_RN_17),
	.b(south_input_NIB_storage_data_f_2__23_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__23_));
   ao22f02 U21748 (.o(n19966),
	.a(FE_OCPN25941_n24965),
	.b(south_input_NIB_storage_data_f_3__23_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__23_));
   ao22f01 U21749 (.o(n24024),
	.a(n25295),
	.b(n24020),
	.c(FE_OFN79_n20501),
	.d(FE_OFN151_n24019));
   ao22f01 U21750 (.o(n23634),
	.a(n25295),
	.b(n23630),
	.c(FE_OFN79_n20501),
	.d(n23629));
   in01s01 U21751 (.o(n18268),
	.a(n18269));
   ao22f01 U21752 (.o(n24735),
	.a(FE_OFN94_n21695),
	.b(n24734),
	.c(n17755),
	.d(FE_OFN530_n24733));
   ao22m02 U21753 (.o(n24548),
	.a(FE_OFN94_n21695),
	.b(FE_OFN223_n24664),
	.c(FE_OFN389_n17786),
	.d(n24665));
   ao22f01 U21754 (.o(n24698),
	.a(FE_OFN94_n21695),
	.b(n24694),
	.c(FE_OFN111_n22773),
	.d(n24693));
   ao22f01 U21755 (.o(n24688),
	.a(FE_OFN94_n21695),
	.b(n24687),
	.c(n17755),
	.d(n24686));
   ao22f01 U21756 (.o(n24707),
	.a(FE_OFN94_n21695),
	.b(n24703),
	.c(n17755),
	.d(FE_OFN515_n24702));
   ao22f01 U21757 (.o(n22355),
	.a(FE_OFN94_n21695),
	.b(n24012),
	.c(n17755),
	.d(FE_OFN487_n24013));
   ao22f01 U21758 (.o(n22343),
	.a(FE_OFN94_n21695),
	.b(n23561),
	.c(FE_OFN389_n17786),
	.d(n23562));
   ao22f01 U21759 (.o(n22359),
	.a(FE_OFN94_n21695),
	.b(n23149),
	.c(FE_OFN111_n22773),
	.d(FE_OFN116_n23148));
   ao22f01 U21760 (.o(n22347),
	.a(FE_OFN94_n21695),
	.b(n23570),
	.c(FE_OFN389_n17786),
	.d(n23571));
   ao22f01 U21761 (.o(n22368),
	.a(FE_OFN94_n21695),
	.b(n23577),
	.c(n17755),
	.d(FE_OFN477_n23578));
   ao22f01 U21762 (.o(n24557),
	.a(FE_OFN94_n21695),
	.b(n24576),
	.c(n17755),
	.d(FE_OFN493_n24577));
   na02f02 U21763 (.o(n24587),
	.a(n24304),
	.b(n24303));
   ao22f01 U21764 (.o(n24573),
	.a(FE_OFN94_n21695),
	.b(n24585),
	.c(n17755),
	.d(FE_OFN497_n24586));
   ao22f01 U21765 (.o(n24537),
	.a(FE_OFN94_n21695),
	.b(n24598),
	.c(FE_OFN389_n17786),
	.d(n24599));
   ao22f01 U21766 (.o(n24565),
	.a(FE_OFN94_n21695),
	.b(n24675),
	.c(n17755),
	.d(n24676));
   ao22f01 U21767 (.o(n24624),
	.a(FE_OFN94_n21695),
	.b(n24620),
	.c(FE_OFN111_n22773),
	.d(FE_OFN207_n24619));
   ao22f01 U21768 (.o(n24632),
	.a(FE_OFN94_n21695),
	.b(n24631),
	.c(FE_OFN111_n22773),
	.d(FE_OFN211_n24630));
   ao22f01 U21769 (.o(n24642),
	.a(FE_OFN94_n21695),
	.b(n24638),
	.c(FE_OFN111_n22773),
	.d(FE_OFN217_n24637));
   na02f02 U21770 (.o(n24752),
	.a(n24396),
	.b(n24395));
   ao22f01 U21771 (.o(n24545),
	.a(FE_OFN94_n21695),
	.b(n24750),
	.c(FE_OFN389_n17786),
	.d(FE_OFN546_n24751));
   ao22f01 U21772 (.o(n24541),
	.a(FE_OFN94_n21695),
	.b(n24740),
	.c(FE_OFN389_n17786),
	.d(n24741));
   ao22f01 U21773 (.o(n24560),
	.a(FE_OFN94_n21695),
	.b(n24722),
	.c(n17755),
	.d(FE_OFN521_n24723));
   na02f04 U21774 (.o(n24713),
	.a(n24329),
	.b(n24328));
   ao22f01 U21775 (.o(n24569),
	.a(FE_OFN94_n21695),
	.b(n24711),
	.c(n17755),
	.d(FE_OFN517_n24712));
   ao22f01 U21776 (.o(n22351),
	.a(FE_OFN94_n21695),
	.b(n24021),
	.c(n17755),
	.d(FE_OFN491_n24022));
   ao22f01 U21777 (.o(n22218),
	.a(FE_OFN94_n21695),
	.b(n23632),
	.c(FE_OFN389_n17786),
	.d(n23630));
   na02f08 U21778 (.o(n22518),
	.a(south_output_current_route_connection_0_),
	.b(n19861));
   ao22f01 U21779 (.o(n24335),
	.a(n19017),
	.b(n24693),
	.c(FE_OFN42_n19022),
	.d(n24694));
   ao22f01 U21780 (.o(n21373),
	.a(n19019),
	.b(FE_OFN485_n24011),
	.c(n19017),
	.d(FE_OFN146_n24010));
   ao22f01 U21781 (.o(n21764),
	.a(n19017),
	.b(FE_OFN116_n23148),
	.c(FE_OFN42_n19022),
	.d(n23149));
   ao22f01 U21782 (.o(n24428),
	.a(n19019),
	.b(n24588),
	.c(n19017),
	.d(n24587));
   na02f02 U21783 (.o(n24600),
	.a(n24284),
	.b(n24283));
   in01f10 U21784 (.o(n18620),
	.a(n18621));
   na02f02 U21785 (.o(n24730),
	.a(n24361),
	.b(n24360));
   na02f02 U21786 (.o(n24662),
	.a(n24098),
	.b(n24097));
   ao22f01 U21787 (.o(n24103),
	.a(FE_OFN366_n17753),
	.b(FE_OFN223_n24664),
	.c(n19057),
	.d(n24665));
   na02f02 U21788 (.o(n24684),
	.a(n24051),
	.b(n24050));
   na02f02 U21789 (.o(n24704),
	.a(n24077),
	.b(n24076));
   na02f03 U21790 (.o(n24578),
	.a(n24122),
	.b(n24121));
   na02f02 U21791 (.o(n24677),
	.a(n24260),
	.b(n24259));
   na02f02 U21792 (.o(n24744),
	.a(n24216),
	.b(n24215));
   ao22f01 U21793 (.o(n24218),
	.a(FE_OFN366_n17753),
	.b(n24740),
	.c(n19057),
	.d(n24741));
   na02f02 U21794 (.o(n24720),
	.a(n24187),
	.b(n24186));
   ao22m02 U21795 (.o(n19958),
	.a(FE_OCPN25943_n24965),
	.b(south_input_NIB_storage_data_f_3__26_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__26_));
   ao22m02 U21796 (.o(n19957),
	.a(n24165),
	.b(south_input_NIB_storage_data_f_2__26_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__26_));
   ao22m02 U21797 (.o(n19959),
	.a(FE_RN_17),
	.b(south_input_NIB_storage_data_f_2__27_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__27_));
   na02f02 U21798 (.o(n19780),
	.a(n19779),
	.b(n19778));
   na02f06 U21799 (.o(n23479),
	.a(n18951),
	.b(n18950));
   ao22f02 U21800 (.o(n18950),
	.a(n18960),
	.b(west_input_NIB_storage_data_f_2__30_),
	.c(n18828),
	.d(west_input_NIB_storage_data_f_1__30_));
   ao22f02 U21801 (.o(n18951),
	.a(FE_RN_5),
	.b(west_input_NIB_storage_data_f_3__30_),
	.c(FE_OFN27_n18974),
	.d(west_input_NIB_storage_data_f_0__30_));
   no03f10 U21802 (.o(n22827),
	.a(n19314),
	.b(n19313),
	.c(n19312));
   na02f04 U21804 (.o(n18368),
	.a(n18370),
	.b(n18369));
   na02f10 U21805 (.o(n23501),
	.a(n19266),
	.b(n19265));
   na02f04 U21806 (.o(n18508),
	.a(n18510),
	.b(n18509));
   na02f10 U21807 (.o(n23302),
	.a(n19212),
	.b(n19211));
   in01f08 U21808 (.o(n23325),
	.a(n18776));
   ao22f08 U21809 (.o(n19276),
	.a(FE_OFN24777_n19932),
	.b(east_input_NIB_storage_data_f_0__47_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__47_));
   ao22f08 U21810 (.o(n19277),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__47_),
	.c(FE_OFN24800_n20506),
	.d(east_input_NIB_storage_data_f_3__47_));
   ao22f10 U21811 (.o(n18909),
	.a(FE_RN_64),
	.b(west_input_NIB_storage_data_f_3__51_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__51_));
   na02f20 U21812 (.o(n23331),
	.a(n19148),
	.b(n19149));
   ao22f20 U21813 (.o(n19149),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__53_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__53_));
   oa12f20 U21814 (.o(n19351),
	.a(n19349),
	.b(n19350),
	.c(n20506));
   ao22f20 U21815 (.o(n18184),
	.a(n18828),
	.b(west_input_NIB_storage_data_f_1__55_),
	.c(FE_OFN27_n18974),
	.d(west_input_NIB_storage_data_f_0__55_));
   ao22f10 U21816 (.o(n19342),
	.a(FE_OFN24780_n19932),
	.b(east_input_NIB_storage_data_f_0__56_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__56_));
   in01f10 U21817 (.o(n18658),
	.a(n18654));
   na02f10 U21818 (.o(n18178),
	.a(n18960),
	.b(west_input_NIB_storage_data_f_2__59_));
   ao22f10 U21819 (.o(n19331),
	.a(FE_OFN24780_n19932),
	.b(east_input_NIB_storage_data_f_0__59_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__59_));
   no03f10 U21820 (.o(n22896),
	.a(n18228),
	.b(n18226),
	.c(n18230));
   na02f10 U21821 (.o(n23510),
	.a(n19190),
	.b(n19189));
   no02f01 U21822 (.o(n22941),
	.a(proc_output_space_yummy_f),
	.b(n22061));
   na02f02 U21823 (.o(n18524),
	.a(n20556),
	.b(n18525));
   no02f04 U21824 (.o(n18521),
	.a(n18523),
	.b(n18522));
   na02f04 U21825 (.o(n18522),
	.a(n20551),
	.b(n20552));
   in01f01 U21826 (.o(n18523),
	.a(n20553));
   no03f04 U21827 (.o(n20552),
	.a(reset),
	.b(n20548),
	.c(n20547));
   oa12f04 U21828 (.o(n20559),
	.a(n18205),
	.b(n18206),
	.c(n18202));
   in01m02 U21829 (.o(n18202),
	.a(n18203));
   no02m02 U21830 (.o(n18203),
	.a(n20237),
	.b(n18204));
   no02f02 U21831 (.o(n25179),
	.a(n25176),
	.b(n25175));
   na03f06 U21832 (.o(n25173),
	.a(n25171),
	.b(n25170),
	.c(n25169));
   no02f02 U21833 (.o(n18429),
	.a(n25160),
	.b(n25161));
   no03f02 U21834 (.o(n25161),
	.a(n25155),
	.b(n25154),
	.c(n25156));
   na02s02 U21835 (.o(n25491),
	.a(west_output_space_valid_f),
	.b(n25436));
   oa22f02 U21836 (.o(n19458),
	.a(n19453),
	.b(n22771),
	.c(n19452),
	.d(n19481));
   in01f02 U21837 (.o(n25106),
	.a(n25124));
   na02f04 U21838 (.o(n25090),
	.a(n25089),
	.b(n25088));
   in01f04 U21839 (.o(n18526),
	.a(n18240));
   oa22f04 U21840 (.o(n20479),
	.a(n20478),
	.b(n20477),
	.c(n25084),
	.d(n20476));
   no02f02 U21841 (.o(n18283),
	.a(n18285),
	.b(n18284));
   in01m01 U21842 (.o(n18284),
	.a(n20470));
   oa12f02 U21843 (.o(n20468),
	.a(n21661),
	.b(FE_OFN25975_n21666),
	.c(n25124));
   in01s01 U21844 (.o(n18456),
	.a(n18457));
   no03f03 U21845 (.o(n18452),
	.a(n18453),
	.b(n25094),
	.c(n25128));
   ao22f02 U21846 (.o(n18453),
	.a(n20462),
	.b(n25129),
	.c(FE_OFN366_n17753),
	.d(n25132));
   ao12f06 U21847 (.o(n18624),
	.a(n20338),
	.b(n18626),
	.c(n18057));
   no02f06 U21848 (.o(n18626),
	.a(n20342),
	.b(n18627));
   na02f04 U21849 (.o(n20341),
	.a(n20340),
	.b(n18078));
   no02f04 U21850 (.o(n18078),
	.a(n17758),
	.b(n18079));
   na02m02 U21851 (.o(n18569),
	.a(n20343),
	.b(n24973));
   oa12f04 U21852 (.o(n24981),
	.a(FE_OFN428_n22902),
	.b(n24954),
	.c(n23482));
   ao22f02 U21853 (.o(n19942),
	.a(FE_RN_69),
	.b(east_input_NIB_storage_data_f_1__29_),
	.c(n19400),
	.d(east_input_NIB_storage_data_f_3__29_));
   ao22f02 U21854 (.o(n19943),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__29_),
	.c(FE_OFN24777_n19932),
	.d(east_input_NIB_storage_data_f_0__29_));
   ao22f02 U21855 (.o(n19939),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__28_),
	.c(n19400),
	.d(east_input_NIB_storage_data_f_3__28_));
   ao22f02 U21856 (.o(n19938),
	.a(FE_OFN24777_n19932),
	.b(east_input_NIB_storage_data_f_0__28_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__28_));
   oa22f01 U21857 (.o(n21904),
	.a(n21900),
	.b(n21570),
	.c(n21899),
	.d(n21154));
   oa12s01 U21858 (.o(n21154),
	.a(n21152),
	.b(n21153),
	.c(n21570));
   ao22s01 U21859 (.o(n20771),
	.a(east_input_control_count_f_4_),
	.b(n21577),
	.c(n20770),
	.d(n21576));
   ao22f02 U21860 (.o(n19940),
	.a(FE_OFN24777_n19932),
	.b(east_input_NIB_storage_data_f_0__24_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__24_));
   ao22m02 U21861 (.o(n19944),
	.a(FE_OFN24777_n19932),
	.b(east_input_NIB_storage_data_f_0__23_),
	.c(n19400),
	.d(east_input_NIB_storage_data_f_3__23_));
   ao22f02 U21862 (.o(n19945),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__23_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__23_));
   oa22f01 U21863 (.o(n21903),
	.a(n21158),
	.b(n21899),
	.c(n21900),
	.d(n21157));
   oa12f02 U21864 (.o(n20622),
	.a(n19448),
	.b(east_input_control_thanks_all_f),
	.c(n19449));
   ao12f02 U21865 (.o(n18196),
	.a(n18598),
	.b(n18601),
	.c(n26008));
   na02f06 U21866 (.o(n23949),
	.a(n19900),
	.b(n19899));
   ao22f02 U21867 (.o(n19906),
	.a(FE_OFN51_n19193),
	.b(north_input_NIB_storage_data_f_3__26_),
	.c(FE_OFN24770_n19075),
	.d(north_input_NIB_storage_data_f_0__26_));
   oa22s01 U21868 (.o(n21890),
	.a(n21887),
	.b(n20716),
	.c(n21886),
	.d(n20715));
   ao22f02 U21869 (.o(n19903),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__25_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__25_));
   ao22f02 U21870 (.o(n19904),
	.a(FE_OFN51_n19193),
	.b(north_input_NIB_storage_data_f_3__25_),
	.c(FE_OFN24770_n19075),
	.d(north_input_NIB_storage_data_f_0__25_));
   ao22f02 U21871 (.o(n19907),
	.a(FE_RN_11),
	.b(north_input_NIB_storage_data_f_2__23_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__23_));
   ao12s01 U21872 (.o(n25280),
	.a(n25283),
	.b(n25279),
	.c(n25288));
   ao12f01 U21873 (.o(n25275),
	.a(FE_OFN25600_reset),
	.b(n25274),
	.c(n25288));
   oa12f02 U21874 (.o(n25398),
	.a(FE_OFN570_n25395),
	.b(n25397),
	.c(n25396));
   ao22f02 U21875 (.o(n19993),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__29_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__29_));
   ao22f02 U21876 (.o(n19996),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__28_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__28_));
   ao22f03 U21877 (.o(n19997),
	.a(FE_OFN28_n18974),
	.b(west_input_NIB_storage_data_f_0__28_),
	.c(n24466),
	.d(west_input_NIB_storage_data_f_2__28_));
   ao12s01 U21878 (.o(n21380),
	.a(n25227),
	.b(n21379),
	.c(west_input_control_count_f_5_));
   na02f06 U21879 (.o(n23525),
	.a(n19990),
	.b(n19989));
   na02f06 U21880 (.o(n23533),
	.a(n19988),
	.b(n19987));
   ao22f02 U21881 (.o(n19995),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__24_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__24_));
   ao22f03 U21882 (.o(n19994),
	.a(FE_OFN24764_n18960),
	.b(west_input_NIB_storage_data_f_2__24_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__24_));
   no02s01 U21883 (.o(n20624),
	.a(west_input_control_count_f_1_),
	.b(west_input_control_count_f_2_));
   ao22f02 U21884 (.o(n19998),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__23_),
	.c(FE_OFN24764_n18960),
	.d(west_input_NIB_storage_data_f_2__23_));
   ao22m02 U21885 (.o(n19979),
	.a(n18127),
	.b(west_input_NIB_storage_data_f_0__22_),
	.c(FE_OFN24764_n18960),
	.d(west_input_NIB_storage_data_f_2__22_));
   na02m01 U21886 (.o(n18639),
	.a(FE_OFN573_n25463),
	.b(FE_OCPN25903_west_input_NIB_head_ptr_f_0));
   na02s01 U21887 (.o(n18635),
	.a(FE_OFN25598_reset),
	.b(n25378));
   ao22s01 U21888 (.o(n25382),
	.a(west_input_NIB_elements_in_array_f_1_),
	.b(n25381),
	.c(n25380),
	.d(n25379));
   na02s01 U21889 (.o(n18637),
	.a(FE_OFN25598_reset),
	.b(n17784));
   oa12f02 U21890 (.o(n20620),
	.a(n19862),
	.b(proc_input_control_thanks_all_f),
	.c(n19863));
   na02f02 U21891 (.o(n20052),
	.a(n20051),
	.b(n20050));
   na02f02 U21892 (.o(n20024),
	.a(n20020),
	.b(n20019));
   na04f08 U21894 (.o(n20102),
	.a(n20101),
	.b(n20100),
	.c(n20099),
	.d(n20098));
   ao22f02 U21895 (.o(n20093),
	.a(FE_OCPN25933_n24342),
	.b(proc_input_NIB_storage_data_f_0__24_),
	.c(n17743),
	.d(proc_input_NIB_storage_data_f_4__24_));
   na02f10 U21896 (.o(n25469),
	.a(thanksIn_P),
	.b(n25978));
   na03f06 U21897 (.o(n25149),
	.a(n18105),
	.b(n17789),
	.c(thanksIn_P));
   ao22m02 U21898 (.o(n19967),
	.a(FE_OCPN25941_n24965),
	.b(south_input_NIB_storage_data_f_3__28_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__28_));
   ao22m02 U21899 (.o(n19961),
	.a(n21365),
	.b(south_input_NIB_storage_data_f_2__25_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__25_));
   ao22m02 U21900 (.o(n19970),
	.a(n24472),
	.b(south_input_NIB_storage_data_f_0__24_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__24_));
   ao22f02 U21901 (.o(n19969),
	.a(FE_OCPN25941_n24965),
	.b(south_input_NIB_storage_data_f_3__24_),
	.c(n17782),
	.d(south_input_NIB_storage_data_f_2__24_));
   in01s01 U21902 (.o(n18609),
	.a(n18610));
   in01s01 U21903 (.o(n18611),
	.a(n25344));
   na02s01 U21904 (.o(n18613),
	.a(FE_OFN575_n25463),
	.b(n25269));
   na02f03 U21905 (.o(n19473),
	.a(south_output_current_route_connection_2_),
	.b(n19911));
   oa12f02 U21906 (.o(n25135),
	.a(n25134),
	.b(north_output_current_route_connection_1_),
	.c(north_output_current_route_connection_2_));
   in01f02 U21907 (.o(n18576),
	.a(n18577));
   na02f04 U21908 (.o(n18572),
	.a(FE_RN_1),
	.b(n18573));
   no02f01 U21909 (.o(north_input_control_N52),
	.a(n21898),
	.b(n22060));
   no02f02 U21910 (.o(proc_input_control_N51),
	.a(n22935),
	.b(proc_input_control_N41));
   na02f02 U21912 (.o(n22903),
	.a(proc_input_control_N41),
	.b(n22934));
   ao12f08 U21913 (.o(n18251),
	.a(n19647),
	.b(n19153),
	.c(n19154));
   in01f02 U21914 (.o(n18424),
	.a(proc_input_NIB_storage_data_f_15__57_));
   no02f08 U21915 (.o(n20374),
	.a(myLocX_f_7_),
	.b(n22826));
   no02f06 U21916 (.o(n20375),
	.a(myLocX_f_6_),
	.b(n22865));
   no02f02 U21917 (.o(n20382),
	.a(n20374),
	.b(n25096));
   na02m02 U21918 (.o(n19816),
	.a(n19815),
	.b(n19814));
   no04f10 U21919 (.o(n19730),
	.a(n19729),
	.b(n19728),
	.c(n19727),
	.d(n19726));
   no02f10 U21920 (.o(n20300),
	.a(n19236),
	.b(n20391));
   na02f10 U21921 (.o(n18177),
	.a(n25516),
	.b(n19622));
   na02f06 U21922 (.o(n18797),
	.a(FE_OFN24742_n18683),
	.b(south_input_NIB_storage_data_f_1__30_));
   ao22f08 U21923 (.o(n18489),
	.a(proc_input_NIB_storage_data_f_10__35_),
	.b(FE_OCPN25952_n18039),
	.c(proc_input_NIB_storage_data_f_11__35_),
	.d(FE_OCPN25914_n19547));
   in01f02 U21924 (.o(n18566),
	.a(proc_input_NIB_storage_data_f_3__35_));
   ao22f08 U21925 (.o(n18704),
	.a(FE_OCPN25943_n24965),
	.b(south_input_NIB_storage_data_f_3__36_),
	.c(n24165),
	.d(south_input_NIB_storage_data_f_2__36_));
   ao22f06 U21926 (.o(n18842),
	.a(n18960),
	.b(west_input_NIB_storage_data_f_2__43_),
	.c(n18828),
	.d(west_input_NIB_storage_data_f_1__43_));
   ao22f06 U21927 (.o(n18831),
	.a(FE_OCPN25810_n18959),
	.b(west_input_NIB_storage_data_f_3__44_),
	.c(FE_OFN27_n18974),
	.d(west_input_NIB_storage_data_f_0__44_));
   ao22f06 U21928 (.o(n18158),
	.a(proc_input_NIB_storage_data_f_15__56_),
	.b(FE_OCPN25947_n19595),
	.c(proc_input_NIB_storage_data_f_8__56_),
	.d(FE_OFN170_n24343));
   ao22f06 U21929 (.o(n18416),
	.a(proc_input_NIB_storage_data_f_3__57_),
	.b(n19707),
	.c(proc_input_NIB_storage_data_f_8__57_),
	.d(FE_OFN170_n24343));
   ao22f06 U21930 (.o(n19604),
	.a(FE_OCPN25841_n24342),
	.b(proc_input_NIB_storage_data_f_0__63_),
	.c(proc_input_NIB_storage_data_f_15__63_),
	.d(FE_OCPN25947_n19595));
   na02f06 U21931 (.o(n19814),
	.a(myLocY_f_5_),
	.b(n22851));
   in01f10 U21932 (.o(n19647),
	.a(myChipID_f_2_));
   in01f20 U21933 (.o(n19666),
	.a(myChipID_f_3_));
   no02f02 U21934 (.o(n20383),
	.a(n20380),
	.b(FE_OFN946_n25096));
   na04f04 U21935 (.o(n20363),
	.a(FE_OFN428_n22902),
	.b(n20362),
	.c(n20378),
	.d(n20361));
   na02m02 U21936 (.o(n20385),
	.a(n20382),
	.b(n20376));
   in01f02 U21937 (.o(n20445),
	.a(n20443));
   na02s02 U21938 (.o(n20204),
	.a(n18422),
	.b(n19738));
   oa12f02 U21939 (.o(n19884),
	.a(n19880),
	.b(n19881),
	.c(n20181));
   ao12f02 U21940 (.o(n19880),
	.a(n19879),
	.b(n20229),
	.c(n18441));
   no02m02 U21941 (.o(n18441),
	.a(n18439),
	.b(n20186));
   in01f01 U21942 (.o(n18444),
	.a(n19802));
   na03f04 U21943 (.o(n20296),
	.a(n20176),
	.b(n20175),
	.c(n20174));
   in01f02 U21944 (.o(n20269),
	.a(n24992));
   ao22f10 U21945 (.o(n18919),
	.a(n18910),
	.b(myChipID_f_2_),
	.c(n19594),
	.d(n21696));
   na02f04 U21947 (.o(n20270),
	.a(n25247),
	.b(n19828));
   in01f02 U21948 (.o(n18340),
	.a(south_input_NIB_storage_data_f_0__22_));
   in01f01 U21950 (.o(n25022),
	.a(n25018));
   in01s01 U21951 (.o(n18338),
	.a(south_input_NIB_storage_data_f_0__2_));
   in01s01 U21952 (.o(n18346),
	.a(south_input_NIB_storage_data_f_2__3_));
   in01s01 U21953 (.o(n18336),
	.a(south_input_NIB_storage_data_f_0__5_));
   na02f10 U21954 (.o(n18725),
	.a(FE_RN_55),
	.b(south_input_NIB_storage_data_f_1__40_));
   na02f10 U21955 (.o(n18621),
	.a(south_input_NIB_storage_data_f_2__40_),
	.b(n24208));
   ao12f01 U21956 (.o(n24042),
	.a(n18563),
	.b(FE_OFN165_n24129),
	.c(proc_input_NIB_storage_data_f_1__3_));
   in01s01 U21957 (.o(n18564),
	.a(proc_input_NIB_storage_data_f_3__3_));
   in01s01 U21958 (.o(n18562),
	.a(proc_input_NIB_storage_data_f_3__8_));
   ao22f01 U21959 (.o(n21797),
	.a(FE_OFN168_n24343),
	.b(proc_input_NIB_storage_data_f_8__9_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__9_));
   ao22f02 U21960 (.o(n21771),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__10_),
	.c(FE_OCPN25834_n),
	.d(proc_input_NIB_storage_data_f_0__10_));
   ao22f01 U21961 (.o(n24108),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__11_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__11_));
   ao22f01 U21962 (.o(n24109),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__11_),
	.c(proc_input_NIB_storage_data_f_5__11_),
	.d(FE_RN_49));
   ao22f01 U21963 (.o(n24114),
	.a(FE_OCPN25814_FE_OFN186_n24453),
	.b(proc_input_NIB_storage_data_f_2__11_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__11_));
   ao22f01 U21964 (.o(n24268),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__13_),
	.c(FE_RN_51),
	.d(proc_input_NIB_storage_data_f_1__13_));
   ao22f01 U21965 (.o(n24269),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__13_),
	.c(FE_OCPN25834_n),
	.d(proc_input_NIB_storage_data_f_0__13_));
   ao22f01 U21966 (.o(n24247),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__14_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__14_));
   ao22f01 U21967 (.o(n24228),
	.a(proc_input_NIB_storage_data_f_13__15_),
	.b(FE_OFN25604_n19530),
	.c(proc_input_NIB_storage_data_f_5__15_),
	.d(FE_RN_49));
   ao22f02 U21968 (.o(n24451),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__16_),
	.c(n21740),
	.d(proc_input_NIB_storage_data_f_0__16_));
   ao22f01 U21969 (.o(n24458),
	.a(proc_input_NIB_storage_data_f_13__16_),
	.b(n24454),
	.c(proc_input_NIB_storage_data_f_5__16_),
	.d(FE_RN_49));
   ao22f01 U21970 (.o(n24154),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__17_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__17_));
   in01s01 U21971 (.o(n18560),
	.a(proc_input_NIB_storage_data_f_3__17_));
   ao22f01 U21972 (.o(n24385),
	.a(FE_OCPN25909_n19547),
	.b(proc_input_NIB_storage_data_f_11__18_),
	.c(proc_input_NIB_storage_data_f_3__18_),
	.d(n17754));
   ao22f01 U21973 (.o(n24383),
	.a(proc_input_NIB_storage_data_f_7__18_),
	.b(FE_OFN20_n17779),
	.c(proc_input_NIB_storage_data_f_5__18_),
	.d(FE_RN_49));
   ao22f01 U21974 (.o(n24381),
	.a(FE_OCPN25814_FE_OFN186_n24453),
	.b(proc_input_NIB_storage_data_f_2__18_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__18_));
   ao22f01 U21975 (.o(n24205),
	.a(proc_input_NIB_storage_data_f_10__19_),
	.b(FE_OCPN25954_n18039),
	.c(proc_input_NIB_storage_data_f_5__19_),
	.d(FE_RN_49));
   ao22f01 U21976 (.o(n24204),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__19_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__19_));
   ao22f01 U21977 (.o(n24202),
	.a(FE_RN_51),
	.b(proc_input_NIB_storage_data_f_1__19_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__19_));
   ao22f01 U21978 (.o(n24177),
	.a(proc_input_NIB_storage_data_f_13__20_),
	.b(n24454),
	.c(proc_input_NIB_storage_data_f_3__20_),
	.d(n21768));
   ao22f01 U21979 (.o(n24183),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__20_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__20_));
   ao22f01 U21980 (.o(n24312),
	.a(FE_OFN25693_n19503),
	.b(proc_input_NIB_storage_data_f_6__21_),
	.c(FE_OFN165_n24129),
	.d(proc_input_NIB_storage_data_f_1__21_));
   ao22f01 U21981 (.o(n24317),
	.a(proc_input_NIB_storage_data_f_15__21_),
	.b(FE_OFN25635_n19595),
	.c(proc_input_NIB_storage_data_f_5__21_),
	.d(n18077));
   ao22f02 U21982 (.o(n19779),
	.a(FE_OCPN25933_n24342),
	.b(proc_input_NIB_storage_data_f_0__30_),
	.c(n24455),
	.d(proc_input_NIB_storage_data_f_11__30_));
   ao22f02 U21983 (.o(n19778),
	.a(FE_OFN156_n24129),
	.b(proc_input_NIB_storage_data_f_1__30_),
	.c(n24343),
	.d(proc_input_NIB_storage_data_f_8__30_));
   ao22f02 U21984 (.o(n19760),
	.a(FE_OCPN25969_n19500),
	.b(proc_input_NIB_storage_data_f_12__31_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__31_));
   ao22m02 U21985 (.o(n19746),
	.a(n18038),
	.b(proc_input_NIB_storage_data_f_10__32_),
	.c(FE_OCPN25933_n24342),
	.d(proc_input_NIB_storage_data_f_0__32_));
   ao22f02 U21986 (.o(n19752),
	.a(n19705),
	.b(proc_input_NIB_storage_data_f_9__32_),
	.c(FE_OFN169_n24343),
	.d(proc_input_NIB_storage_data_f_8__32_));
   ao22f02 U21987 (.o(n19753),
	.a(n19709),
	.b(proc_input_NIB_storage_data_f_3__32_),
	.c(FE_OFN25674_n18033),
	.d(proc_input_NIB_storage_data_f_11__32_));
   ao22f01 U21988 (.o(n21854),
	.a(FE_RN_38),
	.b(proc_input_NIB_storage_data_f_2__33_),
	.c(n17742),
	.d(proc_input_NIB_storage_data_f_4__33_));
   ao22f06 U21989 (.o(n19555),
	.a(n19705),
	.b(proc_input_NIB_storage_data_f_9__34_),
	.c(n18037),
	.d(proc_input_NIB_storage_data_f_10__34_));
   ao22f06 U21990 (.o(n19556),
	.a(proc_input_NIB_storage_data_f_0__34_),
	.b(FE_OCPN25933_n24342),
	.c(proc_input_NIB_storage_data_f_15__34_),
	.d(FE_OFN25636_n19595));
   ao22f04 U21991 (.o(n19553),
	.a(FE_OFN25687_n19500),
	.b(proc_input_NIB_storage_data_f_12__34_),
	.c(FE_OFN25674_n18033),
	.d(proc_input_NIB_storage_data_f_11__34_));
   na02f08 U21992 (.o(n18979),
	.a(n18127),
	.b(west_input_NIB_storage_data_f_0__37_));
   na02f10 U21993 (.o(n18719),
	.a(FE_OFN24742_n18683),
	.b(south_input_NIB_storage_data_f_1__41_));
   na02f08 U21994 (.o(n18718),
	.a(FE_OFN25648_n18762),
	.b(south_input_NIB_storage_data_f_2__41_));
   ao22f04 U21995 (.o(n18520),
	.a(proc_input_NIB_storage_data_f_15__45_),
	.b(FE_OFN25634_n19595),
	.c(proc_input_NIB_storage_data_f_14__45_),
	.d(n19769));
   ao22f20 U21996 (.o(n19585),
	.a(FE_OFN24803_n19500),
	.b(proc_input_NIB_storage_data_f_12__51_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__51_));
   ao22f20 U21997 (.o(n20642),
	.a(FE_OFN24763_n18960),
	.b(west_input_NIB_storage_data_f_2__57_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__57_));
   in01f02 U21998 (.o(n18143),
	.a(south_input_NIB_storage_data_f_2__58_));
   na02s01 U21999 (.o(n18204),
	.a(n21672),
	.b(FE_OFN24833_n25232));
   in01f01 U22000 (.o(n20225),
	.a(n20224));
   in01f10 U22001 (.o(n19346),
	.a(n22889));
   ao22f10 U22002 (.o(n19407),
	.a(n23540),
	.b(myChipID_f_10_),
	.c(n19647),
	.d(n19394));
   no02f01 U22003 (.o(n25162),
	.a(FE_OFN5_reset),
	.b(west_output_current_route_connection_2_));
   na02f02 U22004 (.o(n25088),
	.a(FE_OFN428_n22902),
	.b(n25087));
   in01f02 U22005 (.o(n18492),
	.a(n20151));
   na02m20 U22006 (.o(n25127),
	.a(north_output_current_route_connection_0_),
	.b(n25130));
   no02f06 U22007 (.o(n20478),
	.a(n25087),
	.b(n18527));
   in01f03 U22008 (.o(n18273),
	.a(n20472));
   in01s01 U22009 (.o(n18138),
	.a(n19886));
   ao12f01 U22010 (.o(n25303),
	.a(n25405),
	.b(n25301),
	.c(proc_output_control_planned_f));
   no02f20 U22011 (.o(n25406),
	.a(n20475),
	.b(n20474));
   na02f02 U22012 (.o(n25404),
	.a(n24998),
	.b(n24997));
   oa12m02 U22013 (.o(n20515),
	.a(validIn_E),
	.b(n20514),
	.c(n20513));
   na02s01 U22014 (.o(n18598),
	.a(n18599),
	.b(FE_OFN25596_reset));
   na02s01 U22015 (.o(n20491),
	.a(south_output_space_yummy_f),
	.b(n20480));
   oa22s01 U22016 (.o(n19910),
	.a(north_input_control_thanks_all_f),
	.b(north_input_control_tail_last_f),
	.c(north_input_control_count_one_f),
	.d(n20648));
   no03m02 U22018 (.o(n20254),
	.a(n20242),
	.b(n20241),
	.c(n20240));
   in01f01 U22019 (.o(n18633),
	.a(n20128));
   ao22f02 U22020 (.o(n20084),
	.a(n19709),
	.b(proc_input_NIB_storage_data_f_3__29_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__29_));
   ao22f01 U22021 (.o(n20086),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__29_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__29_));
   ao22f02 U22022 (.o(n20087),
	.a(n24060),
	.b(proc_input_NIB_storage_data_f_9__29_),
	.c(n24343),
	.d(proc_input_NIB_storage_data_f_8__29_));
   ao22f02 U22023 (.o(n20088),
	.a(FE_OFN25637_n19595),
	.b(proc_input_NIB_storage_data_f_15__29_),
	.c(n17743),
	.d(proc_input_NIB_storage_data_f_4__29_));
   ao22f02 U22024 (.o(n20063),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__28_),
	.c(n20097),
	.d(proc_input_NIB_storage_data_f_15__28_));
   ao22f04 U22025 (.o(n20065),
	.a(n21739),
	.b(proc_input_NIB_storage_data_f_12__28_),
	.c(FE_OFN191_n24454),
	.d(proc_input_NIB_storage_data_f_13__28_));
   ao22f02 U22026 (.o(n20064),
	.a(FE_OCPN25823_n21745),
	.b(proc_input_NIB_storage_data_f_2__28_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__28_));
   ao22f02 U22027 (.o(n20067),
	.a(n24060),
	.b(proc_input_NIB_storage_data_f_9__28_),
	.c(n18051),
	.d(proc_input_NIB_storage_data_f_10__28_));
   ao22f02 U22028 (.o(n20068),
	.a(FE_OFN169_n24343),
	.b(proc_input_NIB_storage_data_f_8__28_),
	.c(n17744),
	.d(proc_input_NIB_storage_data_f_4__28_));
   ao22m02 U22029 (.o(n20051),
	.a(FE_OCPN25823_n21745),
	.b(proc_input_NIB_storage_data_f_2__27_),
	.c(n19769),
	.d(proc_input_NIB_storage_data_f_14__27_));
   na02f02 U22030 (.o(n20060),
	.a(n20055),
	.b(n20054));
   ao22f02 U22031 (.o(n20054),
	.a(n21768),
	.b(proc_input_NIB_storage_data_f_3__27_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__27_));
   ao22f02 U22032 (.o(n20055),
	.a(FE_OCPN25933_n24342),
	.b(proc_input_NIB_storage_data_f_0__27_),
	.c(FE_OCPN25915_n19547),
	.d(proc_input_NIB_storage_data_f_11__27_));
   ao22m02 U22033 (.o(n20020),
	.a(proc_input_NIB_storage_data_f_7__26_),
	.b(FE_OFN20_n17779),
	.c(proc_input_NIB_storage_data_f_5__26_),
	.d(FE_RN_49));
   ao22m02 U22034 (.o(n20019),
	.a(n17747),
	.b(proc_input_NIB_storage_data_f_12__26_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__26_));
   ao22f02 U22035 (.o(n20026),
	.a(FE_OCPN25951_n18039),
	.b(proc_input_NIB_storage_data_f_10__26_),
	.c(FE_OFN25604_n19530),
	.d(proc_input_NIB_storage_data_f_13__26_));
   ao22f02 U22036 (.o(n20022),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__26_),
	.c(n19709),
	.d(proc_input_NIB_storage_data_f_3__26_));
   ao22m02 U22037 (.o(n20034),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__25_),
	.c(FE_OFN20_n17779),
	.d(proc_input_NIB_storage_data_f_7__25_));
   ao22f02 U22038 (.o(n20101),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__24_),
	.c(FE_OFN156_n24129),
	.d(proc_input_NIB_storage_data_f_1__24_));
   ao22m02 U22039 (.o(n20094),
	.a(FE_OFN25604_n19530),
	.b(proc_input_NIB_storage_data_f_13__24_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__24_));
   ao22f02 U22040 (.o(n20095),
	.a(n17747),
	.b(proc_input_NIB_storage_data_f_12__24_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__24_));
   ao22f02 U22041 (.o(n20075),
	.a(n17747),
	.b(proc_input_NIB_storage_data_f_12__23_),
	.c(FE_OFN25604_n19530),
	.d(proc_input_NIB_storage_data_f_13__23_));
   ao22f02 U22042 (.o(n20073),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__23_),
	.c(FE_OFN25637_n19595),
	.d(proc_input_NIB_storage_data_f_15__23_));
   ao22m02 U22043 (.o(n20009),
	.a(FE_OCPN25826_n21745),
	.b(proc_input_NIB_storage_data_f_2__22_),
	.c(FE_OCPN25933_n24342),
	.d(proc_input_NIB_storage_data_f_0__22_));
   in01f01 U22045 (.o(n19028),
	.a(n19031));
   no02f01 U22047 (.o(n21385),
	.a(south_input_control_count_f_0_),
	.b(south_input_control_count_f_1_));
   na02s01 U22048 (.o(n25242),
	.a(n25241),
	.b(n25240));
   no04f20 U22049 (.o(n19833),
	.a(n19836),
	.b(n18736),
	.c(n18117),
	.d(n18116));
   no03f04 U22050 (.o(n25033),
	.a(n25017),
	.b(n17759),
	.c(n20501));
   no02f04 U22051 (.o(n25023),
	.a(n25022),
	.b(n25021));
   na02f01 U22052 (.o(n25021),
	.a(n25020),
	.b(n18543));
   no02f06 U22053 (.o(n22957),
	.a(FE_OFN25601_reset),
	.b(east_input_NIB_tail_ptr_f_0_));
   na02f10 U22054 (.o(n24920),
	.a(validIn_E),
	.b(east_input_NIB_tail_ptr_f_0_));
   oa12s01 U22055 (.o(n25769),
	.a(n25766),
	.b(n25768),
	.c(n25767));
   ao22s01 U22056 (.o(n25766),
	.a(ec_thanks_e_to_s_reg),
	.b(n25757),
	.c(ec_thanks_n_to_s_reg),
	.d(n25765));
   ao22m01 U22057 (.o(n24032),
	.a(n25294),
	.b(n24031),
	.c(FE_OFN79_n20501),
	.d(n24030));
   ao22f01 U22058 (.o(n22225),
	.a(FE_OFN526_n24731),
	.b(FE_OFN136_n23623),
	.c(FE_OFN94_n21695),
	.d(n23622));
   ao22f01 U22059 (.o(n22229),
	.a(FE_OFN111_n22773),
	.b(FE_OFN140_n23959),
	.c(FE_OFN94_n21695),
	.d(n23958));
   in01s01 U22060 (.o(n18262),
	.a(n18263));
   in01s01 U22061 (.o(n18265),
	.a(n18266));
   ao22f20 U22062 (.o(n18939),
	.a(FE_OFN24763_n18960),
	.b(west_input_NIB_storage_data_f_2__56_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__56_));
   in01s01 U22063 (.o(n18256),
	.a(n18257));
   in01s01 U22064 (.o(n18259),
	.a(n18260));
   no02f06 U22065 (.o(n19415),
	.a(n19479),
	.b(n19476));
   no02f02 U22066 (.o(n18430),
	.a(FE_OFN250_n25152),
	.b(n25177));
   no02s01 U22067 (.o(n25460),
	.a(n25459),
	.b(n25455));
   ao12s01 U22068 (.o(n25461),
	.a(west_output_space_count_f_0_),
	.b(n25491),
	.c(n25454));
   ao12s01 U22069 (.o(n25444),
	.a(n25439),
	.b(n25459),
	.c(west_output_space_count_f_1_));
   na02f04 U22070 (.o(n25092),
	.a(n25124),
	.b(n25091));
   no02f06 U22072 (.o(n25309),
	.a(n25026),
	.b(n25025));
   na02f02 U22074 (.o(n25418),
	.a(n25414),
	.b(n25413));
   in01f10 U22075 (.o(n25038),
	.a(proc_output_current_route_connection_1_));
   no02f01 U22076 (.o(n25409),
	.a(FE_OFN259_n25295),
	.b(n25294));
   no03f02 U22077 (.o(n21906),
	.a(n21905),
	.b(n21904),
	.c(n21903));
   in01s01 U22078 (.o(n18573),
	.a(n18574));
   no03s01 U22079 (.o(n25328),
	.a(east_input_NIB_elements_in_array_f_0_),
	.b(east_input_NIB_elements_in_array_f_1_),
	.c(validIn_E));
   ao22s01 U22080 (.o(n25319),
	.a(east_input_NIB_elements_in_array_f_0_),
	.b(validIn_E),
	.c(n25316),
	.d(n25315));
   na02f03 U22081 (.o(n20503),
	.a(n25498),
	.b(n19911));
   ao12s01 U22082 (.o(n20500),
	.a(n20491),
	.b(n20495),
	.c(south_output_space_count_f_2_));
   ao22s01 U22083 (.o(n20499),
	.a(n20495),
	.b(n20494),
	.c(n20493),
	.d(n20492));
   ao12s01 U22084 (.o(n20498),
	.a(n20496),
	.b(south_output_space_count_f_0_),
	.c(n20497));
   oa12s01 U22085 (.o(n20484),
	.a(south_output_space_count_f_1_),
	.b(south_output_space_count_f_0_),
	.c(n20493));
   in01s01 U22086 (.o(n20710),
	.a(n20709));
   no03f01 U22087 (.o(n20699),
	.a(north_input_control_count_f_0_),
	.b(north_input_control_count_f_1_),
	.c(n20648));
   ao22s01 U22088 (.o(n20616),
	.a(n20630),
	.b(west_input_control_count_f_1_),
	.c(n20629),
	.d(n20615));
   in01f10 U22089 (.o(n20566),
	.a(west_input_control_thanks_all_f));
   na02s01 U22090 (.o(n20132),
	.a(west_input_NIB_elements_in_array_f_2_),
	.b(FE_OFN25598_reset));
   no02f06 U22091 (.o(n18631),
	.a(n18502),
	.b(n18507));
   in01s01 U22092 (.o(n18502),
	.a(n18503));
   na02f01 U22093 (.o(n18503),
	.a(n18632),
	.b(n18633));
   oa22s01 U22094 (.o(n22391),
	.a(east_output_space_count_f_0_),
	.b(n22390),
	.c(n22389),
	.d(n22388));
   na04f01 U22095 (.o(n22900),
	.a(n22899),
	.b(n22898),
	.c(n22897),
	.d(FE_OFN947_n25096));
   in01s01 U22097 (.o(n18128),
	.a(n18129));
   no03s01 U22098 (.o(n25375),
	.a(n25370),
	.b(n25374),
	.c(n25369));
   ao12s01 U22099 (.o(n25359),
	.a(n25369),
	.b(n25374),
	.c(north_output_space_count_f_1_));
   oa12f10 U22100 (.o(n20590),
	.a(n18794),
	.b(south_input_control_thanks_all_f),
	.c(n18795));
   in01s01 U22101 (.o(n18607),
	.a(n18643));
   na02s01 U22102 (.o(n18643),
	.a(n18645),
	.b(n18644));
   in01s01 U22103 (.o(n18645),
	.a(n19489));
   na02s01 U22104 (.o(n19483),
	.a(south_input_NIB_elements_in_array_f_2_),
	.b(FE_OFN575_n25463));
   no02f06 U22105 (.o(n18615),
	.a(n18616),
	.b(n18399));
   oa22s01 U22106 (.o(n22081),
	.a(proc_output_space_count_f_0_),
	.b(n22080),
	.c(n22941),
	.d(n22079));
   na02f02 U22107 (.o(n22069),
	.a(n22941),
	.b(n22079));
   na02f06 U22108 (.o(n25049),
	.a(n24999),
	.b(n25302));
   na03f04 U22109 (.o(n18493),
	.a(n18495),
	.b(n25311),
	.c(n18494));
   oa12s01 U22110 (.o(n25983),
	.a(FE_OFN574_n25463),
	.b(n25978),
	.c(n25977));
   na02f01 U22111 (.o(n25973),
	.a(proc_input_NIB_tail_ptr_f_1_),
	.b(proc_input_NIB_tail_ptr_f_0_));
   na03f20 U22112 (.o(n24921),
	.a(east_input_NIB_tail_ptr_f_1_),
	.b(FE_OFN25596_reset),
	.c(n25862));
   oa12s01 U22113 (.o(ec_out_3_),
	.a(n25794),
	.b(ec_cfg_11_),
	.c(n25795));
   na02f02 U22115 (.o(n24660),
	.a(n24659),
	.b(n24658));
   oa12f01 U22116 (.o(FE_OFN881_dataOut_P_1),
	.a(n24669),
	.b(n24670),
	.c(FE_OFN524_n24728));
   na02f02 U22117 (.o(n24668),
	.a(n24667),
	.b(n24666));
   ao22m02 U22118 (.o(n24667),
	.a(n25294),
	.b(n24663),
	.c(FE_OFN79_n20501),
	.d(FE_OFN221_n24662));
   oa12f01 U22119 (.o(FE_OFN1072_dataOut_P_2),
	.a(n24649),
	.b(n24701),
	.c(FE_OFN524_n24728));
   na02f02 U22120 (.o(n24648),
	.a(n24647),
	.b(n24646));
   ao22f01 U22121 (.o(n24647),
	.a(n17787),
	.b(n24694),
	.c(FE_OFN79_n20501),
	.d(n24693));
   oa12f01 U22122 (.o(FE_OFN1070_dataOut_P_3),
	.a(n24653),
	.b(n24692),
	.c(FE_OFN524_n24728));
   na02f02 U22123 (.o(n24652),
	.a(n24651),
	.b(n24650));
   oa12f01 U22124 (.o(FE_OFN1068_dataOut_P_4),
	.a(n24657),
	.b(FE_OFN937_n24710),
	.c(FE_OFN524_n24728));
   na02f02 U22125 (.o(n24656),
	.a(n24655),
	.b(n24654));
   na02f02 U22126 (.o(n23980),
	.a(n23979),
	.b(n23978));
   ao22f01 U22127 (.o(n23978),
	.a(n25294),
	.b(n23977),
	.c(n17787),
	.d(n23976));
   oa12m02 U22128 (.o(FE_OFN879_dataOut_P_6),
	.a(n24017),
	.b(n24018),
	.c(FE_OFN524_n24728));
   ao22f01 U22129 (.o(n24015),
	.a(n25295),
	.b(FE_OFN485_n24011),
	.c(FE_OFN79_n20501),
	.d(FE_OFN146_n24010));
   oa12f01 U22130 (.o(FE_OFN1064_dataOut_P_7),
	.a(n23566),
	.b(n23567),
	.c(FE_OFN524_n24728));
   ao22f01 U22131 (.o(n23564),
	.a(n25294),
	.b(FE_OFN473_n23560),
	.c(FE_OFN79_n20501),
	.d(FE_OFN130_n23559));
   oa12f01 U22132 (.o(FE_OFN1062_dataOut_P_8),
	.a(n23153),
	.b(n23154),
	.c(FE_OFN524_n24728));
   ao22f01 U22133 (.o(n23150),
	.a(n17787),
	.b(n23149),
	.c(FE_OFN79_n20501),
	.d(FE_OFN116_n23148));
   oa12f01 U22134 (.o(FE_OFN25731_dataOut_P_9),
	.a(n23575),
	.b(FE_OFN923_n23576),
	.c(FE_OFN524_n24728));
   ao22f01 U22135 (.o(n23573),
	.a(FE_OFN257_n25294),
	.b(n23569),
	.c(FE_OFN79_n20501),
	.d(n23568));
   oa12f01 U22136 (.o(FE_OFN877_dataOut_P_10),
	.a(n23584),
	.b(n23585),
	.c(FE_OFN523_n24728));
   oa12f01 U22137 (.o(FE_OFN875_dataOut_P_11),
	.a(n24583),
	.b(FE_OFN201_n24584),
	.c(FE_OFN524_n24728));
   na02f02 U22139 (.o(n24591),
	.a(n24590),
	.b(n24589));
   oa12f01 U22140 (.o(FE_OFN873_dataOut_P_13),
	.a(n24605),
	.b(n24606),
	.c(FE_OFN524_n24728));
   na02f02 U22141 (.o(n24604),
	.a(n24603),
	.b(n24602));
   ao22f01 U22142 (.o(n24602),
	.a(n25294),
	.b(FE_OFN499_n24601),
	.c(FE_OFN79_n20501),
	.d(FE_OFN203_n24600));
   oa12f01 U22143 (.o(FE_OFN1056_dataOut_P_14),
	.a(n24682),
	.b(n24683),
	.c(n24728));
   na02f02 U22144 (.o(n24681),
	.a(n24680),
	.b(n24679));
   oa12f01 U22145 (.o(FE_OFN871_dataOut_P_15),
	.a(n24614),
	.b(n24627),
	.c(n24728));
   na02f02 U22146 (.o(n24613),
	.a(n24612),
	.b(n24611));
   ao22f01 U22147 (.o(n24612),
	.a(n17787),
	.b(n24620),
	.c(FE_OFN79_n20501),
	.d(FE_OFN207_n24619));
   oa12m02 U22148 (.o(FE_OFN869_dataOut_P_16),
	.a(n24610),
	.b(FE_OFN215_n24636),
	.c(FE_OFN524_n24728));
   na02f02 U22149 (.o(n24609),
	.a(n24608),
	.b(n24607));
   ao22f01 U22150 (.o(n24607),
	.a(n17787),
	.b(n24631),
	.c(FE_OFN79_n20501),
	.d(FE_OFN211_n24630));
   oa12f01 U22151 (.o(FE_OFN867_dataOut_P_17),
	.a(n24618),
	.b(FE_OFN219_n24645),
	.c(FE_OFN524_n24728));
   na02f02 U22152 (.o(n24617),
	.a(n24616),
	.b(n24615));
   ao22f01 U22153 (.o(n24616),
	.a(n17787),
	.b(n24638),
	.c(FE_OFN79_n20501),
	.d(FE_OFN217_n24637));
   oa12f01 U22154 (.o(FE_OFN1054_dataOut_P_18),
	.a(n24758),
	.b(n24759),
	.c(FE_OFN524_n24728));
   na02f02 U22155 (.o(n24757),
	.a(n24756),
	.b(n24755));
   ao22f01 U22156 (.o(n24755),
	.a(FE_OFN257_n25294),
	.b(n24754),
	.c(FE_OFN79_n20501),
	.d(n24752));
   oa12f01 U22157 (.o(FE_OFN865_dataOut_P_19),
	.a(n24597),
	.b(n24749),
	.c(FE_OFN524_n24728));
   na02f02 U22158 (.o(n24596),
	.a(n24595),
	.b(n24594));
   oa12f01 U22159 (.o(FE_OFN863_dataOut_P_20),
	.a(n24727),
	.b(FE_OFN235_n24729),
	.c(n24728));
   na02f02 U22160 (.o(n24726),
	.a(n24725),
	.b(n24724));
   oa12f01 U22161 (.o(FE_OFN861_dataOut_P_21),
	.a(n24718),
	.b(FE_OFN233_n24719),
	.c(FE_OFN524_n24728));
   na02f02 U22162 (.o(n24717),
	.a(n24716),
	.b(n24715));
   no02f01 U22163 (.o(n23990),
	.a(n23989),
	.b(n23988));
   oa22f01 U22164 (.o(n23988),
	.a(FE_OFN483_n23987),
	.b(n25411),
	.c(n23986),
	.d(n20501));
   ao22m01 U22165 (.o(n23624),
	.a(FE_OFN79_n20501),
	.b(FE_OFN136_n23623),
	.c(n17787),
	.d(n23622));
   na03f02 U22166 (.o(FE_OFN853_dataOut_P_25),
	.a(n23539),
	.b(n23538),
	.c(n23537));
   na03f04 U22167 (.o(dataOut_P_26_),
	.a(n23531),
	.b(n23530),
	.c(n23529));
   na03f04 U22168 (.o(dataOut_P_27_),
	.a(n23523),
	.b(n23522),
	.c(n23521));
   ao22m01 U22169 (.o(n23960),
	.a(FE_OFN79_n20501),
	.b(FE_OFN140_n23959),
	.c(n17787),
	.d(n23958));
   na03f02 U22170 (.o(dataOut_P_30_),
	.a(n23485),
	.b(n23484),
	.c(n23483));
   ao22f01 U22171 (.o(n23484),
	.a(n17787),
	.b(n23481),
	.c(n25294),
	.d(n23480));
   no02f02 U22172 (.o(n23039),
	.a(n23038),
	.b(n23037));
   oa12f01 U22173 (.o(FE_OFN843_dataOut_P_33),
	.a(n24026),
	.b(FE_OFN153_n24027),
	.c(FE_OFN524_n24728));
   oa12f01 U22174 (.o(FE_OFN25707_dataOut_P_35),
	.a(n22841),
	.b(n18097),
	.c(n24728));
   no02f01 U22175 (.o(n22849),
	.a(n22848),
	.b(n22847));
   na03f01 U22176 (.o(FE_OFN827_dataOut_P_43),
	.a(n23499),
	.b(n23498),
	.c(n23497));
   na03f06 U22177 (.o(dataOut_P_44_),
	.a(n23507),
	.b(n23506),
	.c(n23505));
   na03f04 U22178 (.o(dataOut_P_45_),
	.a(n23307),
	.b(n23306),
	.c(n23305));
   na03f03 U22179 (.o(dataOut_P_46_),
	.a(n23299),
	.b(n23298),
	.c(n23297));
   na03f03 U22180 (.o(dataOut_P_47_),
	.a(n23329),
	.b(n23328),
	.c(n23327));
   na03m02 U22181 (.o(dataOut_P_51_),
	.a(n23339),
	.b(n23338),
	.c(n23337));
   oa12f01 U22182 (.o(dataOut_P_52_),
	.a(n23636),
	.b(n18103),
	.c(FE_OFN24730_n));
   na03m02 U22183 (.o(dataOut_P_53_),
	.a(n23336),
	.b(n23335),
	.c(n23334));
   na03f02 U22184 (.o(dataOut_P_55_),
	.a(n23321),
	.b(n23320),
	.c(n23319));
   oa12f02 U22185 (.o(dataOut_P_58_),
	.a(n23593),
	.b(FE_OFN134_n23594),
	.c(FE_OFN524_n24728));
   na03f02 U22186 (.o(dataOut_P_59_),
	.a(n23350),
	.b(n23349),
	.c(n23348));
   oa12f02 U22187 (.o(dataOut_P_61_),
	.a(n24008),
	.b(n24009),
	.c(FE_OFN524_n24728));
   no02f01 U22188 (.o(n24008),
	.a(n24007),
	.b(n24006));
   no02f01 U22189 (.o(n22895),
	.a(n22894),
	.b(n22893));
   oa22f01 U22190 (.o(n22893),
	.a(n22892),
	.b(n25029),
	.c(n22891),
	.d(n25411));
   na03m02 U22191 (.o(dataOut_P_63_),
	.a(n23515),
	.b(n23514),
	.c(n23513));
   oa12f01 U22192 (.o(FE_OFN809_dataOut_W_0),
	.a(n24738),
	.b(FE_OFN239_n24739),
	.c(FE_OFN25878_n19446));
   oa12f01 U22193 (.o(FE_OFN807_dataOut_W_1),
	.a(n24551),
	.b(n24670),
	.c(FE_OFN25878_n19446));
   ao22f01 U22194 (.o(n24549),
	.a(n17755),
	.b(n24663),
	.c(FE_OFN111_n22773),
	.d(FE_OFN221_n24662));
   oa12f01 U22195 (.o(FE_OFN1050_dataOut_W_2),
	.a(n24700),
	.b(n24701),
	.c(FE_OFN25878_n19446));
   oa12f01 U22196 (.o(FE_OFN1048_dataOut_W_3),
	.a(n24691),
	.b(n24692),
	.c(FE_OFN394_n19446));
   oa12f01 U22197 (.o(FE_OFN1046_dataOut_W_4),
	.a(n24709),
	.b(FE_OFN937_n24710),
	.c(FE_OFN25878_n19446));
   oa12f01 U22198 (.o(FE_OFN1044_dataOut_W_5),
	.a(n22366),
	.b(n23982),
	.c(FE_OFN25878_n19446));
   oa12f01 U22199 (.o(FE_OFN805_dataOut_W_6),
	.a(n22358),
	.b(n24018),
	.c(FE_OFN25878_n19446));
   oa12f01 U22200 (.o(FE_OFN1042_dataOut_W_7),
	.a(n22346),
	.b(n23567),
	.c(FE_OFN394_n19446));
   oa12f01 U22201 (.o(FE_OFN1040_dataOut_W_8),
	.a(n22362),
	.b(n23154),
	.c(FE_OFN25878_n19446));
   oa12f01 U22202 (.o(FE_OFN25729_dataOut_W_9),
	.a(n22350),
	.b(FE_OFN923_n23576),
	.c(FE_OFN394_n19446));
   oa12f01 U22203 (.o(FE_OFN803_dataOut_W_10),
	.a(n22370),
	.b(n23585),
	.c(FE_OFN25879_n19446));
   oa12f01 U22204 (.o(FE_OFN801_dataOut_W_11),
	.a(n24559),
	.b(FE_OFN201_n24584),
	.c(FE_OFN25878_n19446));
   oa12f01 U22205 (.o(FE_OFN1036_dataOut_W_12),
	.a(n24575),
	.b(n24593),
	.c(FE_OFN25880_n19446));
   ao22f01 U22207 (.o(n24536),
	.a(n17755),
	.b(FE_OFN499_n24601),
	.c(FE_OFN111_n22773),
	.d(FE_OFN203_n24600));
   oa12f01 U22208 (.o(FE_OFN1034_dataOut_W_14),
	.a(n24567),
	.b(n24683),
	.c(FE_OFN25881_n19446));
   oa12f01 U22209 (.o(FE_OFN797_dataOut_W_15),
	.a(n24626),
	.b(n24627),
	.c(FE_OFN25880_n19446));
   oa12f01 U22210 (.o(FE_OFN795_dataOut_W_16),
	.a(n24635),
	.b(FE_OFN215_n24636),
	.c(FE_OFN25878_n19446));
   oa12f01 U22211 (.o(FE_OFN793_dataOut_W_17),
	.a(n24644),
	.b(FE_OFN219_n24645),
	.c(FE_OFN25878_n19446));
   ao22f01 U22213 (.o(n24544),
	.a(n17755),
	.b(n24754),
	.c(FE_OFN111_n22773),
	.d(n24752));
   oa12f01 U22214 (.o(FE_OFN791_dataOut_W_19),
	.a(n24543),
	.b(n24749),
	.c(FE_OFN25878_n19446));
   ao22f01 U22215 (.o(n24540),
	.a(n17755),
	.b(n24742),
	.c(FE_OFN111_n22773),
	.d(FE_OFN242_n24744));
   oa12m02 U22216 (.o(FE_OFN789_dataOut_W_20),
	.a(n24563),
	.b(FE_OFN235_n24729),
	.c(FE_OFN25880_n19446));
   oa12f02 U22218 (.o(dataOut_W_22_),
	.a(n21548),
	.b(FE_OFN144_n23991),
	.c(FE_OFN25880_n19446));
   no02f01 U22219 (.o(n21548),
	.a(n21547),
	.b(n21546));
   ao22f01 U22220 (.o(n21707),
	.a(FE_OFN526_n24731),
	.b(n23478),
	.c(n17755),
	.d(n23480));
   no02f02 U22221 (.o(n22659),
	.a(n22658),
	.b(n22657));
   oa12f01 U22222 (.o(FE_OFN769_dataOut_W_33),
	.a(n22354),
	.b(FE_OFN153_n24027),
	.c(FE_OFN25878_n19446));
   no02f01 U22223 (.o(n22776),
	.a(n22775),
	.b(n22774));
   oa12f01 U22224 (.o(FE_OFN25701_dataOut_W_35),
	.a(n22525),
	.b(n18097),
	.c(FE_OFN25880_n19446));
   no02f01 U22225 (.o(n22525),
	.a(n22524),
	.b(n22523));
   no02f01 U22226 (.o(n22770),
	.a(n22769),
	.b(n22768));
   no02f01 U22227 (.o(n22759),
	.a(n22758),
	.b(n22757));
   oa22f01 U22228 (.o(n22758),
	.a(n22852),
	.b(FE_OFN110_n22771),
	.c(n17751),
	.d(n21695));
   na02f01 U22229 (.o(FE_OFN362_dataOut_W_40),
	.a(n21495),
	.b(n21494));
   no02f01 U22230 (.o(n21495),
	.a(n21493),
	.b(n21492));
   na02f02 U22231 (.o(dataOut_W_41_),
	.a(n21526),
	.b(n21525));
   no02f01 U22232 (.o(n21526),
	.a(n21524),
	.b(n21523));
   no02f02 U22233 (.o(n22628),
	.a(n22627),
	.b(n22626));
   no02f01 U22234 (.o(n22662),
	.a(n22661),
	.b(n22660));
   no02f01 U22235 (.o(n22491),
	.a(n22490),
	.b(n22489));
   oa12f01 U22236 (.o(dataOut_W_52_),
	.a(n22220),
	.b(n18103),
	.c(FE_OFN25883_n19446));
   ao22f01 U22237 (.o(n22217),
	.a(FE_OFN111_n22773),
	.b(n23629),
	.c(n17755),
	.d(FE_OFN479_n23631));
   oa12f01 U22238 (.o(dataOut_W_54_),
	.a(n22764),
	.b(n24000),
	.c(FE_OFN25883_n19446));
   no02f01 U22239 (.o(n22764),
	.a(n22763),
	.b(n22762));
   no02f01 U22240 (.o(n22539),
	.a(n22538),
	.b(n22537));
   no02f02 U22241 (.o(n22767),
	.a(FE_OFN424_n22766),
	.b(n22765));
   oa12f01 U22242 (.o(FE_OFN733_dataOut_S_0),
	.a(n24487),
	.b(FE_OFN239_n24739),
	.c(FE_OFN25652_n25499));
   oa12f01 U22243 (.o(FE_OFN731_dataOut_S_1),
	.a(n24507),
	.b(n24670),
	.c(FE_OFN25652_n25499));
   oa12f01 U22244 (.o(FE_OFN1026_dataOut_S_2),
	.a(n24555),
	.b(n24701),
	.c(FE_OFN266_n25499));
   oa12f01 U22245 (.o(FE_OFN1024_dataOut_S_3),
	.a(n24519),
	.b(n24692),
	.c(FE_OFN25652_n25499));
   oa12f01 U22246 (.o(FE_OFN1022_dataOut_S_4),
	.a(n24523),
	.b(FE_OFN937_n24710),
	.c(FE_OFN266_n25499));
   oa12f01 U22247 (.o(FE_OFN1020_dataOut_S_5),
	.a(n22601),
	.b(n23982),
	.c(FE_OFN266_n25499));
   oa12f01 U22248 (.o(FE_OFN729_dataOut_S_6),
	.a(n22617),
	.b(n24018),
	.c(FE_OFN266_n25499));
   oa12f01 U22249 (.o(FE_OFN1018_dataOut_S_7),
	.a(n22609),
	.b(n23567),
	.c(FE_OFN25652_n25499));
   oa12f01 U22250 (.o(FE_OFN1016_dataOut_S_8),
	.a(n22605),
	.b(n23154),
	.c(FE_OFN25652_n25499));
   oa12m02 U22251 (.o(FE_OFN1014_dataOut_S_9),
	.a(n22613),
	.b(FE_OFN923_n23576),
	.c(FE_OFN25652_n25499));
   oa12f01 U22252 (.o(FE_OFN727_dataOut_S_10),
	.a(n22621),
	.b(n23585),
	.c(FE_OFN266_n25499));
   oa12f01 U22253 (.o(FE_OFN725_dataOut_S_11),
	.a(n24499),
	.b(FE_OFN201_n24584),
	.c(FE_OFN266_n25499));
   oa12f01 U22254 (.o(FE_OFN1012_dataOut_S_12),
	.a(n24495),
	.b(n24593),
	.c(FE_OFN266_n25499));
   oa12f01 U22255 (.o(FE_OFN723_dataOut_S_13),
	.a(n24511),
	.b(n24606),
	.c(FE_OFN266_n25499));
   oa12f01 U22256 (.o(FE_OFN1010_dataOut_S_14),
	.a(n24503),
	.b(n24683),
	.c(FE_OFN266_n25499));
   oa12m02 U22257 (.o(FE_OFN721_dataOut_S_15),
	.a(n24515),
	.b(n24627),
	.c(FE_OFN266_n25499));
   oa12f01 U22258 (.o(FE_OFN719_dataOut_S_16),
	.a(n24491),
	.b(FE_OFN215_n24636),
	.c(FE_OFN25652_n25499));
   oa12f01 U22259 (.o(FE_OFN717_dataOut_S_17),
	.a(n24527),
	.b(FE_OFN219_n24645),
	.c(FE_OFN266_n25499));
   oa12m02 U22261 (.o(FE_OFN715_dataOut_S_19),
	.a(n24748),
	.b(n24749),
	.c(FE_OFN266_n25499));
   oa12f01 U22262 (.o(FE_OFN713_dataOut_S_20),
	.a(n24535),
	.b(FE_OFN235_n24729),
	.c(FE_OFN266_n25499));
   oa12f01 U22263 (.o(FE_OFN711_dataOut_S_21),
	.a(n24531),
	.b(FE_OFN233_n24719),
	.c(FE_OFN25652_n25499));
   no02f02 U22264 (.o(n21635),
	.a(n21634),
	.b(n21633));
   oa22f01 U22265 (.o(n21633),
	.a(FE_OFN483_n23987),
	.b(FE_OFN92_n21667),
	.c(n23986),
	.d(n22518));
   oa12f01 U22266 (.o(FE_OFN693_dataOut_S_33),
	.a(n22434),
	.b(FE_OFN153_n24027),
	.c(FE_OFN266_n25499));
   oa12f01 U22267 (.o(FE_OFN689_dataOut_S_35),
	.a(n21625),
	.b(n18097),
	.c(FE_OFN25651_n25499));
   oa22f01 U22268 (.o(n21624),
	.a(n22835),
	.b(n22518),
	.c(n22838),
	.d(n22517));
   oa12m02 U22269 (.o(dataOut_S_52_),
	.a(n22516),
	.b(n18103),
	.c(FE_OFN25652_n25499));
   ao22f01 U22270 (.o(n22513),
	.a(FE_OFN396_n19493),
	.b(n23630),
	.c(FE_OFN93_n21667),
	.d(FE_OFN479_n23631));
   oa22f01 U22271 (.o(n21617),
	.a(n23589),
	.b(FE_OFN540_n24743),
	.c(n21616),
	.d(FE_OFN247_n24982));
   ao22f01 U22272 (.o(n25502),
	.a(FE_OFN105_n22517),
	.b(n18028),
	.c(FE_OFN577_n25498),
	.d(n25497));
   na02f02 U22274 (.o(n24370),
	.a(n24369),
	.b(n24368));
   ao22f01 U22275 (.o(n24368),
	.a(FE_OFN42_n19022),
	.b(n24734),
	.c(n19020),
	.d(FE_OFN530_n24733));
   oa12f02 U22276 (.o(dataOut_E_1_),
	.a(n24341),
	.b(n24670),
	.c(FE_OFN25895_n25395));
   na02f01 U22277 (.o(n24340),
	.a(n24339),
	.b(n24338));
   ao22f01 U22278 (.o(n24338),
	.a(n19019),
	.b(n24665),
	.c(FE_OFN42_n19022),
	.d(FE_OFN223_n24664));
   oa12f01 U22279 (.o(FE_OFN1004_dataOut_E_2),
	.a(n24337),
	.b(n24701),
	.c(FE_OFN25892_n25395));
   na02f02 U22280 (.o(n24336),
	.a(n24335),
	.b(n24334));
   ao22f01 U22281 (.o(n24334),
	.a(n19019),
	.b(n24696),
	.c(n19020),
	.d(FE_OFN513_n24695));
   oa12f01 U22282 (.o(FE_OFN1002_dataOut_E_3),
	.a(n24059),
	.b(n24692),
	.c(FE_OFN25895_n25395));
   na02f02 U22283 (.o(n24058),
	.a(n24057),
	.b(n24056));
   ao22f01 U22284 (.o(n24056),
	.a(FE_OFN42_n19022),
	.b(n24687),
	.c(n19020),
	.d(n24686));
   oa12f01 U22285 (.o(FE_OFN1000_dataOut_E_4),
	.a(n24443),
	.b(FE_OFN937_n24710),
	.c(FE_OFN25892_n25395));
   na02f02 U22286 (.o(n24442),
	.a(n24441),
	.b(n24440));
   ao22f01 U22287 (.o(n24441),
	.a(n19022),
	.b(n24703),
	.c(n19020),
	.d(FE_OFN515_n24702));
   na02f01 U22289 (.o(n21324),
	.a(n21323),
	.b(n21322));
   ao22f01 U22290 (.o(n21322),
	.a(FE_OFN42_n19022),
	.b(n23976),
	.c(n19020),
	.d(n23977));
   oa12f01 U22291 (.o(FE_OFN655_dataOut_E_6),
	.a(n21375),
	.b(n24018),
	.c(FE_OFN25895_n25395));
   ao22f01 U22292 (.o(n21372),
	.a(FE_OFN42_n19022),
	.b(n24012),
	.c(n19020),
	.d(FE_OFN487_n24013));
   oa12f01 U22293 (.o(FE_OFN996_dataOut_E_7),
	.a(n21837),
	.b(n23567),
	.c(FE_OFN25895_n25395));
   na02f02 U22294 (.o(n21836),
	.a(n21835),
	.b(n21834));
   ao22f01 U22295 (.o(n21835),
	.a(n19017),
	.b(FE_OFN130_n23559),
	.c(n19020),
	.d(FE_OFN473_n23560));
   ao22f01 U22296 (.o(n21765),
	.a(n19019),
	.b(n23147),
	.c(n19020),
	.d(n23146));
   oa12f01 U22297 (.o(FE_OFN992_dataOut_E_9),
	.a(n21885),
	.b(FE_OFN923_n23576),
	.c(FE_OFN25895_n25395));
   na02f02 U22298 (.o(n21884),
	.a(n21883),
	.b(n21882));
   ao22f01 U22299 (.o(n21883),
	.a(n19017),
	.b(n23568),
	.c(n19020),
	.d(n23569));
   oa12f01 U22300 (.o(FE_OFN653_dataOut_E_10),
	.a(n21790),
	.b(n23585),
	.c(n25395));
   na02f02 U22301 (.o(n21789),
	.a(n21788),
	.b(n21787));
   ao22f01 U22302 (.o(n21788),
	.a(n19022),
	.b(n23577),
	.c(n19020),
	.d(FE_OFN477_n23578));
   oa12m02 U22303 (.o(FE_OFN651_dataOut_E_11),
	.a(n24435),
	.b(FE_OFN201_n24584),
	.c(FE_OFN25895_n25395));
   na02f02 U22304 (.o(n24434),
	.a(n24433),
	.b(n24432));
   ao22f01 U22305 (.o(n24433),
	.a(FE_OFN42_n19022),
	.b(n24576),
	.c(n19020),
	.d(FE_OFN493_n24577));
   oa12m02 U22306 (.o(FE_OFN990_dataOut_E_12),
	.a(n24431),
	.b(n24593),
	.c(FE_OFN25891_n25395));
   na02f02 U22307 (.o(n24430),
	.a(n24429),
	.b(n24428));
   ao22f01 U22308 (.o(n24429),
	.a(n19022),
	.b(n24585),
	.c(n19020),
	.d(FE_OFN497_n24586));
   oa12f01 U22309 (.o(FE_OFN649_dataOut_E_13),
	.a(n24427),
	.b(n24606),
	.c(FE_OFN25892_n25395));
   na02f02 U22310 (.o(n24426),
	.a(n24425),
	.b(n24424));
   ao22f01 U22311 (.o(n24424),
	.a(n19017),
	.b(FE_OFN203_n24600),
	.c(n19020),
	.d(FE_OFN499_n24601));
   oa12f01 U22312 (.o(FE_OFN988_dataOut_E_14),
	.a(n24423),
	.b(n24683),
	.c(n25395));
   na02f02 U22313 (.o(n24422),
	.a(n24421),
	.b(n24420));
   ao22f01 U22314 (.o(n24421),
	.a(FE_OFN42_n19022),
	.b(n24675),
	.c(n19020),
	.d(n24676));
   oa12f01 U22315 (.o(FE_OFN647_dataOut_E_15),
	.a(n24415),
	.b(n24627),
	.c(FE_OFN25891_n25395));
   na02f02 U22316 (.o(n24414),
	.a(n24413),
	.b(n24412));
   ao22f01 U22317 (.o(n24412),
	.a(n19019),
	.b(n24622),
	.c(n19020),
	.d(n24621));
   oa12f02 U22318 (.o(dataOut_E_16_),
	.a(n24483),
	.b(FE_OFN215_n24636),
	.c(FE_OFN25895_n25395));
   oa12f01 U22321 (.o(FE_OFN641_dataOut_E_19),
	.a(n24379),
	.b(n24749),
	.c(FE_OFN25892_n25395));
   ao22f01 U22322 (.o(n24377),
	.a(n19019),
	.b(n24741),
	.c(FE_OFN42_n19022),
	.d(n24740));
   oa12f01 U22323 (.o(FE_OFN639_dataOut_E_20),
	.a(n24375),
	.b(FE_OFN235_n24729),
	.c(n25395));
   ao22f01 U22324 (.o(n24372),
	.a(FE_OFN42_n19022),
	.b(n24722),
	.c(n19020),
	.d(FE_OFN521_n24723));
   oa12m02 U22325 (.o(FE_OFN637_dataOut_E_21),
	.a(n24333),
	.b(FE_OFN233_n24719),
	.c(FE_OFN25895_n25395));
   ao22f01 U22326 (.o(n24331),
	.a(FE_OFN42_n19022),
	.b(n24711),
	.c(n19020),
	.d(FE_OFN517_n24712));
   oa12m02 U22327 (.o(FE_OFN25719_dataOut_E_22),
	.a(n21434),
	.b(FE_OFN144_n23991),
	.c(FE_OFN569_n25395));
   no02f02 U22328 (.o(n21434),
	.a(n21433),
	.b(n21432));
   na02f02 U22329 (.o(n21401),
	.a(n21400),
	.b(n21399));
   na02f01 U22330 (.o(n21451),
	.a(n21450),
	.b(n21449));
   na02f01 U22331 (.o(n21132),
	.a(n21131),
	.b(n21130));
   na02f02 U22332 (.o(n20967),
	.a(n20966),
	.b(n20965));
   no02f01 U22333 (.o(n21480),
	.a(n21479),
	.b(n21478));
   oa12f01 U22334 (.o(FE_OFN621_dataOut_E_33),
	.a(n21877),
	.b(FE_OFN153_n24027),
	.c(FE_OFN25892_n25395));
   ao22f01 U22335 (.o(n21874),
	.a(FE_OFN42_n19022),
	.b(n24021),
	.c(n19020),
	.d(FE_OFN491_n24022));
   oa12f02 U22336 (.o(dataOut_E_35_),
	.a(n20915),
	.b(n18097),
	.c(FE_OFN569_n25395));
   oa22f01 U22337 (.o(n20761),
	.a(n22852),
	.b(n21672),
	.c(n17751),
	.d(FE_OFN412_n21671));
   oa12f01 U22338 (.o(dataOut_E_52_),
	.a(n21171),
	.b(n18103),
	.c(FE_OFN25895_n25395));
   no02f01 U22339 (.o(n20794),
	.a(n20793),
	.b(n20792));
   oa12f01 U22340 (.o(FE_OFN342_dataOut_N_0),
	.a(n24419),
	.b(FE_OFN239_n24739),
	.c(n21666));
   oa12f01 U22342 (.o(FE_OFN340_dataOut_N_1),
	.a(n24106),
	.b(n24670),
	.c(n21666));
   oa12m02 U22343 (.o(FE_OFN980_dataOut_N_2),
	.a(n24152),
	.b(n24701),
	.c(n21666));
   oa12f01 U22344 (.o(FE_OFN978_dataOut_N_3),
	.a(n24407),
	.b(n24692),
	.c(n21666));
   ao22f01 U22345 (.o(n24405),
	.a(FE_OFN44_n19054),
	.b(FE_OFN229_n24684),
	.c(n19057),
	.d(n24685));
   oa12f01 U22346 (.o(FE_OFN976_dataOut_N_4),
	.a(n24083),
	.b(FE_OFN937_n24710),
	.c(n21666));
   ao22f01 U22347 (.o(n24080),
	.a(FE_OFN44_n19054),
	.b(FE_OFN231_n24704),
	.c(n19057),
	.d(n24705));
   oa12f01 U22348 (.o(FE_OFN974_dataOut_N_5),
	.a(n21321),
	.b(n23982),
	.c(n21666));
   ao22f01 U22349 (.o(n21319),
	.a(FE_OFN44_n19054),
	.b(n23974),
	.c(n19057),
	.d(n23975));
   oa12f01 U22350 (.o(FE_OFN338_dataOut_N_6),
	.a(n21371),
	.b(n24018),
	.c(n21666));
   ao22f01 U22351 (.o(n21369),
	.a(FE_OFN44_n19054),
	.b(FE_OFN146_n24010),
	.c(n19057),
	.d(FE_OFN485_n24011));
   oa12f01 U22352 (.o(FE_OFN972_dataOut_N_7),
	.a(n21881),
	.b(n23567),
	.c(n21666));
   oa12f01 U22353 (.o(FE_OFN970_dataOut_N_8),
	.a(n21845),
	.b(n23154),
	.c(n21666));
   ao22f01 U22354 (.o(n21843),
	.a(FE_OFN47_n19056),
	.b(n23146),
	.c(n19057),
	.d(n23147));
   oa12f01 U22355 (.o(FE_OFN968_dataOut_N_9),
	.a(n21814),
	.b(FE_OFN923_n23576),
	.c(n21666));
   ao22f01 U22356 (.o(n21812),
	.a(FE_OFN47_n19056),
	.b(n23569),
	.c(FE_OFN44_n19054),
	.d(n23568));
   oa12f01 U22357 (.o(FE_OFN336_dataOut_N_10),
	.a(n21841),
	.b(n23585),
	.c(n21666));
   ao22f01 U22358 (.o(n21838),
	.a(FE_OFN45_n19054),
	.b(n23579),
	.c(n19057),
	.d(n23580));
   oa12m02 U22359 (.o(FE_OFN334_dataOut_N_11),
	.a(n24128),
	.b(FE_OFN201_n24584),
	.c(n21666));
   ao22f01 U22360 (.o(n24125),
	.a(FE_OFN44_n19054),
	.b(n24578),
	.c(n19057),
	.d(FE_OFN495_n24579));
   oa12m02 U22361 (.o(FE_OFN966_dataOut_N_12),
	.a(n24310),
	.b(n24593),
	.c(n21666));
   oa12f01 U22362 (.o(FE_OFN332_dataOut_N_13),
	.a(n24288),
	.b(n24606),
	.c(n21666));
   oa12f01 U22363 (.o(FE_OFN964_dataOut_N_14),
	.a(n24266),
	.b(n24683),
	.c(n21666));
   ao22f01 U22364 (.o(n24263),
	.a(n19054),
	.b(FE_OFN227_n24677),
	.c(n19057),
	.d(n24678));
   oa12f01 U22365 (.o(FE_OFN330_dataOut_N_15),
	.a(n24243),
	.b(n24627),
	.c(n21666));
   ao22f01 U22366 (.o(n24240),
	.a(n19056),
	.b(n24621),
	.c(n19057),
	.d(n24622));
   oa12f01 U22367 (.o(FE_OFN328_dataOut_N_16),
	.a(n24479),
	.b(FE_OFN215_n24636),
	.c(n21666));
   ao22f01 U22368 (.o(n24477),
	.a(FE_OFN47_n19056),
	.b(n24628),
	.c(n19057),
	.d(n24629));
   oa12f01 U22369 (.o(FE_OFN326_dataOut_N_17),
	.a(n24175),
	.b(FE_OFN219_n24645),
	.c(n21666));
   ao22f01 U22370 (.o(n24172),
	.a(n19056),
	.b(n24639),
	.c(n19057),
	.d(n24640));
   oa12m02 U22371 (.o(FE_OFN962_dataOut_N_18),
	.a(n24439),
	.b(n24759),
	.c(n21666));
   oa12f01 U22372 (.o(FE_OFN324_dataOut_N_19),
	.a(n24220),
	.b(n24749),
	.c(n21666));
   oa12m02 U22373 (.o(FE_OFN322_dataOut_N_20),
	.a(n24197),
	.b(FE_OFN235_n24729),
	.c(n21666));
   ao22f01 U22374 (.o(n24195),
	.a(n19054),
	.b(n24720),
	.c(n19057),
	.d(n24721));
   oa12m02 U22375 (.o(FE_OFN320_dataOut_N_21),
	.a(n24447),
	.b(FE_OFN233_n24719),
	.c(n21666));
   ao22f01 U22376 (.o(n21556),
	.a(n19056),
	.b(n23535),
	.c(n19054),
	.d(n23534));
   ao22f01 U22377 (.o(n21520),
	.a(n19054),
	.b(n23527),
	.c(n19059),
	.d(n23526));
   ao22f01 U22378 (.o(n21563),
	.a(n19054),
	.b(n23519),
	.c(n19059),
	.d(n23518));
   ao22f01 U22379 (.o(n21463),
	.a(n19054),
	.b(n23478),
	.c(n19056),
	.d(n23480));
   oa12f01 U22380 (.o(FE_OFN304_dataOut_N_33),
	.a(n21873),
	.b(FE_OFN153_n24027),
	.c(n21666));
   ao22f01 U22381 (.o(n21870),
	.a(n19056),
	.b(FE_OFN491_n24022),
	.c(FE_OFN366_n17753),
	.d(n24021));
   oa12m02 U22382 (.o(FE_OFN25705_dataOut_N_35),
	.a(n20918),
	.b(n18097),
	.c(FE_OFN25976_n21666));
   oa22f01 U22383 (.o(n20764),
	.a(n17751),
	.b(n25095),
	.c(n22852),
	.d(n21661));
   oa12f01 U22384 (.o(dataOut_N_52_),
	.a(n21167),
	.b(n18103),
	.c(FE_OFN25980_n21666));
   ao22f01 U22385 (.o(n21164),
	.a(FE_OFN44_n19054),
	.b(n23629),
	.c(FE_OFN47_n19056),
	.d(FE_OFN479_n23631));
   no02f01 U22386 (.o(n20751),
	.a(FE_OFN904_n20750),
	.b(n20749));
   na03f02 U22387 (.o(n20562),
	.a(FE_OFN25598_reset),
	.b(n25396),
	.c(n20546));
   oa12f02 U22388 (.o(n20561),
	.a(n18521),
	.b(n25396),
	.c(n18524));
   na02f04 U22389 (.o(n19494),
	.a(n19493),
	.b(n19911));
   na02f02 U22390 (.o(n20543),
	.a(n20537),
	.b(n20536));
   no02f01 U22391 (.o(west_output_control_N72),
	.a(n25496),
	.b(n25495));
   oa12s01 U22392 (.o(n25492),
	.a(n25491),
	.b(west_output_space_is_one_f),
	.c(west_output_space_yummy_f));
   in01f02 U22393 (.o(n18277),
	.a(n18278));
   na02f04 U22395 (.o(n18451),
	.a(n18142),
	.b(n18452));
   oa22s01 U22396 (.o(east_input_control_N48),
	.a(n21575),
	.b(n21588),
	.c(n21574),
	.d(FE_OFN906_n21586));
   ao22s01 U22397 (.o(n21574),
	.a(east_input_control_count_f_7_),
	.b(n21573),
	.c(n21572),
	.d(n21901));
   oa12f01 U22398 (.o(east_input_control_N41),
	.a(n20574),
	.b(n20575),
	.c(n21586));
   no02f02 U22399 (.o(n20527),
	.a(n20525),
	.b(n20511));
   oa12m01 U22400 (.o(south_output_space_N44),
	.a(FE_OFN25599_reset),
	.b(n20483),
	.c(n20482));
   ao12s01 U22401 (.o(n20482),
	.a(n20494),
	.b(n20489),
	.c(n20486));
   na02f01 U22402 (.o(n25273),
	.a(validOut_S),
	.b(FE_OFN25599_reset));
   oa22s01 U22403 (.o(n20739),
	.a(n21893),
	.b(north_input_control_count_f_5_),
	.c(n20736),
	.d(n21886));
   no02f01 U22404 (.o(n26009),
	.a(n20572),
	.b(n20571));
   ao22s01 U22405 (.o(n20572),
	.a(north_input_control_count_f_0_),
	.b(n21886),
	.c(n20719),
	.d(n21887));
   ao12f01 U22406 (.o(north_input_control_N51),
	.a(n26009),
	.b(FE_OFN575_n25463),
	.c(n22060));
   oa22s01 U22407 (.o(n25278),
	.a(north_input_NIB_elements_in_array_f_1_),
	.b(validIn_N),
	.c(n25288),
	.d(n25281));
   ao22s01 U22408 (.o(n25276),
	.a(n25279),
	.b(north_input_NIB_elements_in_array_f_1_),
	.c(validIn_N),
	.d(n25288));
   ao22m04 U22409 (.o(n20333),
	.a(north_input_NIB_elements_in_array_f_0_),
	.b(n25830),
	.c(validIn_N),
	.d(n25289));
   oa12f02 U22410 (.o(n25068),
	.a(FE_OFN25598_reset),
	.b(east_output_current_route_connection_2_),
	.c(n25384));
   na02f08 U22411 (.o(n19026),
	.a(n25506),
	.b(n20213));
   na02f02 U22412 (.o(n20328),
	.a(FE_OFN25598_reset),
	.b(n25384));
   ao12f01 U22414 (.o(n25233),
	.a(n25230),
	.b(FE_OFN24831_n25232),
	.c(n25231));
   ao22m01 U22415 (.o(n25229),
	.a(west_input_control_count_f_7_),
	.b(n25228),
	.c(n25227),
	.d(n25226));
   ao22m01 U22416 (.o(n23041),
	.a(west_input_control_count_f_6_),
	.b(n25227),
	.c(n23040),
	.d(n25225));
   na02f03 U22417 (.o(n18504),
	.a(n18505),
	.b(n18507));
   in01s01 U22418 (.o(n18505),
	.a(n18506));
   in01f01 U22419 (.o(n25426),
	.a(n18638));
   na02f04 U22420 (.o(n25425),
	.a(n26013),
	.b(FE_OFN24761_west_input_NIB_head_ptr_f_0));
   na02f04 U22421 (.o(n18546),
	.a(n20130),
	.b(n20131));
   na02f04 U22422 (.o(n18547),
	.a(n20133),
	.b(n20134));
   na02f04 U22423 (.o(n20130),
	.a(n20129),
	.b(n18507));
   na02f02 U22424 (.o(n25988),
	.a(n25383),
	.b(n18545));
   in01f02 U22425 (.o(n25383),
	.a(n18634));
   na02f04 U22426 (.o(n18545),
	.a(n26013),
	.b(n25382));
   in01f02 U22427 (.o(n25236),
	.a(n18636));
   no02s01 U22428 (.o(n18501),
	.a(reset),
	.b(n17784));
   no02s01 U22429 (.o(east_output_space_N47),
	.a(n25817),
	.b(east_output_space_N48));
   na02f01 U22430 (.o(east_output_space_N44),
	.a(FE_OFN25599_reset),
	.b(n22374));
   oa22m02 U22431 (.o(n22374),
	.a(east_output_space_count_f_2_),
	.b(n22376),
	.c(n22373),
	.d(n22384));
   no02s01 U22432 (.o(n22373),
	.a(n22376),
	.b(n22372));
   oa22f01 U22433 (.o(n21692),
	.a(FE_OFN428_n22902),
	.b(n21691),
	.c(n21690),
	.d(n21689));
   oa22f01 U22434 (.o(proc_input_control_N46),
	.a(FE_OFN122_n23520),
	.b(n21694),
	.c(n21641),
	.d(n21689));
   oa22f01 U22435 (.o(proc_input_control_N45),
	.a(n21649),
	.b(n21694),
	.c(n21648),
	.d(n21689));
   oa22f01 U22436 (.o(proc_input_control_N41),
	.a(n20576),
	.b(n21689),
	.c(n23991),
	.d(n21694));
   na02f10 U22437 (.o(proc_input_valid),
	.a(FE_OFN25684_n25474),
	.b(n25486));
   na03f02 U22439 (.o(n25143),
	.a(n25142),
	.b(proc_input_NIB_head_ptr_f_1_),
	.c(n25463));
   na02f04 U22440 (.o(n25144),
	.a(n25995),
	.b(n25141));
   na03f04 U22441 (.o(n20510),
	.a(n25142),
	.b(proc_input_NIB_head_ptr_f_0_),
	.c(FE_OFN573_n25463));
   na02f06 U22442 (.o(n20509),
	.a(n25995),
	.b(n20508));
   no02f10 U22443 (.o(n25995),
	.a(reset),
	.b(n25142));
   na03s01 U22444 (.o(n18594),
	.a(n18597),
	.b(n18596),
	.c(n18595));
   in01s01 U22445 (.o(n18595),
	.a(north_output_space_is_two_or_more_f));
   in01s01 U22446 (.o(n18597),
	.a(n22938));
   na03f01 U22447 (.o(north_output_space_N48),
	.a(n25815),
	.b(n17888),
	.c(n25816));
   no03f01 U22448 (.o(n20758),
	.a(n20757),
	.b(n20756),
	.c(n20755));
   no03f02 U22449 (.o(n26026),
	.a(n20565),
	.b(FE_OFN5_reset),
	.c(n20564));
   ao22s01 U22450 (.o(n20565),
	.a(south_input_control_count_f_0_),
	.b(n25250),
	.c(n20752),
	.d(n23550));
   na02f02 U22451 (.o(n2988),
	.a(n24966),
	.b(n18592));
   in01s01 U22453 (.o(n18397),
	.a(n18398));
   in01f02 U22454 (.o(n25350),
	.a(n18608));
   in01f02 U22455 (.o(n25272),
	.a(n18612));
   no02s01 U22456 (.o(proc_output_space_N47),
	.a(n25824),
	.b(proc_output_space_N48));
   oa12s01 U22457 (.o(n3093),
	.a(n23825),
	.b(FE_OFN25618_n23789),
	.c(n23827));
   na02s01 U22458 (.o(n23825),
	.a(proc_input_NIB_storage_data_f_0__63_),
	.b(FE_OFN25618_n23789));
   oa12s01 U22459 (.o(n3098),
	.a(n23794),
	.b(FE_OFN25618_n23789),
	.c(n23810));
   na02s01 U22460 (.o(n23794),
	.a(proc_input_NIB_storage_data_f_0__62_),
	.b(FE_OFN25618_n23789));
   oa12s01 U22461 (.o(n3103),
	.a(n23828),
	.b(FE_OFN25618_n23789),
	.c(n23918));
   oa12s01 U22462 (.o(n3108),
	.a(n23835),
	.b(FE_OFN25618_n23789),
	.c(n23926));
   na02s01 U22463 (.o(n23835),
	.a(proc_input_NIB_storage_data_f_0__60_),
	.b(FE_OFN25618_n23789));
   oa12s01 U22464 (.o(n3113),
	.a(n23846),
	.b(FE_OFN25618_n23789),
	.c(n23938));
   na02s01 U22465 (.o(n23846),
	.a(proc_input_NIB_storage_data_f_0__59_),
	.b(FE_OFN25618_n23789));
   oa12s01 U22466 (.o(n3118),
	.a(n23832),
	.b(FE_OFN25618_n23789),
	.c(n23936));
   na02s01 U22467 (.o(n23832),
	.a(proc_input_NIB_storage_data_f_0__58_),
	.b(FE_OFN25618_n23789));
   oa12f01 U22468 (.o(n3123),
	.a(n23852),
	.b(FE_OFN25620_n23789),
	.c(n23932));
   na02s01 U22469 (.o(n23852),
	.a(proc_input_NIB_storage_data_f_0__57_),
	.b(FE_OFN25620_n23789));
   oa12f01 U22470 (.o(n3128),
	.a(n23853),
	.b(FE_OFN25620_n23789),
	.c(n23930));
   na02f01 U22471 (.o(n23853),
	.a(proc_input_NIB_storage_data_f_0__56_),
	.b(FE_OFN25620_n23789));
   oa12f01 U22472 (.o(n3133),
	.a(n23830),
	.b(FE_OFN25620_n23789),
	.c(n23910));
   na02f01 U22473 (.o(n23830),
	.a(proc_input_NIB_storage_data_f_0__55_),
	.b(FE_OFN25620_n23789));
   oa12f01 U22474 (.o(n3138),
	.a(n23861),
	.b(FE_OFN25620_n23789),
	.c(n23924));
   na02f01 U22475 (.o(n23861),
	.a(proc_input_NIB_storage_data_f_0__54_),
	.b(FE_OFN25620_n23789));
   oa12f01 U22476 (.o(n3143),
	.a(n23845),
	.b(FE_OFN25620_n23789),
	.c(n23922));
   na02f01 U22477 (.o(n23845),
	.a(proc_input_NIB_storage_data_f_0__53_),
	.b(FE_OFN25620_n23789));
   oa12f01 U22478 (.o(n3148),
	.a(n23847),
	.b(FE_OFN25620_n23789),
	.c(n23890));
   na02f01 U22479 (.o(n23847),
	.a(proc_input_NIB_storage_data_f_0__52_),
	.b(FE_OFN25620_n23789));
   oa12s01 U22480 (.o(n3153),
	.a(n23946),
	.b(FE_OFN25618_n23789),
	.c(n23947));
   na02s01 U22481 (.o(n23946),
	.a(proc_input_NIB_storage_data_f_0__51_),
	.b(FE_OFN25618_n23789));
   oa12s01 U22482 (.o(n3158),
	.a(n23848),
	.b(FE_OFN25618_n23789),
	.c(n23903));
   na02s01 U22483 (.o(n23848),
	.a(proc_input_NIB_storage_data_f_0__50_),
	.b(FE_OFN25618_n23789));
   oa12f01 U22484 (.o(n3163),
	.a(n23849),
	.b(n25547),
	.c(n23908));
   na02f01 U22485 (.o(n23849),
	.a(proc_input_NIB_storage_data_f_0__49_),
	.b(n25547));
   oa12f01 U22486 (.o(n3168),
	.a(n23850),
	.b(n25547),
	.c(n23912));
   na02f01 U22487 (.o(n23850),
	.a(proc_input_NIB_storage_data_f_0__48_),
	.b(n25547));
   oa12f01 U22488 (.o(n3173),
	.a(n23851),
	.b(n17765),
	.c(n23914));
   na02f01 U22489 (.o(n23851),
	.a(proc_input_NIB_storage_data_f_0__47_),
	.b(n17765));
   oa12f01 U22490 (.o(n3178),
	.a(n23891),
	.b(n25547),
	.c(n23916));
   oa12f01 U22491 (.o(n3183),
	.a(n23854),
	.b(FE_OFN25622_n23789),
	.c(n23942));
   na02f01 U22492 (.o(n23854),
	.a(proc_input_NIB_storage_data_f_0__45_),
	.b(FE_OFN25622_n23789));
   oa12f01 U22493 (.o(n3188),
	.a(n23855),
	.b(FE_OFN25622_n23789),
	.c(n23920));
   na02f01 U22494 (.o(n23855),
	.a(proc_input_NIB_storage_data_f_0__44_),
	.b(FE_OFN25622_n23789));
   oa12f01 U22495 (.o(n3193),
	.a(n23805),
	.b(n17765),
	.c(n23806));
   na02f01 U22496 (.o(n23805),
	.a(proc_input_NIB_storage_data_f_0__43_),
	.b(n17765));
   oa12f01 U22497 (.o(n3198),
	.a(n23807),
	.b(n25547),
	.c(n23808));
   na02f01 U22498 (.o(n23807),
	.a(proc_input_NIB_storage_data_f_0__42_),
	.b(n25547));
   oa12f01 U22499 (.o(n3203),
	.a(n23863),
	.b(n17765),
	.c(n23928));
   na02f01 U22500 (.o(n23863),
	.a(proc_input_NIB_storage_data_f_0__41_),
	.b(n17765));
   oa12f01 U22501 (.o(n3208),
	.a(n23799),
	.b(FE_OFN25622_n23789),
	.c(n23800));
   na02f01 U22502 (.o(n23799),
	.a(proc_input_NIB_storage_data_f_0__40_),
	.b(FE_OFN25622_n23789));
   oa12f01 U22503 (.o(n3213),
	.a(n23868),
	.b(FE_OFN25619_n23789),
	.c(n23934));
   na02f01 U22504 (.o(n23868),
	.a(proc_input_NIB_storage_data_f_0__39_),
	.b(FE_OFN25619_n23789));
   oa12f01 U22505 (.o(n3218),
	.a(n23811),
	.b(n17765),
	.c(n23812));
   na02f01 U22506 (.o(n23811),
	.a(proc_input_NIB_storage_data_f_0__38_),
	.b(n17765));
   oa12f01 U22507 (.o(n3223),
	.a(n23795),
	.b(n17765),
	.c(n23796));
   na02f01 U22508 (.o(n23795),
	.a(proc_input_NIB_storage_data_f_0__37_),
	.b(n17765));
   oa12f01 U22509 (.o(n3228),
	.a(n23875),
	.b(n17765),
	.c(n23940));
   na02f01 U22510 (.o(n23875),
	.a(proc_input_NIB_storage_data_f_0__36_),
	.b(n17765));
   oa12f01 U22511 (.o(n3233),
	.a(n23876),
	.b(n17765),
	.c(n23944));
   na02f01 U22512 (.o(n23876),
	.a(proc_input_NIB_storage_data_f_0__35_),
	.b(n17765));
   oa12f01 U22513 (.o(n3238),
	.a(n23815),
	.b(n17765),
	.c(n23816));
   na02f01 U22514 (.o(n23815),
	.a(proc_input_NIB_storage_data_f_0__34_),
	.b(n17765));
   oa22f01 U22515 (.o(n25525),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_0__33_),
	.d(FE_OFN580_n25547));
   oa12f01 U22516 (.o(n3248),
	.a(n23878),
	.b(n17765),
	.c(n23905));
   na02f01 U22517 (.o(n23878),
	.a(proc_input_NIB_storage_data_f_0__32_),
	.b(n17765));
   oa12f01 U22518 (.o(n3253),
	.a(n23790),
	.b(FE_OFN25622_n23789),
	.c(n23791));
   oa12f01 U22519 (.o(n3258),
	.a(n23881),
	.b(n25547),
	.c(n23894));
   na02f01 U22520 (.o(n23881),
	.a(proc_input_NIB_storage_data_f_0__30_),
	.b(n25547));
   oa12f01 U22521 (.o(n3263),
	.a(n23803),
	.b(n25547),
	.c(n23804));
   na02s01 U22522 (.o(n23803),
	.a(proc_input_NIB_storage_data_f_0__29_),
	.b(n25547));
   oa12f01 U22523 (.o(n3268),
	.a(n23813),
	.b(FE_OFN25619_n23789),
	.c(n23814));
   na02f01 U22524 (.o(n23813),
	.a(proc_input_NIB_storage_data_f_0__28_),
	.b(FE_OFN25619_n23789));
   oa12f01 U22525 (.o(n3273),
	.a(n23821),
	.b(FE_OFN25619_n23789),
	.c(n23822));
   na02f01 U22526 (.o(n23821),
	.a(proc_input_NIB_storage_data_f_0__27_),
	.b(FE_OFN25619_n23789));
   oa12f01 U22527 (.o(n3278),
	.a(n23817),
	.b(n25547),
	.c(n23818));
   na02f01 U22528 (.o(n23817),
	.a(proc_input_NIB_storage_data_f_0__26_),
	.b(n25547));
   oa12f01 U22529 (.o(n3283),
	.a(n23801),
	.b(FE_OFN25619_n23789),
	.c(n23802));
   na02f01 U22530 (.o(n23801),
	.a(proc_input_NIB_storage_data_f_0__25_),
	.b(FE_OFN25619_n23789));
   oa12f01 U22531 (.o(n3288),
	.a(n23797),
	.b(n25547),
	.c(n23798));
   na02f01 U22532 (.o(n23797),
	.a(proc_input_NIB_storage_data_f_0__24_),
	.b(n25547));
   oa12f01 U22533 (.o(n3293),
	.a(n23792),
	.b(n17765),
	.c(n23793));
   na02f01 U22534 (.o(n23792),
	.a(proc_input_NIB_storage_data_f_0__23_),
	.b(n17765));
   oa12f01 U22535 (.o(n3298),
	.a(n23819),
	.b(FE_OFN25619_n23789),
	.c(n23820));
   na02f01 U22536 (.o(n23819),
	.a(proc_input_NIB_storage_data_f_0__22_),
	.b(FE_OFN25619_n23789));
   oa22s01 U22537 (.o(n25526),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_0__21_),
	.d(FE_OFN580_n25547));
   oa22f01 U22538 (.o(n25527),
	.a(FE_OFN25622_n23789),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_0__20_),
	.d(FE_OFN580_n25547));
   oa22s01 U22539 (.o(n25528),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_0__19_),
	.d(FE_OFN580_n25547));
   oa22s01 U22540 (.o(n25530),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_0__17_),
	.d(FE_OFN580_n25547));
   oa22f01 U22541 (.o(n25531),
	.a(FE_OFN25620_n23789),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_0__16_),
	.d(FE_OFN580_n25547));
   oa22f01 U22542 (.o(n25532),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_0__15_),
	.d(FE_OFN580_n25547));
   oa22f01 U22543 (.o(n25533),
	.a(FE_OFN25622_n23789),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_0__14_),
	.d(FE_OFN580_n25547));
   oa22s01 U22544 (.o(n25534),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_0__13_),
	.d(FE_OFN580_n25547));
   oa22f01 U22545 (.o(n25535),
	.a(FE_OFN25622_n23789),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_0__12_),
	.d(FE_OFN580_n25547));
   oa22f01 U22546 (.o(n25536),
	.a(FE_OFN25622_n23789),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_0__11_),
	.d(FE_OFN580_n25547));
   oa22s01 U22547 (.o(n25537),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_0__10_),
	.d(FE_OFN580_n25547));
   oa22s01 U22548 (.o(n25538),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_0__9_),
	.d(FE_OFN580_n25547));
   oa22s01 U22549 (.o(n25539),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_0__8_),
	.d(FE_OFN580_n25547));
   oa22s01 U22550 (.o(n25540),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_0__7_),
	.d(FE_OFN580_n25547));
   oa22s01 U22551 (.o(n25541),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_0__6_),
	.d(FE_OFN580_n25547));
   oa22s01 U22552 (.o(n25542),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_0__5_),
	.d(FE_OFN580_n25547));
   oa22f01 U22553 (.o(n25543),
	.a(FE_OFN25622_n23789),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_0__4_),
	.d(FE_OFN580_n25547));
   oa22f01 U22554 (.o(n25545),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_0__2_),
	.d(FE_OFN580_n25547));
   oa22f01 U22555 (.o(n25546),
	.a(FE_OFN25620_n23789),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_0__1_),
	.d(FE_OFN580_n25547));
   oa22f01 U22556 (.o(n25548),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_0__0_),
	.d(FE_OFN580_n25547));
   oa22s01 U22557 (.o(n25572),
	.a(n17762),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_1__0_),
	.d(n25571));
   oa12f01 U22558 (.o(n3733),
	.a(n23826),
	.b(FE_OFN272_n25595),
	.c(n23827));
   na02s01 U22559 (.o(n23826),
	.a(proc_input_NIB_storage_data_f_2__63_),
	.b(FE_OFN272_n25595));
   oa12f01 U22560 (.o(n3738),
	.a(n23786),
	.b(FE_OFN272_n25595),
	.c(n23810));
   na02s01 U22561 (.o(n23786),
	.a(proc_input_NIB_storage_data_f_2__62_),
	.b(FE_OFN272_n25595));
   oa12f01 U22562 (.o(n3743),
	.a(n23917),
	.b(FE_OFN272_n25595),
	.c(n23918));
   na02s01 U22563 (.o(n23917),
	.a(proc_input_NIB_storage_data_f_2__61_),
	.b(FE_OFN272_n25595));
   oa12f01 U22564 (.o(n3748),
	.a(n23906),
	.b(FE_OFN272_n25595),
	.c(n23926));
   na02s01 U22565 (.o(n23906),
	.a(proc_input_NIB_storage_data_f_2__60_),
	.b(FE_OFN272_n25595));
   oa12f01 U22566 (.o(n3753),
	.a(n23901),
	.b(FE_OFN272_n25595),
	.c(n23938));
   na02s01 U22567 (.o(n23901),
	.a(proc_input_NIB_storage_data_f_2__59_),
	.b(FE_OFN272_n25595));
   oa12f01 U22568 (.o(n3758),
	.a(n23899),
	.b(FE_OFN272_n25595),
	.c(n23936));
   oa12s01 U22569 (.o(n3763),
	.a(n23898),
	.b(FE_OFN272_n25595),
	.c(n23932));
   na02s01 U22570 (.o(n23898),
	.a(proc_input_NIB_storage_data_f_2__57_),
	.b(FE_OFN272_n25595));
   oa12s01 U22571 (.o(n3768),
	.a(n23897),
	.b(FE_OFN272_n25595),
	.c(n23930));
   na02s01 U22572 (.o(n23897),
	.a(proc_input_NIB_storage_data_f_2__56_),
	.b(FE_OFN272_n25595));
   oa12s01 U22573 (.o(n3773),
	.a(n23896),
	.b(FE_OFN272_n25595),
	.c(n23910));
   na02s01 U22574 (.o(n23896),
	.a(proc_input_NIB_storage_data_f_2__55_),
	.b(FE_OFN272_n25595));
   oa12f01 U22575 (.o(n3778),
	.a(n23895),
	.b(FE_OFN272_n25595),
	.c(n23924));
   na02s01 U22576 (.o(n23895),
	.a(proc_input_NIB_storage_data_f_2__54_),
	.b(FE_OFN272_n25595));
   oa12s01 U22577 (.o(n3783),
	.a(n23892),
	.b(FE_OFN272_n25595),
	.c(n23922));
   na02s01 U22578 (.o(n23892),
	.a(proc_input_NIB_storage_data_f_2__53_),
	.b(FE_OFN272_n25595));
   oa12f01 U22579 (.o(n3788),
	.a(n23889),
	.b(FE_OFN272_n25595),
	.c(n23890));
   na02s01 U22580 (.o(n23889),
	.a(proc_input_NIB_storage_data_f_2__52_),
	.b(FE_OFN272_n25595));
   oa12f01 U22581 (.o(n3793),
	.a(n23888),
	.b(FE_OFN272_n25595),
	.c(n23947));
   na02s01 U22582 (.o(n23888),
	.a(proc_input_NIB_storage_data_f_2__51_),
	.b(FE_OFN272_n25595));
   oa12f01 U22583 (.o(n3798),
	.a(n23887),
	.b(FE_OFN272_n25595),
	.c(n23903));
   na02s01 U22584 (.o(n23887),
	.a(proc_input_NIB_storage_data_f_2__50_),
	.b(FE_OFN272_n25595));
   oa12f01 U22585 (.o(n3803),
	.a(n23886),
	.b(n17764),
	.c(n23908));
   na02s01 U22586 (.o(n23886),
	.a(proc_input_NIB_storage_data_f_2__49_),
	.b(n17764));
   oa12f01 U22587 (.o(n3808),
	.a(n23885),
	.b(n17764),
	.c(n23912));
   na02s01 U22588 (.o(n23885),
	.a(proc_input_NIB_storage_data_f_2__48_),
	.b(n17764));
   oa12f01 U22589 (.o(n3813),
	.a(n23884),
	.b(n17764),
	.c(n23914));
   na02s01 U22590 (.o(n23884),
	.a(proc_input_NIB_storage_data_f_2__47_),
	.b(n17764));
   oa12f01 U22591 (.o(n3818),
	.a(n23883),
	.b(n17764),
	.c(n23916));
   na02s01 U22592 (.o(n23883),
	.a(proc_input_NIB_storage_data_f_2__46_),
	.b(n17764));
   oa12f01 U22593 (.o(n3823),
	.a(n23882),
	.b(n17764),
	.c(n23942));
   na02s01 U22594 (.o(n23882),
	.a(proc_input_NIB_storage_data_f_2__45_),
	.b(n17764));
   oa12f01 U22595 (.o(n3828),
	.a(n23880),
	.b(n17764),
	.c(n23920));
   na02s01 U22596 (.o(n23880),
	.a(proc_input_NIB_storage_data_f_2__44_),
	.b(n17764));
   oa12f01 U22597 (.o(n3833),
	.a(n23774),
	.b(n17764),
	.c(n23806));
   oa12f01 U22598 (.o(n3838),
	.a(n23773),
	.b(n17764),
	.c(n23808));
   na02s01 U22599 (.o(n23773),
	.a(proc_input_NIB_storage_data_f_2__42_),
	.b(n17764));
   oa12f01 U22600 (.o(n3843),
	.a(n23871),
	.b(n17764),
	.c(n23928));
   na02s01 U22601 (.o(n23871),
	.a(proc_input_NIB_storage_data_f_2__41_),
	.b(n17764));
   oa12f01 U22602 (.o(n3848),
	.a(n23772),
	.b(n17764),
	.c(n23800));
   na02s01 U22603 (.o(n23772),
	.a(proc_input_NIB_storage_data_f_2__40_),
	.b(n17764));
   oa12f01 U22604 (.o(n3853),
	.a(n23869),
	.b(n17764),
	.c(n23934));
   na02s01 U22605 (.o(n23869),
	.a(proc_input_NIB_storage_data_f_2__39_),
	.b(n17764));
   oa12f01 U22606 (.o(n3858),
	.a(n23744),
	.b(n17764),
	.c(n23812));
   na02s01 U22607 (.o(n23744),
	.a(proc_input_NIB_storage_data_f_2__38_),
	.b(n17764));
   oa12f01 U22608 (.o(n3863),
	.a(n23745),
	.b(n17764),
	.c(n23796));
   na02s01 U22609 (.o(n23745),
	.a(proc_input_NIB_storage_data_f_2__37_),
	.b(n17764));
   oa12f01 U22610 (.o(n3868),
	.a(n23865),
	.b(n17764),
	.c(n23940));
   na02s01 U22611 (.o(n23865),
	.a(proc_input_NIB_storage_data_f_2__36_),
	.b(n17764));
   oa12f01 U22612 (.o(n3873),
	.a(n23864),
	.b(n17764),
	.c(n23944));
   na02s01 U22613 (.o(n23864),
	.a(proc_input_NIB_storage_data_f_2__35_),
	.b(n17764));
   oa12f01 U22614 (.o(n3878),
	.a(n23742),
	.b(n17764),
	.c(n23816));
   na02s01 U22615 (.o(n23742),
	.a(proc_input_NIB_storage_data_f_2__34_),
	.b(n17764));
   oa12f01 U22616 (.o(n3888),
	.a(n23862),
	.b(n17764),
	.c(n23905));
   na02s01 U22617 (.o(n23862),
	.a(proc_input_NIB_storage_data_f_2__32_),
	.b(n17764));
   oa12f01 U22618 (.o(n3893),
	.a(n23751),
	.b(n17764),
	.c(n23791));
   na02s01 U22619 (.o(n23751),
	.a(proc_input_NIB_storage_data_f_2__31_),
	.b(n17764));
   oa12f01 U22620 (.o(n3898),
	.a(n23857),
	.b(n17764),
	.c(n23894));
   na02s01 U22621 (.o(n23857),
	.a(proc_input_NIB_storage_data_f_2__30_),
	.b(n17764));
   oa12f01 U22622 (.o(n3903),
	.a(n23746),
	.b(n17764),
	.c(n23804));
   na02s01 U22623 (.o(n23746),
	.a(proc_input_NIB_storage_data_f_2__29_),
	.b(n17764));
   oa12f01 U22624 (.o(n3908),
	.a(n23758),
	.b(n17764),
	.c(n23814));
   oa12f01 U22625 (.o(n3913),
	.a(n23738),
	.b(n17764),
	.c(n23822));
   na02s01 U22626 (.o(n23738),
	.a(proc_input_NIB_storage_data_f_2__27_),
	.b(n17764));
   oa12f01 U22627 (.o(n3918),
	.a(n23756),
	.b(n17764),
	.c(n23818));
   na02s01 U22628 (.o(n23756),
	.a(proc_input_NIB_storage_data_f_2__26_),
	.b(n17764));
   oa12f01 U22629 (.o(n3923),
	.a(n23755),
	.b(n17764),
	.c(n23802));
   na02s01 U22630 (.o(n23755),
	.a(proc_input_NIB_storage_data_f_2__25_),
	.b(n17764));
   oa12f01 U22631 (.o(n3928),
	.a(n23754),
	.b(n17764),
	.c(n23798));
   na02s01 U22632 (.o(n23754),
	.a(proc_input_NIB_storage_data_f_2__24_),
	.b(n17764));
   oa12f01 U22633 (.o(n3933),
	.a(n23753),
	.b(n17764),
	.c(n23793));
   na02s01 U22634 (.o(n23753),
	.a(proc_input_NIB_storage_data_f_2__23_),
	.b(n17764));
   oa12f01 U22635 (.o(n3938),
	.a(n23759),
	.b(n17764),
	.c(n23820));
   na02s01 U22636 (.o(n23759),
	.a(proc_input_NIB_storage_data_f_2__22_),
	.b(n17764));
   oa22f01 U22637 (.o(n25585),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_2__10_),
	.d(n25595));
   oa22f01 U22638 (.o(n25586),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_2__9_),
	.d(n25595));
   oa22f01 U22639 (.o(n25587),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_2__8_),
	.d(n25595));
   oa22f01 U22640 (.o(n25588),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_2__7_),
	.d(n25595));
   oa22f01 U22641 (.o(n25589),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_2__6_),
	.d(n25595));
   oa22f01 U22642 (.o(n25590),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_2__5_),
	.d(n25595));
   oa22f01 U22643 (.o(n25591),
	.a(n17764),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_2__4_),
	.d(n25595));
   oa22f01 U22644 (.o(n25592),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_2__3_),
	.d(n25595));
   oa22f01 U22645 (.o(n25593),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_2__2_),
	.d(n25595));
   oa22f01 U22646 (.o(n25594),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_2__1_),
	.d(n25595));
   oa12s01 U22647 (.o(n4053),
	.a(n23824),
	.b(FE_OFN25775_FE_OFN582_n25619),
	.c(n23827));
   na02s01 U22648 (.o(n23824),
	.a(proc_input_NIB_storage_data_f_3__63_),
	.b(FE_OFN25775_FE_OFN582_n25619));
   oa12s01 U22649 (.o(n4058),
	.a(n23787),
	.b(FE_OFN25773_FE_OFN582_n25619),
	.c(n23810));
   na02s01 U22650 (.o(n23787),
	.a(proc_input_NIB_storage_data_f_3__62_),
	.b(FE_OFN25773_FE_OFN582_n25619));
   oa12s01 U22651 (.o(n4063),
	.a(n23844),
	.b(FE_OFN582_n25619),
	.c(n23918));
   na02s01 U22652 (.o(n23844),
	.a(proc_input_NIB_storage_data_f_3__61_),
	.b(FE_OFN582_n25619));
   oa12s01 U22653 (.o(n4068),
	.a(n23860),
	.b(FE_OFN25774_FE_OFN582_n25619),
	.c(n23926));
   na02s01 U22654 (.o(n23860),
	.a(proc_input_NIB_storage_data_f_3__60_),
	.b(FE_OFN25774_FE_OFN582_n25619));
   oa12s01 U22655 (.o(n4073),
	.a(n23842),
	.b(FE_OFN582_n25619),
	.c(n23938));
   na02s01 U22656 (.o(n23842),
	.a(proc_input_NIB_storage_data_f_3__59_),
	.b(FE_OFN582_n25619));
   oa12s01 U22657 (.o(n4078),
	.a(n23879),
	.b(FE_OFN25775_FE_OFN582_n25619),
	.c(n23936));
   na02s01 U22658 (.o(n23879),
	.a(proc_input_NIB_storage_data_f_3__58_),
	.b(FE_OFN25775_FE_OFN582_n25619));
   oa12s01 U22659 (.o(n4083),
	.a(n23840),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23932));
   na02f01 U22660 (.o(n23840),
	.a(proc_input_NIB_storage_data_f_3__57_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22661 (.o(n4088),
	.a(n23874),
	.b(FE_OFN25775_FE_OFN582_n25619),
	.c(n23930));
   na02s01 U22662 (.o(n23874),
	.a(proc_input_NIB_storage_data_f_3__56_),
	.b(FE_OFN25775_FE_OFN582_n25619));
   oa12s01 U22663 (.o(n4093),
	.a(n23873),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23910));
   na02s01 U22664 (.o(n23873),
	.a(proc_input_NIB_storage_data_f_3__55_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22665 (.o(n4098),
	.a(n23872),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23924));
   na02f01 U22666 (.o(n23872),
	.a(proc_input_NIB_storage_data_f_3__54_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22667 (.o(n4103),
	.a(n23833),
	.b(FE_OFN25775_FE_OFN582_n25619),
	.c(n23922));
   na02s01 U22668 (.o(n23833),
	.a(proc_input_NIB_storage_data_f_3__53_),
	.b(FE_OFN25775_FE_OFN582_n25619));
   oa12s01 U22669 (.o(n4108),
	.a(n23870),
	.b(FE_OFN25775_FE_OFN582_n25619),
	.c(n23890));
   na02s01 U22670 (.o(n23870),
	.a(proc_input_NIB_storage_data_f_3__52_),
	.b(FE_OFN25775_FE_OFN582_n25619));
   oa12s01 U22671 (.o(n4113),
	.a(n23838),
	.b(FE_OFN25774_FE_OFN582_n25619),
	.c(n23947));
   na02f02 U22672 (.o(n23838),
	.a(proc_input_NIB_storage_data_f_3__51_),
	.b(FE_OFN25774_FE_OFN582_n25619));
   oa12s01 U22673 (.o(n4118),
	.a(n23837),
	.b(FE_OFN25775_FE_OFN582_n25619),
	.c(n23903));
   na02s01 U22674 (.o(n23837),
	.a(proc_input_NIB_storage_data_f_3__50_),
	.b(FE_OFN25775_FE_OFN582_n25619));
   oa12f01 U22675 (.o(n4123),
	.a(n23867),
	.b(FE_OFN25778_FE_OFN582_n25619),
	.c(n23908));
   oa12s01 U22676 (.o(n4128),
	.a(n23866),
	.b(FE_OFN25778_FE_OFN582_n25619),
	.c(n23912));
   na02f01 U22677 (.o(n23866),
	.a(proc_input_NIB_storage_data_f_3__48_),
	.b(FE_OFN25778_FE_OFN582_n25619));
   oa12s01 U22678 (.o(n4133),
	.a(n23829),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23914));
   na02s01 U22679 (.o(n23829),
	.a(proc_input_NIB_storage_data_f_3__47_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22680 (.o(n4138),
	.a(n23843),
	.b(FE_OFN25778_FE_OFN582_n25619),
	.c(n23916));
   na02f01 U22681 (.o(n23843),
	.a(proc_input_NIB_storage_data_f_3__46_),
	.b(FE_OFN25778_FE_OFN582_n25619));
   oa12s01 U22682 (.o(n4143),
	.a(n23839),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23942));
   na02s01 U22683 (.o(n23839),
	.a(proc_input_NIB_storage_data_f_3__45_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22684 (.o(n4148),
	.a(n23841),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23920));
   na02s01 U22685 (.o(n23841),
	.a(proc_input_NIB_storage_data_f_3__44_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22686 (.o(n4153),
	.a(n23747),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23806));
   na02s01 U22687 (.o(n23747),
	.a(proc_input_NIB_storage_data_f_3__43_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22688 (.o(n4158),
	.a(n23741),
	.b(FE_OFN25778_FE_OFN582_n25619),
	.c(n23808));
   na02s01 U22689 (.o(n23741),
	.a(proc_input_NIB_storage_data_f_3__42_),
	.b(FE_OFN25778_FE_OFN582_n25619));
   oa12s01 U22690 (.o(n4163),
	.a(n23877),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23928));
   na02s01 U22691 (.o(n23877),
	.a(proc_input_NIB_storage_data_f_3__41_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22692 (.o(n4168),
	.a(n23740),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23800));
   na02s01 U22693 (.o(n23740),
	.a(proc_input_NIB_storage_data_f_3__40_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22694 (.o(n4173),
	.a(n23859),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23934));
   na02s01 U22695 (.o(n23859),
	.a(proc_input_NIB_storage_data_f_3__39_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22696 (.o(n4178),
	.a(n23743),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23812));
   na02s01 U22697 (.o(n23743),
	.a(proc_input_NIB_storage_data_f_3__38_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22698 (.o(n4183),
	.a(n23752),
	.b(FE_OFN25778_FE_OFN582_n25619),
	.c(n23796));
   na02f01 U22699 (.o(n23752),
	.a(proc_input_NIB_storage_data_f_3__37_),
	.b(FE_OFN25778_FE_OFN582_n25619));
   oa12s01 U22700 (.o(n4188),
	.a(n23858),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23940));
   na02s01 U22701 (.o(n23858),
	.a(proc_input_NIB_storage_data_f_3__36_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22702 (.o(n4193),
	.a(n23836),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23944));
   na02s01 U22703 (.o(n23836),
	.a(proc_input_NIB_storage_data_f_3__35_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22704 (.o(n4198),
	.a(n23748),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23816));
   oa12s01 U22705 (.o(n4208),
	.a(n23856),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23905));
   na02s01 U22706 (.o(n23856),
	.a(proc_input_NIB_storage_data_f_3__32_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22707 (.o(n4213),
	.a(n23749),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23791));
   na02s01 U22708 (.o(n23749),
	.a(proc_input_NIB_storage_data_f_3__31_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22709 (.o(n4218),
	.a(n23834),
	.b(FE_OFN25778_FE_OFN582_n25619),
	.c(n23894));
   na02f01 U22710 (.o(n23834),
	.a(proc_input_NIB_storage_data_f_3__30_),
	.b(FE_OFN25778_FE_OFN582_n25619));
   oa12s01 U22711 (.o(n4223),
	.a(n23750),
	.b(FE_OFN582_n25619),
	.c(n23804));
   na02s01 U22712 (.o(n23750),
	.a(proc_input_NIB_storage_data_f_3__29_),
	.b(FE_OFN582_n25619));
   oa12s01 U22713 (.o(n4228),
	.a(n23778),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23814));
   na02s01 U22714 (.o(n23778),
	.a(proc_input_NIB_storage_data_f_3__28_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22715 (.o(n4233),
	.a(n23779),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23822));
   na02s01 U22716 (.o(n23779),
	.a(proc_input_NIB_storage_data_f_3__27_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22717 (.o(n4238),
	.a(n23780),
	.b(FE_OFN25778_FE_OFN582_n25619),
	.c(n23818));
   na02s01 U22718 (.o(n23780),
	.a(proc_input_NIB_storage_data_f_3__26_),
	.b(FE_OFN25778_FE_OFN582_n25619));
   oa12s01 U22719 (.o(n4243),
	.a(n23781),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23802));
   na02s01 U22720 (.o(n23781),
	.a(proc_input_NIB_storage_data_f_3__25_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa12s01 U22721 (.o(n4248),
	.a(n23782),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23798));
   na02s01 U22722 (.o(n23782),
	.a(proc_input_NIB_storage_data_f_3__24_),
	.b(FE_OFN582_n25619));
   oa12s01 U22723 (.o(n4253),
	.a(n23783),
	.b(FE_OFN25778_FE_OFN582_n25619),
	.c(n23793));
   na02f01 U22724 (.o(n23783),
	.a(proc_input_NIB_storage_data_f_3__23_),
	.b(FE_OFN25778_FE_OFN582_n25619));
   oa12s01 U22725 (.o(n4258),
	.a(n23757),
	.b(FE_OFN25777_FE_OFN582_n25619),
	.c(n23820));
   na02s01 U22726 (.o(n23757),
	.a(proc_input_NIB_storage_data_f_3__22_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa22s01 U22727 (.o(n25609),
	.a(FE_OFN25776_FE_OFN582_n25619),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_3__10_),
	.d(n25619));
   oa22s01 U22728 (.o(n25610),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_3__9_),
	.d(n25619));
   oa22s01 U22729 (.o(n25611),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_3__8_),
	.d(n25619));
   oa22s01 U22730 (.o(n25612),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_3__7_),
	.d(n25619));
   oa22s01 U22731 (.o(n25614),
	.a(FE_OFN25776_FE_OFN582_n25619),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_3__5_),
	.d(n25619));
   oa22s01 U22732 (.o(n25615),
	.a(FE_OFN25777_FE_OFN582_n25619),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_3__4_),
	.d(n17763));
   oa22s01 U22733 (.o(n25616),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_3__3_),
	.d(n25619));
   oa22s01 U22734 (.o(n25617),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_3__2_),
	.d(n25619));
   oa22s01 U22735 (.o(n25618),
	.a(FE_OFN25777_FE_OFN582_n25619),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_3__1_),
	.d(n17763));
   oa22s01 U22736 (.o(n25620),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_3__0_),
	.d(n25619));
   oa12m01 U22737 (.o(n4373),
	.a(n23654),
	.b(n23827),
	.c(FE_OFN25763_FE_OFN1077_n17766));
   oa12m01 U22738 (.o(n4378),
	.a(n23655),
	.b(n23810),
	.c(FE_OFN25763_FE_OFN1077_n17766));
   oa12m01 U22739 (.o(n4383),
	.a(n23656),
	.b(FE_OFN25763_FE_OFN1077_n17766),
	.c(n23918));
   oa12m01 U22740 (.o(n4388),
	.a(n23659),
	.b(n23926),
	.c(FE_OFN25763_FE_OFN1077_n17766));
   oa12m01 U22741 (.o(n4393),
	.a(n23660),
	.b(n23938),
	.c(FE_OFN25763_FE_OFN1077_n17766));
   oa12m01 U22742 (.o(n4398),
	.a(n23726),
	.b(FE_OFN25763_FE_OFN1077_n17766),
	.c(n23936));
   oa12m01 U22743 (.o(n4403),
	.a(n23595),
	.b(n23932),
	.c(FE_OFN25763_FE_OFN1077_n17766));
   oa12m01 U22744 (.o(n4408),
	.a(n23662),
	.b(FE_OFN25763_FE_OFN1077_n17766),
	.c(n23930));
   oa12m01 U22745 (.o(n4413),
	.a(n23723),
	.b(n23910),
	.c(FE_OFN25763_FE_OFN1077_n17766));
   oa12m01 U22746 (.o(n4418),
	.a(n23663),
	.b(n23924),
	.c(FE_OFN25765_FE_OFN1077_n17766));
   oa12m01 U22747 (.o(n4423),
	.a(n23724),
	.b(FE_OFN25763_FE_OFN1077_n17766),
	.c(n23922));
   oa12m01 U22748 (.o(n4428),
	.a(n23666),
	.b(FE_OFN25763_FE_OFN1077_n17766),
	.c(n23890));
   oa12m01 U22749 (.o(n4433),
	.a(n23725),
	.b(n23947),
	.c(FE_OFN25763_FE_OFN1077_n17766));
   oa12m01 U22750 (.o(n4438),
	.a(n23597),
	.b(FE_OFN25763_FE_OFN1077_n17766),
	.c(n23903));
   oa12m01 U22751 (.o(n4443),
	.a(n23602),
	.b(FE_OFN25768_FE_OFN1077_n17766),
	.c(n23908));
   oa12m01 U22752 (.o(n4448),
	.a(n23677),
	.b(FE_OFN25768_FE_OFN1077_n17766),
	.c(n23912));
   oa12m01 U22753 (.o(n4453),
	.a(n23166),
	.b(n23914),
	.c(n17766));
   oa12m01 U22754 (.o(n4458),
	.a(n23670),
	.b(FE_OFN25768_FE_OFN1077_n17766),
	.c(n23916));
   oa12m01 U22755 (.o(n4463),
	.a(n23180),
	.b(n17766),
	.c(n23942));
   oa12m01 U22756 (.o(n4468),
	.a(n23177),
	.b(n17766),
	.c(n23920));
   oa12m01 U22757 (.o(n4473),
	.a(n23172),
	.b(n23806),
	.c(FE_OFN1074_n17766));
   oa12m01 U22758 (.o(n4478),
	.a(n23161),
	.b(n23808),
	.c(FE_OFN25768_FE_OFN1077_n17766));
   oa12m01 U22759 (.o(n4483),
	.a(n23165),
	.b(n17766),
	.c(n23928));
   oa12m01 U22760 (.o(n4488),
	.a(n23176),
	.b(n17766),
	.c(n23800));
   oa12m01 U22761 (.o(n4493),
	.a(n23715),
	.b(n17766),
	.c(n23934));
   oa12m01 U22762 (.o(n4498),
	.a(n23355),
	.b(FE_OFN25768_FE_OFN1077_n17766),
	.c(n23812));
   oa12m01 U22763 (.o(n4503),
	.a(n23159),
	.b(FE_OFN25768_FE_OFN1077_n17766),
	.c(n23796));
   oa12m01 U22764 (.o(n4508),
	.a(n23352),
	.b(n23940),
	.c(FE_OFN25768_FE_OFN1077_n17766));
   oa12m01 U22765 (.o(n4513),
	.a(n23351),
	.b(FE_OFN25768_FE_OFN1077_n17766),
	.c(n23944));
   oa12m01 U22766 (.o(n4518),
	.a(n23359),
	.b(n23816),
	.c(FE_OFN25768_FE_OFN1077_n17766));
   oa12m01 U22767 (.o(n4528),
	.a(n23596),
	.b(FE_OFN25768_FE_OFN1077_n17766),
	.c(n23905));
   oa12m01 U22768 (.o(n4533),
	.a(n23357),
	.b(FE_OFN25765_FE_OFN1077_n17766),
	.c(n23791));
   oa12m01 U22769 (.o(n4538),
	.a(n23354),
	.b(n23894),
	.c(FE_OFN25768_FE_OFN1077_n17766));
   oa12m01 U22770 (.o(n4543),
	.a(n23669),
	.b(FE_OFN1076_n17766),
	.c(n23804));
   oa12m01 U22771 (.o(n4548),
	.a(n23651),
	.b(FE_OFN1075_n17766),
	.c(n23814));
   oa12m01 U22772 (.o(n4553),
	.a(n23641),
	.b(n17766),
	.c(n23822));
   oa12m01 U22773 (.o(n4558),
	.a(n23638),
	.b(n17766),
	.c(n23818));
   oa12m01 U22774 (.o(n4563),
	.a(n23639),
	.b(FE_OFN25768_FE_OFN1077_n17766),
	.c(n23802));
   oa12m01 U22775 (.o(n4568),
	.a(n23644),
	.b(n23798),
	.c(n17766));
   oa12m01 U22776 (.o(n4573),
	.a(n23657),
	.b(n17766),
	.c(n23793));
   oa12m01 U22777 (.o(n4578),
	.a(n23642),
	.b(FE_OFN1075_n17766),
	.c(n23820));
   oa22m01 U22778 (.o(n23121),
	.a(FE_OFN25761_FE_OFN1077_n17766),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_4__14_),
	.d(n23090));
   oa22m01 U22779 (.o(n23145),
	.a(FE_OFN25760_FE_OFN1077_n17766),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_4__2_),
	.d(n23090));
   oa22m01 U22780 (.o(n23144),
	.a(FE_OFN1077_n17766),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_4__1_),
	.d(n23090));
   oa22m01 U22781 (.o(n23135),
	.a(FE_OFN25760_FE_OFN1077_n17766),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_4__0_),
	.d(n23090));
   oa12f01 U22782 (.o(n4693),
	.a(n23647),
	.b(n23827),
	.c(FE_OFN368_n17761));
   oa12f01 U22783 (.o(n4698),
	.a(n23648),
	.b(n23810),
	.c(FE_OFN368_n17761));
   oa12s01 U22784 (.o(n4703),
	.a(n23649),
	.b(n23918),
	.c(FE_OFN368_n17761));
   oa12f01 U22785 (.o(n4708),
	.a(n23645),
	.b(n23926),
	.c(FE_OFN368_n17761));
   oa12s01 U22786 (.o(n4713),
	.a(n23643),
	.b(n23938),
	.c(FE_OFN368_n17761));
   oa12s01 U22787 (.o(n4718),
	.a(n23713),
	.b(n23936),
	.c(FE_OFN368_n17761));
   oa12f01 U22788 (.o(n4723),
	.a(n23608),
	.b(n23932),
	.c(FE_OFN368_n17761));
   oa12f01 U22789 (.o(n4728),
	.a(n23665),
	.b(n23930),
	.c(FE_OFN368_n17761));
   oa12f01 U22790 (.o(n4733),
	.a(n23714),
	.b(n23910),
	.c(FE_OFN368_n17761));
   oa12f01 U22791 (.o(n4738),
	.a(n23646),
	.b(n23924),
	.c(FE_OFN368_n17761));
   oa12f01 U22792 (.o(n4743),
	.a(n23721),
	.b(n23922),
	.c(FE_OFN368_n17761));
   oa12f01 U22793 (.o(n4748),
	.a(n23650),
	.b(n23890),
	.c(FE_OFN368_n17761));
   oa12f01 U22794 (.o(n4753),
	.a(n23719),
	.b(n23947),
	.c(FE_OFN368_n17761));
   oa12f01 U22795 (.o(n4758),
	.a(n23606),
	.b(n23903),
	.c(FE_OFN368_n17761));
   oa12s01 U22796 (.o(n4763),
	.a(n23607),
	.b(n23908),
	.c(FE_OFN369_n17761));
   oa12s01 U22797 (.o(n4768),
	.a(n23652),
	.b(n23912),
	.c(FE_OFN369_n17761));
   oa12f01 U22798 (.o(n4773),
	.a(n23167),
	.b(n23914),
	.c(FE_OFN369_n17761));
   oa12s01 U22799 (.o(n4778),
	.a(n23653),
	.b(n23916),
	.c(FE_OFN369_n17761));
   oa12f01 U22800 (.o(n4783),
	.a(n23178),
	.b(n23942),
	.c(FE_OFN368_n17761));
   oa12f01 U22801 (.o(n4788),
	.a(n23160),
	.b(n23920),
	.c(FE_OFN368_n17761));
   oa12f01 U22802 (.o(n4793),
	.a(n23168),
	.b(n23806),
	.c(FE_OFN369_n17761));
   oa12s01 U22803 (.o(n4798),
	.a(n23173),
	.b(n23808),
	.c(FE_OFN369_n17761));
   oa12f01 U22804 (.o(n4803),
	.a(n23156),
	.b(n23928),
	.c(FE_OFN369_n17761));
   oa12f01 U22805 (.o(n4808),
	.a(n23171),
	.b(n23800),
	.c(FE_OFN368_n17761));
   oa12f01 U22806 (.o(n4813),
	.a(n23353),
	.b(n23934),
	.c(FE_OFN368_n17761));
   oa12f01 U22807 (.o(n4818),
	.a(n23356),
	.b(n23812),
	.c(FE_OFN369_n17761));
   oa12s01 U22808 (.o(n4823),
	.a(n23182),
	.b(n23796),
	.c(FE_OFN369_n17761));
   oa12f01 U22809 (.o(n4828),
	.a(n23727),
	.b(n23940),
	.c(FE_OFN368_n17761));
   oa12f01 U22810 (.o(n4833),
	.a(n23363),
	.b(n23944),
	.c(FE_OFN369_n17761));
   oa12s01 U22811 (.o(n4838),
	.a(n23364),
	.b(n23816),
	.c(FE_OFN369_n17761));
   oa12f01 U22812 (.o(n4848),
	.a(n23609),
	.b(FE_OFN369_n17761),
	.c(n23905));
   oa12f01 U22813 (.o(n4853),
	.a(n23366),
	.b(n23791),
	.c(FE_OFN368_n17761));
   oa12s01 U22814 (.o(n4858),
	.a(n23367),
	.b(n23894),
	.c(FE_OFN369_n17761));
   oa12s01 U22815 (.o(n4863),
	.a(n23658),
	.b(n23804),
	.c(n17761));
   oa12f01 U22816 (.o(n4868),
	.a(n23661),
	.b(n23814),
	.c(FE_OFN368_n17761));
   oa12f01 U22817 (.o(n4873),
	.a(n23664),
	.b(n23822),
	.c(FE_OFN368_n17761));
   oa12s01 U22818 (.o(n4878),
	.a(n23667),
	.b(n23818),
	.c(FE_OFN113_n23102));
   oa12s01 U22819 (.o(n4883),
	.a(n23668),
	.b(n23802),
	.c(FE_OFN369_n17761));
   oa12s01 U22820 (.o(n4888),
	.a(n23672),
	.b(n23798),
	.c(FE_OFN114_n23102));
   oa12s01 U22821 (.o(n4893),
	.a(n23680),
	.b(n23793),
	.c(FE_OFN369_n17761));
   oa12s01 U22822 (.o(n4898),
	.a(n23683),
	.b(n23820),
	.c(FE_OFN370_n17761));
   oa22m01 U22823 (.o(n23132),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_5__21_),
	.d(n23102));
   oa22m01 U22824 (.o(n23130),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_5__19_),
	.d(n23102));
   oa22m01 U22825 (.o(n23127),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_5__18_),
	.d(n23102));
   oa22m01 U22826 (.o(n23126),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_5__17_),
	.d(n23102));
   oa22m01 U22827 (.o(n23125),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_5__16_),
	.d(n23102));
   oa22m01 U22828 (.o(n23124),
	.a(FE_OFN369_n17761),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_5__15_),
	.d(n23102));
   oa22m01 U22829 (.o(n23122),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_5__14_),
	.d(n23102));
   oa22m01 U22830 (.o(n23120),
	.a(FE_OFN369_n17761),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_5__13_),
	.d(n23102));
   oa22m01 U22831 (.o(n23118),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_5__12_),
	.d(n23102));
   oa22m01 U22832 (.o(n23117),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_5__11_),
	.d(n23102));
   oa22m01 U22833 (.o(n23115),
	.a(FE_OFN369_n17761),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_5__10_),
	.d(n23102));
   oa22m01 U22834 (.o(n23113),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_5__9_),
	.d(n23102));
   oa22m01 U22835 (.o(n23112),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_5__8_),
	.d(n23102));
   oa22m01 U22836 (.o(n23111),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_5__7_),
	.d(n23102));
   oa22m01 U22837 (.o(n23110),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_5__6_),
	.d(n23102));
   oa22m01 U22838 (.o(n23108),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_5__4_),
	.d(n23102));
   oa22m01 U22839 (.o(n23107),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_5__3_),
	.d(n23102));
   oa22m01 U22840 (.o(n23106),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_5__2_),
	.d(n23102));
   oa22m01 U22841 (.o(n23105),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_5__1_),
	.d(n23102));
   oa22m01 U22842 (.o(n23103),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_5__0_),
	.d(n23102));
   oa12f01 U22843 (.o(n5013),
	.a(n23686),
	.b(n23827),
	.c(FE_OFN442_n23051));
   na02s01 U22844 (.o(n23686),
	.a(proc_input_NIB_storage_data_f_6__63_),
	.b(FE_OFN442_n23051));
   oa12f01 U22845 (.o(n5018),
	.a(n23692),
	.b(n23810),
	.c(FE_OFN442_n23051));
   na02s01 U22846 (.o(n23692),
	.a(proc_input_NIB_storage_data_f_6__62_),
	.b(FE_OFN442_n23051));
   oa12s01 U22847 (.o(n5023),
	.a(n23694),
	.b(n23918),
	.c(FE_OFN442_n23051));
   na02s01 U22848 (.o(n23694),
	.a(proc_input_NIB_storage_data_f_6__61_),
	.b(FE_OFN442_n23051));
   oa12f01 U22849 (.o(n5028),
	.a(n23682),
	.b(n23926),
	.c(FE_OFN442_n23051));
   na02s01 U22850 (.o(n23682),
	.a(proc_input_NIB_storage_data_f_6__60_),
	.b(FE_OFN442_n23051));
   oa12s01 U22851 (.o(n5033),
	.a(n23720),
	.b(n23938),
	.c(FE_OFN442_n23051));
   oa12s01 U22852 (.o(n5038),
	.a(n23698),
	.b(n23936),
	.c(FE_OFN442_n23051));
   na02s01 U22853 (.o(n23698),
	.a(proc_input_NIB_storage_data_f_6__58_),
	.b(FE_OFN442_n23051));
   oa12f01 U22854 (.o(n5043),
	.a(n23610),
	.b(n23932),
	.c(FE_OFN442_n23051));
   oa12f01 U22855 (.o(n5048),
	.a(n23688),
	.b(n23930),
	.c(FE_OFN442_n23051));
   na02s01 U22856 (.o(n23688),
	.a(proc_input_NIB_storage_data_f_6__56_),
	.b(FE_OFN442_n23051));
   oa12f01 U22857 (.o(n5053),
	.a(n23640),
	.b(n23910),
	.c(FE_OFN442_n23051));
   na02f01 U22858 (.o(n23640),
	.a(proc_input_NIB_storage_data_f_6__55_),
	.b(FE_OFN442_n23051));
   oa12f01 U22859 (.o(n5058),
	.a(n23722),
	.b(n23924),
	.c(FE_OFN442_n23051));
   oa12f01 U22860 (.o(n5063),
	.a(n23684),
	.b(n23922),
	.c(FE_OFN442_n23051));
   na02f01 U22861 (.o(n23684),
	.a(proc_input_NIB_storage_data_f_6__53_),
	.b(FE_OFN442_n23051));
   oa12f01 U22862 (.o(n5068),
	.a(n23718),
	.b(n23890),
	.c(FE_OFN442_n23051));
   oa12f01 U22863 (.o(n5073),
	.a(n23605),
	.b(n23947),
	.c(FE_OFN442_n23051));
   oa12f01 U22864 (.o(n5078),
	.a(n23604),
	.b(n23903),
	.c(FE_OFN442_n23051));
   oa12f01 U22865 (.o(n5083),
	.a(n23691),
	.b(n23908),
	.c(FE_OFN25806_n23051));
   na02f01 U22866 (.o(n23691),
	.a(proc_input_NIB_storage_data_f_6__49_),
	.b(FE_OFN25806_n23051));
   oa12f01 U22867 (.o(n5088),
	.a(n23693),
	.b(n23912),
	.c(FE_OFN25806_n23051));
   na02f01 U22868 (.o(n23693),
	.a(proc_input_NIB_storage_data_f_6__48_),
	.b(FE_OFN25806_n23051));
   oa12f01 U22869 (.o(n5093),
	.a(n23365),
	.b(n23914),
	.c(FE_OFN25801_n23051));
   oa12f01 U22870 (.o(n5098),
	.a(n23716),
	.b(n23916),
	.c(FE_OFN25806_n23051));
   oa12f01 U22871 (.o(n5103),
	.a(n23361),
	.b(n23942),
	.c(FE_OFN25798_n23051));
   oa12f01 U22872 (.o(n5108),
	.a(n23368),
	.b(n23920),
	.c(FE_OFN25798_n23051));
   oa12f01 U22873 (.o(n5113),
	.a(n23370),
	.b(n23806),
	.c(FE_OFN25801_n23051));
   oa12f01 U22874 (.o(n5118),
	.a(n23358),
	.b(n23808),
	.c(FE_OFN25798_n23051));
   oa12f01 U22875 (.o(n5123),
	.a(n23369),
	.b(n23928),
	.c(FE_OFN25802_n23051));
   oa12f01 U22876 (.o(n5128),
	.a(n23362),
	.b(n23800),
	.c(FE_OFN25798_n23051));
   oa12f01 U22877 (.o(n5133),
	.a(n23179),
	.b(n23934),
	.c(FE_OFN25801_n23051));
   oa12f01 U22878 (.o(n5138),
	.a(n23155),
	.b(n23812),
	.c(FE_OFN25801_n23051));
   oa12f01 U22879 (.o(n5143),
	.a(n23360),
	.b(n23796),
	.c(FE_OFN25802_n23051));
   oa12f01 U22880 (.o(n5148),
	.a(n23717),
	.b(n23940),
	.c(FE_OFN25801_n23051));
   oa12f01 U22881 (.o(n5153),
	.a(n23174),
	.b(n23944),
	.c(FE_OFN25801_n23051));
   oa12f01 U22882 (.o(n5158),
	.a(n23175),
	.b(n23816),
	.c(FE_OFN25801_n23051));
   oa22f01 U22883 (.o(n23096),
	.a(FE_OFN25798_n23051),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_6__33_),
	.d(FE_OFN440_n23051));
   oa12f01 U22884 (.o(n5168),
	.a(n23603),
	.b(FE_OFN25802_n23051),
	.c(n23905));
   oa12f01 U22885 (.o(n5173),
	.a(n23181),
	.b(n23791),
	.c(FE_OFN25798_n23051));
   oa12f01 U22886 (.o(n5178),
	.a(n23170),
	.b(n23894),
	.c(FE_OFN25806_n23051));
   oa12f01 U22887 (.o(n5183),
	.a(n23701),
	.b(n23804),
	.c(FE_OFN25798_n23051));
   na02f01 U22888 (.o(n23701),
	.a(proc_input_NIB_storage_data_f_6__29_),
	.b(FE_OFN25798_n23051));
   oa12f01 U22889 (.o(n5188),
	.a(n23704),
	.b(n23814),
	.c(FE_OFN25801_n23051));
   na02s01 U22890 (.o(n23704),
	.a(proc_input_NIB_storage_data_f_6__28_),
	.b(FE_OFN25801_n23051));
   oa12f01 U22891 (.o(n5193),
	.a(n23685),
	.b(n23822),
	.c(FE_OFN25801_n23051));
   na02s01 U22892 (.o(n23685),
	.a(proc_input_NIB_storage_data_f_6__27_),
	.b(FE_OFN25801_n23051));
   oa12f01 U22893 (.o(n5198),
	.a(n23702),
	.b(n23818),
	.c(FE_OFN25806_n23051));
   na02f01 U22894 (.o(n23702),
	.a(proc_input_NIB_storage_data_f_6__26_),
	.b(FE_OFN25806_n23051));
   oa12f01 U22895 (.o(n5203),
	.a(n23707),
	.b(n23802),
	.c(FE_OFN25801_n23051));
   oa12f01 U22896 (.o(n5208),
	.a(n23705),
	.b(n23798),
	.c(FE_OFN25798_n23051));
   na02f01 U22897 (.o(n23705),
	.a(proc_input_NIB_storage_data_f_6__24_),
	.b(FE_OFN25798_n23051));
   oa12f01 U22898 (.o(n5213),
	.a(n23706),
	.b(n23793),
	.c(FE_OFN25802_n23051));
   na02f01 U22899 (.o(n23706),
	.a(proc_input_NIB_storage_data_f_6__23_),
	.b(FE_OFN25802_n23051));
   oa12f01 U22900 (.o(n5218),
	.a(n23696),
	.b(n23820),
	.c(FE_OFN25801_n23051));
   na02s01 U22901 (.o(n23696),
	.a(proc_input_NIB_storage_data_f_6__22_),
	.b(FE_OFN25801_n23051));
   oa22s01 U22902 (.o(n23095),
	.a(n23051),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_6__21_),
	.d(FE_OFN440_n23051));
   oa22f01 U22903 (.o(n23094),
	.a(FE_OFN25798_n23051),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_6__20_),
	.d(FE_OFN440_n23051));
   oa22s01 U22904 (.o(n23093),
	.a(n23051),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_6__19_),
	.d(FE_OFN440_n23051));
   oa22f01 U22905 (.o(n23092),
	.a(n23051),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_6__18_),
	.d(FE_OFN440_n23051));
   oa22s01 U22906 (.o(n23088),
	.a(n23051),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_6__17_),
	.d(FE_OFN440_n23051));
   oa22s01 U22907 (.o(n23075),
	.a(n23051),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_6__16_),
	.d(FE_OFN440_n23051));
   oa22f01 U22908 (.o(n23086),
	.a(FE_OFN25798_n23051),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_6__15_),
	.d(FE_OFN440_n23051));
   oa22f01 U22909 (.o(n23084),
	.a(FE_OFN25798_n23051),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_6__14_),
	.d(FE_OFN440_n23051));
   oa22f01 U22910 (.o(n23081),
	.a(FE_OFN25798_n23051),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_6__13_),
	.d(FE_OFN440_n23051));
   oa22f01 U22911 (.o(n23073),
	.a(n23051),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_6__11_),
	.d(FE_OFN440_n23051));
   oa22f01 U22912 (.o(n23072),
	.a(FE_OFN25798_n23051),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_6__10_),
	.d(FE_OFN440_n23051));
   oa22s01 U22913 (.o(n23071),
	.a(n23051),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_6__9_),
	.d(FE_OFN440_n23051));
   oa22s01 U22914 (.o(n23060),
	.a(n23051),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_6__8_),
	.d(FE_OFN440_n23051));
   oa22s01 U22915 (.o(n23068),
	.a(n23051),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_6__7_),
	.d(FE_OFN440_n23051));
   oa22s01 U22916 (.o(n23087),
	.a(n23051),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_6__6_),
	.d(FE_OFN440_n23051));
   oa22f01 U22917 (.o(n23057),
	.a(FE_OFN25798_n23051),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_6__5_),
	.d(FE_OFN440_n23051));
   oa22f01 U22918 (.o(n23085),
	.a(FE_OFN25798_n23051),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_6__4_),
	.d(FE_OFN440_n23051));
   oa22s01 U22919 (.o(n23063),
	.a(n23051),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_6__3_),
	.d(FE_OFN440_n23051));
   oa22s01 U22920 (.o(n23082),
	.a(n23051),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_6__2_),
	.d(FE_OFN440_n23051));
   oa22s01 U22921 (.o(n23052),
	.a(n23051),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_6__1_),
	.d(FE_OFN440_n23051));
   oa22f01 U22922 (.o(n23076),
	.a(FE_OFN25798_n23051),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_6__0_),
	.d(FE_OFN440_n23051));
   oa12s01 U22923 (.o(n5333),
	.a(n23687),
	.b(FE_OFN1081_n17767),
	.c(n23827));
   oa12s01 U22924 (.o(n5338),
	.a(n23708),
	.b(n17767),
	.c(n23810));
   oa12s01 U22925 (.o(n5343),
	.a(n23709),
	.b(n23918),
	.c(n17767));
   oa12f01 U22926 (.o(n5348),
	.a(n23695),
	.b(n17767),
	.c(n23926));
   oa12s01 U22927 (.o(n5353),
	.a(n23730),
	.b(FE_OFN1081_n17767),
	.c(n23938));
   oa12s01 U22928 (.o(n5358),
	.a(n23703),
	.b(n23936),
	.c(n17767));
   oa12s01 U22929 (.o(n5363),
	.a(n23601),
	.b(FE_OFN1081_n17767),
	.c(n23932));
   oa12s01 U22930 (.o(n5368),
	.a(n23700),
	.b(n23930),
	.c(FE_OFN1081_n17767));
   oa12s01 U22931 (.o(n5373),
	.a(n23699),
	.b(FE_OFN1081_n17767),
	.c(n23910));
   oa12s01 U22932 (.o(n5378),
	.a(n23731),
	.b(FE_OFN1081_n17767),
	.c(n23924));
   oa12s01 U22933 (.o(n5383),
	.a(n23697),
	.b(n23922),
	.c(FE_OFN1081_n17767));
   oa12s01 U22934 (.o(n5388),
	.a(n23729),
	.b(n23890),
	.c(FE_OFN1081_n17767));
   oa12s01 U22935 (.o(n5393),
	.a(n23599),
	.b(n17767),
	.c(n23947));
   oa12s01 U22936 (.o(n5398),
	.a(n23598),
	.b(n23903),
	.c(FE_OFN1081_n17767));
   oa12s01 U22937 (.o(n5403),
	.a(n23690),
	.b(n23908),
	.c(n17767));
   oa12s01 U22938 (.o(n5408),
	.a(n23689),
	.b(n23912),
	.c(n17767));
   oa12s01 U22939 (.o(n5413),
	.a(n23371),
	.b(n17767),
	.c(n23914));
   oa12s01 U22940 (.o(n5418),
	.a(n23728),
	.b(n23916),
	.c(n17767));
   oa12s01 U22941 (.o(n5423),
	.a(n23373),
	.b(n23942),
	.c(FE_OFN1081_n17767));
   oa12s01 U22942 (.o(n5428),
	.a(n23375),
	.b(n23920),
	.c(FE_OFN1081_n17767));
   oa12s01 U22943 (.o(n5433),
	.a(n23376),
	.b(n17767),
	.c(n23806));
   oa12s01 U22944 (.o(n5438),
	.a(n23377),
	.b(n17767),
	.c(n23808));
   oa12f01 U22945 (.o(n5443),
	.a(n23374),
	.b(n23928),
	.c(n17767));
   oa12s01 U22946 (.o(n5448),
	.a(n23378),
	.b(n23800),
	.c(FE_OFN1081_n17767));
   oa12s01 U22947 (.o(n5453),
	.a(n23169),
	.b(n23934),
	.c(FE_OFN1081_n17767));
   oa12s01 U22948 (.o(n5458),
	.a(n23157),
	.b(n23812),
	.c(n17767));
   oa12s01 U22949 (.o(n5463),
	.a(n23372),
	.b(n23796),
	.c(n17767));
   oa12s01 U22950 (.o(n5468),
	.a(n23732),
	.b(FE_OFN907_n23046),
	.c(n23940));
   oa12s01 U22951 (.o(n5473),
	.a(n23158),
	.b(n23944),
	.c(n17767));
   oa12s01 U22952 (.o(n5478),
	.a(n23162),
	.b(n17767),
	.c(n23816));
   oa22s01 U22953 (.o(n23142),
	.a(n17767),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_7__33_),
	.d(n23046));
   oa12s01 U22954 (.o(n5488),
	.a(n23600),
	.b(n17767),
	.c(n23905));
   oa12s01 U22955 (.o(n5493),
	.a(n23163),
	.b(n23791),
	.c(FE_OFN1081_n17767));
   oa12s01 U22956 (.o(n5498),
	.a(n23164),
	.b(n17767),
	.c(n23894));
   oa12s01 U22957 (.o(n5503),
	.a(n23681),
	.b(n23804),
	.c(FE_OFN1080_n17767));
   oa12s01 U22958 (.o(n5508),
	.a(n23679),
	.b(n23814),
	.c(FE_OFN907_n23046));
   oa12s01 U22959 (.o(n5513),
	.a(n23678),
	.b(n23822),
	.c(FE_OFN907_n23046));
   oa12s01 U22960 (.o(n5518),
	.a(n23676),
	.b(n23818),
	.c(n17767));
   oa12s01 U22961 (.o(n5523),
	.a(n23675),
	.b(n23802),
	.c(n17767));
   oa12s01 U22962 (.o(n5528),
	.a(n23674),
	.b(n17767),
	.c(n23798));
   oa12s01 U22963 (.o(n5533),
	.a(n23673),
	.b(n23793),
	.c(n17767));
   oa12s01 U22964 (.o(n5538),
	.a(n23671),
	.b(n23820),
	.c(n17767));
   oa22s01 U22965 (.o(n23083),
	.a(FE_OFN1081_n17767),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_7__21_),
	.d(n23046));
   oa22s01 U22966 (.o(n23077),
	.a(FE_OFN1081_n17767),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_7__20_),
	.d(n23046));
   oa22s01 U22967 (.o(n23074),
	.a(n17767),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_7__19_),
	.d(n23046));
   oa22s01 U22968 (.o(n23070),
	.a(n17767),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_7__17_),
	.d(n23046));
   oa22s01 U22969 (.o(n23069),
	.a(FE_OFN1081_n17767),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_7__16_),
	.d(n23046));
   oa22s01 U22970 (.o(n23067),
	.a(n17767),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_7__15_),
	.d(n23046));
   oa22s01 U22971 (.o(n23066),
	.a(n17767),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_7__14_),
	.d(n23046));
   oa22s01 U22972 (.o(n23053),
	.a(n17767),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_7__13_),
	.d(n23046));
   oa22s01 U22973 (.o(n23059),
	.a(FE_OFN1081_n17767),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_7__12_),
	.d(n23046));
   oa22s01 U22974 (.o(n23056),
	.a(FE_OFN1081_n17767),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_7__11_),
	.d(n23046));
   oa22s01 U22975 (.o(n23048),
	.a(n17767),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_7__10_),
	.d(n23046));
   oa22s01 U22976 (.o(n23058),
	.a(n17767),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_7__9_),
	.d(n23046));
   oa22s01 U22977 (.o(n23055),
	.a(n17767),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_7__8_),
	.d(n23046));
   oa22s01 U22978 (.o(n23047),
	.a(n17767),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_7__7_),
	.d(n23046));
   oa22s01 U22979 (.o(n23054),
	.a(n17767),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_7__6_),
	.d(n23046));
   oa22s01 U22980 (.o(n23049),
	.a(n17767),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_7__5_),
	.d(n23046));
   oa22s01 U22981 (.o(n23061),
	.a(n17767),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_7__4_),
	.d(n23046));
   oa22s01 U22982 (.o(n23078),
	.a(n17767),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_7__2_),
	.d(n23046));
   oa22s01 U22983 (.o(n23064),
	.a(FE_OFN1081_n17767),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_7__1_),
	.d(n23046));
   oa22s01 U22984 (.o(n23080),
	.a(n17767),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_7__0_),
	.d(n23046));
   oa12s01 U22985 (.o(n6613),
	.a(n23392),
	.b(FE_OFN1085_n22923),
	.c(n23827));
   na02s01 U22986 (.o(n23392),
	.a(proc_input_NIB_storage_data_f_11__63_),
	.b(FE_OFN1085_n22923));
   oa12s01 U22987 (.o(n6618),
	.a(n23394),
	.b(FE_OFN1085_n22923),
	.c(n23810));
   oa12s01 U22988 (.o(n6623),
	.a(n23393),
	.b(FE_OFN1085_n22923),
	.c(n23918));
   oa12s01 U22989 (.o(n6628),
	.a(n23389),
	.b(FE_OFN1085_n22923),
	.c(n23926));
   na02s01 U22990 (.o(n23389),
	.a(proc_input_NIB_storage_data_f_11__60_),
	.b(FE_OFN1085_n22923));
   oa12s01 U22991 (.o(n6633),
	.a(n23396),
	.b(FE_OFN1085_n22923),
	.c(n23938));
   oa12s01 U22992 (.o(n6638),
	.a(n23404),
	.b(FE_OFN1085_n22923),
	.c(n23936));
   na02s01 U22993 (.o(n23404),
	.a(proc_input_NIB_storage_data_f_11__58_),
	.b(FE_OFN1085_n22923));
   oa12s01 U22994 (.o(n6643),
	.a(n23290),
	.b(n22923),
	.c(n23932));
   na02s01 U22995 (.o(n23290),
	.a(proc_input_NIB_storage_data_f_11__57_),
	.b(FE_OFN1085_n22923));
   oa12s01 U22996 (.o(n6648),
	.a(n23391),
	.b(FE_OFN1085_n22923),
	.c(n23930));
   na02s01 U22997 (.o(n23391),
	.a(proc_input_NIB_storage_data_f_11__56_),
	.b(FE_OFN1085_n22923));
   oa12s01 U22998 (.o(n6653),
	.a(n23403),
	.b(FE_OFN1085_n22923),
	.c(n23910));
   na02s01 U22999 (.o(n23403),
	.a(proc_input_NIB_storage_data_f_11__55_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23000 (.o(n6658),
	.a(n23395),
	.b(FE_OFN1085_n22923),
	.c(n23924));
   oa12s01 U23001 (.o(n6663),
	.a(n23405),
	.b(FE_OFN1085_n22923),
	.c(n23922));
   na02s01 U23002 (.o(n23405),
	.a(proc_input_NIB_storage_data_f_11__53_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23003 (.o(n6668),
	.a(n23380),
	.b(FE_OFN1085_n22923),
	.c(n23890));
   oa12s01 U23004 (.o(n6673),
	.a(n23401),
	.b(FE_OFN1085_n22923),
	.c(n23947));
   na02s01 U23005 (.o(n23401),
	.a(proc_input_NIB_storage_data_f_11__51_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23006 (.o(n6678),
	.a(n23291),
	.b(FE_OFN1085_n22923),
	.c(n23903));
   na02s01 U23007 (.o(n23291),
	.a(proc_input_NIB_storage_data_f_11__50_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23008 (.o(n6683),
	.a(n23289),
	.b(n22778),
	.c(n23908));
   na02s01 U23009 (.o(n23289),
	.a(proc_input_NIB_storage_data_f_11__49_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23010 (.o(n6688),
	.a(n23382),
	.b(FE_OFN1085_n22923),
	.c(n23912));
   na02s01 U23011 (.o(n23382),
	.a(proc_input_NIB_storage_data_f_11__48_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23012 (.o(n6693),
	.a(n22815),
	.b(FE_OFN1086_n22923),
	.c(n23914));
   na02s01 U23013 (.o(n22815),
	.a(proc_input_NIB_storage_data_f_11__47_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23014 (.o(n6698),
	.a(n23381),
	.b(FE_OFN1085_n22923),
	.c(n23916));
   na02s01 U23015 (.o(n23381),
	.a(proc_input_NIB_storage_data_f_11__46_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23016 (.o(n6703),
	.a(n22814),
	.b(FE_OFN1086_n22923),
	.c(n23942));
   na02s01 U23017 (.o(n22814),
	.a(proc_input_NIB_storage_data_f_11__45_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23018 (.o(n6708),
	.a(n22812),
	.b(FE_OFN1086_n22923),
	.c(n23920));
   na02s01 U23019 (.o(n22812),
	.a(proc_input_NIB_storage_data_f_11__44_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23020 (.o(n6713),
	.a(n22816),
	.b(FE_OFN1086_n22923),
	.c(n23806));
   na02s01 U23021 (.o(n22816),
	.a(proc_input_NIB_storage_data_f_11__43_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23022 (.o(n6718),
	.a(n22818),
	.b(FE_OFN1085_n22923),
	.c(n23808));
   na02s01 U23023 (.o(n22818),
	.a(proc_input_NIB_storage_data_f_11__42_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23024 (.o(n6723),
	.a(n22813),
	.b(FE_OFN1086_n22923),
	.c(n23928));
   na02s01 U23025 (.o(n22813),
	.a(proc_input_NIB_storage_data_f_11__41_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23026 (.o(n6728),
	.a(n22811),
	.b(FE_OFN1086_n22923),
	.c(n23800));
   na02s01 U23027 (.o(n22811),
	.a(proc_input_NIB_storage_data_f_11__40_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23028 (.o(n6733),
	.a(n22924),
	.b(FE_OFN426_n22778),
	.c(n23934));
   na02s01 U23029 (.o(n22924),
	.a(proc_input_NIB_storage_data_f_11__39_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23030 (.o(n6738),
	.a(n22921),
	.b(FE_OFN427_n22778),
	.c(n23812));
   oa12s01 U23031 (.o(n6743),
	.a(n22817),
	.b(FE_OFN1085_n22923),
	.c(n23796));
   na02s01 U23032 (.o(n22817),
	.a(proc_input_NIB_storage_data_f_11__37_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23033 (.o(n6748),
	.a(n23402),
	.b(FE_OFN1086_n22923),
	.c(n23940));
   na02s01 U23034 (.o(n23402),
	.a(proc_input_NIB_storage_data_f_11__36_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23035 (.o(n6753),
	.a(n22918),
	.b(FE_OFN426_n22778),
	.c(n23944));
   na02s01 U23036 (.o(n22918),
	.a(proc_input_NIB_storage_data_f_11__35_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23037 (.o(n6758),
	.a(n22920),
	.b(FE_OFN427_n22778),
	.c(n23816));
   na02s01 U23038 (.o(n22920),
	.a(proc_input_NIB_storage_data_f_11__34_),
	.b(FE_OFN1086_n22923));
   oa22s01 U23039 (.o(n22795),
	.a(FE_OFN1086_n22923),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_11__33_),
	.d(n22779));
   oa12s01 U23040 (.o(n6768),
	.a(n23288),
	.b(FE_OFN427_n22778),
	.c(n23905));
   na02s01 U23041 (.o(n23288),
	.a(proc_input_NIB_storage_data_f_11__32_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23042 (.o(n6773),
	.a(n22919),
	.b(n22923),
	.c(n23791));
   na02s01 U23043 (.o(n22919),
	.a(proc_input_NIB_storage_data_f_11__31_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23044 (.o(n6778),
	.a(n22922),
	.b(n22778),
	.c(n23894));
   na02s01 U23045 (.o(n22922),
	.a(proc_input_NIB_storage_data_f_11__30_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23046 (.o(n6783),
	.a(n23390),
	.b(FE_OFN1085_n22923),
	.c(n23804));
   na02s01 U23047 (.o(n23390),
	.a(proc_input_NIB_storage_data_f_11__29_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23048 (.o(n6788),
	.a(n23379),
	.b(n22778),
	.c(n23814));
   na02s01 U23049 (.o(n23379),
	.a(proc_input_NIB_storage_data_f_11__28_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23050 (.o(n6793),
	.a(n23383),
	.b(FE_OFN426_n22778),
	.c(n23822));
   na02s01 U23051 (.o(n23383),
	.a(proc_input_NIB_storage_data_f_11__27_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23052 (.o(n6798),
	.a(n23387),
	.b(FE_OFN1085_n22923),
	.c(n23818));
   na02s01 U23053 (.o(n23387),
	.a(proc_input_NIB_storage_data_f_11__26_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23054 (.o(n6803),
	.a(n23386),
	.b(FE_OFN426_n22778),
	.c(n23802));
   na02s01 U23055 (.o(n23386),
	.a(proc_input_NIB_storage_data_f_11__25_),
	.b(FE_OFN1086_n22923));
   oa12s01 U23056 (.o(n6808),
	.a(n23385),
	.b(FE_OFN1085_n22923),
	.c(n23798));
   na02s01 U23057 (.o(n23385),
	.a(proc_input_NIB_storage_data_f_11__24_),
	.b(FE_OFN1085_n22923));
   oa12s01 U23058 (.o(n6813),
	.a(n23384),
	.b(FE_OFN427_n22778),
	.c(n23793));
   oa12s01 U23059 (.o(n6818),
	.a(n23388),
	.b(FE_OFN1086_n22923),
	.c(n23820));
   na02s01 U23060 (.o(n23388),
	.a(proc_input_NIB_storage_data_f_11__22_),
	.b(FE_OFN1086_n22923));
   oa22s01 U23061 (.o(n22789),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_11__21_),
	.d(n22779));
   oa22s01 U23062 (.o(n22780),
	.a(FE_OFN1086_n22923),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_11__20_),
	.d(n22779));
   oa22s01 U23063 (.o(n22798),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_11__19_),
	.d(n22779));
   oa22s01 U23064 (.o(n22782),
	.a(FE_OFN1086_n22923),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_11__18_),
	.d(n22779));
   oa22s01 U23065 (.o(n22785),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_11__17_),
	.d(n22779));
   oa22s01 U23066 (.o(n22790),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_11__16_),
	.d(n22779));
   oa22s01 U23067 (.o(n22801),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_11__15_),
	.d(n22779));
   oa22s01 U23068 (.o(n22796),
	.a(FE_OFN1086_n22923),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_11__14_),
	.d(n22779));
   oa22s01 U23069 (.o(n22794),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_11__13_),
	.d(n22779));
   oa22s01 U23070 (.o(n22793),
	.a(FE_OFN1086_n22923),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_11__12_),
	.d(n22779));
   oa22s01 U23071 (.o(n22787),
	.a(FE_OFN1086_n22923),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_11__11_),
	.d(n22779));
   oa22s01 U23072 (.o(n22797),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_11__9_),
	.d(n22779));
   oa22s01 U23073 (.o(n22788),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_11__8_),
	.d(n22779));
   oa22s01 U23074 (.o(n22800),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_11__7_),
	.d(n22779));
   oa22s01 U23075 (.o(n22781),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_11__6_),
	.d(n22779));
   oa22s01 U23076 (.o(n22783),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_11__5_),
	.d(n22779));
   oa22s01 U23077 (.o(n22792),
	.a(FE_OFN1086_n22923),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_11__4_),
	.d(n22779));
   oa22s01 U23078 (.o(n22786),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_11__3_),
	.d(n22779));
   oa22s01 U23079 (.o(n22791),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_11__2_),
	.d(n22779));
   oa22s01 U23080 (.o(n22799),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_11__1_),
	.d(n22779));
   oa22s01 U23081 (.o(n22802),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_11__0_),
	.d(n22779));
   oa12s01 U23082 (.o(n7893),
	.a(n22282),
	.b(FE_OFN585_n25643),
	.c(n23827));
   na02s01 U23083 (.o(n22282),
	.a(proc_input_NIB_storage_data_f_15__63_),
	.b(FE_OFN585_n25643));
   oa12s01 U23084 (.o(n7898),
	.a(n22276),
	.b(n17768),
	.c(n23810));
   na02s01 U23085 (.o(n22276),
	.a(proc_input_NIB_storage_data_f_15__62_),
	.b(n17768));
   oa12s01 U23086 (.o(n7903),
	.a(n23284),
	.b(n17768),
	.c(n23918));
   oa12s01 U23087 (.o(n7908),
	.a(n23271),
	.b(n17768),
	.c(n23926));
   na02s01 U23088 (.o(n23271),
	.a(proc_input_NIB_storage_data_f_15__60_),
	.b(n17768));
   oa12s01 U23089 (.o(n7913),
	.a(n23269),
	.b(n17768),
	.c(n23938));
   na02s01 U23090 (.o(n23269),
	.a(proc_input_NIB_storage_data_f_15__59_),
	.b(n17768));
   oa12s01 U23091 (.o(n7918),
	.a(n23267),
	.b(n17768),
	.c(n23936));
   na02s01 U23092 (.o(n23267),
	.a(proc_input_NIB_storage_data_f_15__58_),
	.b(n17768));
   oa12s01 U23093 (.o(n7923),
	.a(n23283),
	.b(FE_OFN585_n25643),
	.c(n23932));
   na02s01 U23094 (.o(n23283),
	.a(proc_input_NIB_storage_data_f_15__57_),
	.b(FE_OFN585_n25643));
   oa12s01 U23095 (.o(n7928),
	.a(n23277),
	.b(FE_OFN585_n25643),
	.c(n23930));
   na02s01 U23096 (.o(n23277),
	.a(proc_input_NIB_storage_data_f_15__56_),
	.b(FE_OFN585_n25643));
   oa12s01 U23097 (.o(n7933),
	.a(n23285),
	.b(FE_OFN585_n25643),
	.c(n23910));
   na02s01 U23098 (.o(n23285),
	.a(proc_input_NIB_storage_data_f_15__55_),
	.b(FE_OFN585_n25643));
   oa12s01 U23099 (.o(n7938),
	.a(n23279),
	.b(FE_OFN585_n25643),
	.c(n23924));
   na02s01 U23100 (.o(n23279),
	.a(proc_input_NIB_storage_data_f_15__54_),
	.b(FE_OFN585_n25643));
   oa12s01 U23101 (.o(n7943),
	.a(n23274),
	.b(FE_OFN585_n25643),
	.c(n23922));
   na02s01 U23102 (.o(n23274),
	.a(proc_input_NIB_storage_data_f_15__53_),
	.b(FE_OFN585_n25643));
   oa12s01 U23103 (.o(n7948),
	.a(n23276),
	.b(FE_OFN585_n25643),
	.c(n23890));
   na02s01 U23104 (.o(n23276),
	.a(proc_input_NIB_storage_data_f_15__52_),
	.b(FE_OFN585_n25643));
   oa12s01 U23105 (.o(n7953),
	.a(n23287),
	.b(n17768),
	.c(n23947));
   na02s01 U23106 (.o(n23287),
	.a(proc_input_NIB_storage_data_f_15__51_),
	.b(n17768));
   oa12s01 U23107 (.o(n7958),
	.a(n23282),
	.b(FE_OFN585_n25643),
	.c(n23903));
   na02s01 U23108 (.o(n23282),
	.a(proc_input_NIB_storage_data_f_15__50_),
	.b(FE_OFN585_n25643));
   oa12f01 U23109 (.o(n7963),
	.a(n23266),
	.b(n17768),
	.c(n23908));
   na02s01 U23110 (.o(n23266),
	.a(proc_input_NIB_storage_data_f_15__49_),
	.b(n17768));
   oa12f01 U23111 (.o(n7968),
	.a(n23268),
	.b(n17768),
	.c(n23912));
   na02s01 U23112 (.o(n23268),
	.a(proc_input_NIB_storage_data_f_15__48_),
	.b(n17768));
   oa12s01 U23113 (.o(n7973),
	.a(n23280),
	.b(FE_OFN585_n25643),
	.c(n23914));
   na02s01 U23114 (.o(n23280),
	.a(proc_input_NIB_storage_data_f_15__47_),
	.b(FE_OFN585_n25643));
   oa12f01 U23115 (.o(n7978),
	.a(n23270),
	.b(n17768),
	.c(n23916));
   oa12s01 U23116 (.o(n7983),
	.a(n23265),
	.b(FE_OFN585_n25643),
	.c(n23942));
   na02s01 U23117 (.o(n23265),
	.a(proc_input_NIB_storage_data_f_15__45_),
	.b(FE_OFN585_n25643));
   oa12s01 U23118 (.o(n7988),
	.a(n23272),
	.b(FE_OFN585_n25643),
	.c(n23920));
   na02s01 U23119 (.o(n23272),
	.a(proc_input_NIB_storage_data_f_15__44_),
	.b(FE_OFN585_n25643));
   oa12f01 U23120 (.o(n7993),
	.a(n22274),
	.b(FE_OFN585_n25643),
	.c(n23806));
   na02s01 U23121 (.o(n22274),
	.a(proc_input_NIB_storage_data_f_15__43_),
	.b(FE_OFN585_n25643));
   oa12f01 U23122 (.o(n7998),
	.a(n22809),
	.b(n17768),
	.c(n23808));
   na02s01 U23123 (.o(n22809),
	.a(proc_input_NIB_storage_data_f_15__42_),
	.b(n17768));
   oa12s01 U23124 (.o(n8003),
	.a(n23273),
	.b(FE_OFN585_n25643),
	.c(n23928));
   na02s01 U23125 (.o(n23273),
	.a(proc_input_NIB_storage_data_f_15__41_),
	.b(FE_OFN585_n25643));
   oa12s01 U23126 (.o(n8008),
	.a(n22806),
	.b(FE_OFN585_n25643),
	.c(n23800));
   na02s01 U23127 (.o(n22806),
	.a(proc_input_NIB_storage_data_f_15__40_),
	.b(FE_OFN585_n25643));
   oa12s01 U23128 (.o(n8013),
	.a(n23286),
	.b(FE_OFN585_n25643),
	.c(n23934));
   na02s01 U23129 (.o(n23286),
	.a(proc_input_NIB_storage_data_f_15__39_),
	.b(FE_OFN585_n25643));
   oa12f01 U23130 (.o(n8018),
	.a(n23275),
	.b(FE_OFN585_n25643),
	.c(n23812));
   na02s01 U23131 (.o(n23275),
	.a(proc_input_NIB_storage_data_f_15__38_),
	.b(FE_OFN585_n25643));
   oa12f01 U23132 (.o(n8023),
	.a(n22807),
	.b(n17768),
	.c(n23796));
   na02s01 U23133 (.o(n22807),
	.a(proc_input_NIB_storage_data_f_15__37_),
	.b(n17768));
   oa12s01 U23134 (.o(n8028),
	.a(n22803),
	.b(FE_OFN585_n25643),
	.c(n23940));
   na02s01 U23135 (.o(n22803),
	.a(proc_input_NIB_storage_data_f_15__36_),
	.b(FE_OFN585_n25643));
   oa12f01 U23136 (.o(n8033),
	.a(n22275),
	.b(FE_OFN585_n25643),
	.c(n23944));
   na02s01 U23137 (.o(n22275),
	.a(proc_input_NIB_storage_data_f_15__35_),
	.b(FE_OFN585_n25643));
   oa12s01 U23138 (.o(n8038),
	.a(n23281),
	.b(FE_OFN585_n25643),
	.c(n23816));
   na02s01 U23139 (.o(n23281),
	.a(proc_input_NIB_storage_data_f_15__34_),
	.b(FE_OFN585_n25643));
   oa12s01 U23140 (.o(n8048),
	.a(n23264),
	.b(FE_OFN585_n25643),
	.c(n23905));
   na02s01 U23141 (.o(n23264),
	.a(proc_input_NIB_storage_data_f_15__32_),
	.b(FE_OFN585_n25643));
   oa12s01 U23142 (.o(n8053),
	.a(n22278),
	.b(FE_OFN585_n25643),
	.c(n23791));
   na02s01 U23143 (.o(n22278),
	.a(proc_input_NIB_storage_data_f_15__31_),
	.b(FE_OFN585_n25643));
   oa12f01 U23144 (.o(n8058),
	.a(n23278),
	.b(n17768),
	.c(n23894));
   na02s01 U23145 (.o(n23278),
	.a(proc_input_NIB_storage_data_f_15__30_),
	.b(n17768));
   oa12f01 U23146 (.o(n8063),
	.a(n22277),
	.b(n17768),
	.c(n23804));
   na02s01 U23147 (.o(n22277),
	.a(proc_input_NIB_storage_data_f_15__29_),
	.b(n17768));
   oa12s01 U23148 (.o(n8068),
	.a(n22281),
	.b(FE_OFN585_n25643),
	.c(n23814));
   na02s01 U23149 (.o(n22281),
	.a(proc_input_NIB_storage_data_f_15__28_),
	.b(FE_OFN585_n25643));
   oa12s01 U23150 (.o(n8073),
	.a(n22808),
	.b(FE_OFN585_n25643),
	.c(n23822));
   na02s01 U23151 (.o(n22808),
	.a(proc_input_NIB_storage_data_f_15__27_),
	.b(FE_OFN585_n25643));
   oa12f01 U23152 (.o(n8078),
	.a(n22279),
	.b(n17768),
	.c(n23818));
   na02s01 U23153 (.o(n22279),
	.a(proc_input_NIB_storage_data_f_15__26_),
	.b(n17768));
   oa12s01 U23154 (.o(n8083),
	.a(n22280),
	.b(FE_OFN585_n25643),
	.c(n23802));
   na02s01 U23155 (.o(n22280),
	.a(proc_input_NIB_storage_data_f_15__25_),
	.b(FE_OFN585_n25643));
   oa12f01 U23156 (.o(n8088),
	.a(n22805),
	.b(n17768),
	.c(n23798));
   na02s01 U23157 (.o(n22805),
	.a(proc_input_NIB_storage_data_f_15__24_),
	.b(n17768));
   oa12f01 U23158 (.o(n8093),
	.a(n22804),
	.b(FE_OFN585_n25643),
	.c(n23793));
   na02s01 U23159 (.o(n22804),
	.a(proc_input_NIB_storage_data_f_15__23_),
	.b(FE_OFN585_n25643));
   oa12s01 U23160 (.o(n8098),
	.a(n22810),
	.b(FE_OFN585_n25643),
	.c(n23820));
   na02s01 U23161 (.o(n22810),
	.a(proc_input_NIB_storage_data_f_15__22_),
	.b(FE_OFN585_n25643));
   oa22s01 U23162 (.o(n25624),
	.a(n17768),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_15__19_),
	.d(n25643));
   oa22s01 U23163 (.o(n25625),
	.a(FE_OFN585_n25643),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_15__18_),
	.d(n25643));
   oa22s01 U23164 (.o(n25626),
	.a(n17768),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_15__17_),
	.d(n25643));
   oa22s01 U23165 (.o(n25627),
	.a(FE_OFN585_n25643),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_15__16_),
	.d(n25643));
   oa22f01 U23166 (.o(n25628),
	.a(n17768),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_15__15_),
	.d(n25643));
   oa22s01 U23167 (.o(n25629),
	.a(FE_OFN585_n25643),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_15__14_),
	.d(n25643));
   oa22f01 U23168 (.o(n25630),
	.a(n17768),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_15__13_),
	.d(n25643));
   oa22s01 U23169 (.o(n25632),
	.a(FE_OFN585_n25643),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_15__11_),
	.d(n25643));
   ao22s01 U23170 (.o(n25927),
	.a(validIn_W),
	.b(n25928),
	.c(west_input_NIB_tail_ptr_f_0_),
	.d(n25929));
   oa22s01 U23171 (.o(n24847),
	.a(FE_OFN896_n17769),
	.b(dataIn_S_21_),
	.c(south_input_NIB_storage_data_f_3__21_),
	.d(n20996));
   oa22s01 U23172 (.o(n24838),
	.a(n17769),
	.b(dataIn_S_19_),
	.c(south_input_NIB_storage_data_f_3__19_),
	.d(n20996));
   oa22s01 U23173 (.o(n24848),
	.a(n17769),
	.b(dataIn_S_18_),
	.c(south_input_NIB_storage_data_f_3__18_),
	.d(n20996));
   oa22s01 U23174 (.o(n24837),
	.a(n17769),
	.b(dataIn_S_16_),
	.c(south_input_NIB_storage_data_f_3__16_),
	.d(n20996));
   oa22s01 U23175 (.o(n24844),
	.a(n17769),
	.b(dataIn_S_14_),
	.c(south_input_NIB_storage_data_f_3__14_),
	.d(n20996));
   oa22s01 U23176 (.o(n24841),
	.a(n17769),
	.b(dataIn_S_13_),
	.c(south_input_NIB_storage_data_f_3__13_),
	.d(n20996));
   oa22s01 U23177 (.o(n22401),
	.a(n17769),
	.b(dataIn_S_11_),
	.c(south_input_NIB_storage_data_f_3__11_),
	.d(n20996));
   oa22s01 U23178 (.o(n22411),
	.a(n17769),
	.b(dataIn_S_10_),
	.c(south_input_NIB_storage_data_f_3__10_),
	.d(n20996));
   oa22s01 U23179 (.o(n22395),
	.a(FE_OFN896_n17769),
	.b(dataIn_S_9_),
	.c(south_input_NIB_storage_data_f_3__9_),
	.d(n20996));
   oa22s01 U23180 (.o(n22404),
	.a(FE_OFN896_n17769),
	.b(dataIn_S_7_),
	.c(south_input_NIB_storage_data_f_3__7_),
	.d(n20996));
   oa22s01 U23181 (.o(n22403),
	.a(n17769),
	.b(dataIn_S_6_),
	.c(south_input_NIB_storage_data_f_3__6_),
	.d(n20996));
   oa22s01 U23182 (.o(n22402),
	.a(FE_OFN896_n17769),
	.b(dataIn_S_5_),
	.c(south_input_NIB_storage_data_f_3__5_),
	.d(n20996));
   oa22s01 U23183 (.o(n22412),
	.a(n17769),
	.b(dataIn_S_4_),
	.c(south_input_NIB_storage_data_f_3__4_),
	.d(n20996));
   oa22s01 U23184 (.o(n22399),
	.a(FE_OFN896_n17769),
	.b(dataIn_S_3_),
	.c(south_input_NIB_storage_data_f_3__3_),
	.d(n20996));
   oa22s01 U23185 (.o(n22398),
	.a(n17769),
	.b(dataIn_S_2_),
	.c(south_input_NIB_storage_data_f_3__2_),
	.d(n20996));
   oa22s01 U23186 (.o(n22396),
	.a(n17769),
	.b(dataIn_S_1_),
	.c(south_input_NIB_storage_data_f_3__1_),
	.d(n20996));
   oa22s01 U23187 (.o(n22405),
	.a(FE_OFN896_n17769),
	.b(dataIn_S_0_),
	.c(south_input_NIB_storage_data_f_3__0_),
	.d(n20996));
   oa22s01 U23188 (.o(n25662),
	.a(n25881),
	.b(dataIn_E_33_),
	.c(east_input_NIB_storage_data_f_1__33_),
	.d(n24761));
   oa12s01 U23189 (.o(n11288),
	.a(n24886),
	.b(n24761),
	.c(n24887));
   oa12s01 U23190 (.o(n11303),
	.a(n24884),
	.b(n24761),
	.c(n24885));
   oa12s01 U23191 (.o(n11308),
	.a(n24870),
	.b(n24761),
	.c(n24871));
   oa12s01 U23192 (.o(n11318),
	.a(n24880),
	.b(n24761),
	.c(n24881));
   oa12s01 U23193 (.o(n11323),
	.a(n24878),
	.b(n24761),
	.c(n24879));
   oa12s01 U23194 (.o(n11328),
	.a(n24876),
	.b(n24761),
	.c(n24877));
   oa12s01 U23195 (.o(n11333),
	.a(n24874),
	.b(n24761),
	.c(n24875));
   oa12s01 U23196 (.o(n11338),
	.a(n24872),
	.b(n24761),
	.c(n24873));
   oa22s01 U23197 (.o(n25663),
	.a(n25881),
	.b(dataIn_E_21_),
	.c(east_input_NIB_storage_data_f_1__21_),
	.d(n24761));
   oa22s01 U23198 (.o(n25664),
	.a(n25881),
	.b(dataIn_E_20_),
	.c(east_input_NIB_storage_data_f_1__20_),
	.d(n24761));
   oa22s01 U23199 (.o(n25665),
	.a(n25881),
	.b(dataIn_E_19_),
	.c(east_input_NIB_storage_data_f_1__19_),
	.d(n24761));
   oa22s01 U23200 (.o(n25666),
	.a(n25881),
	.b(dataIn_E_18_),
	.c(east_input_NIB_storage_data_f_1__18_),
	.d(FE_OFN556_n24761));
   oa22s01 U23201 (.o(n25667),
	.a(n25881),
	.b(dataIn_E_17_),
	.c(east_input_NIB_storage_data_f_1__17_),
	.d(n24761));
   oa22s01 U23202 (.o(n25668),
	.a(n25881),
	.b(dataIn_E_15_),
	.c(east_input_NIB_storage_data_f_1__15_),
	.d(n24761));
   oa22s01 U23203 (.o(n25669),
	.a(n25881),
	.b(dataIn_E_13_),
	.c(east_input_NIB_storage_data_f_1__13_),
	.d(n24761));
   oa22s01 U23204 (.o(n25670),
	.a(n25881),
	.b(dataIn_E_12_),
	.c(east_input_NIB_storage_data_f_1__12_),
	.d(n24761));
   oa22s01 U23205 (.o(n25671),
	.a(n25881),
	.b(dataIn_E_11_),
	.c(east_input_NIB_storage_data_f_1__11_),
	.d(n24761));
   oa22s01 U23206 (.o(n25672),
	.a(n25881),
	.b(dataIn_E_10_),
	.c(east_input_NIB_storage_data_f_1__10_),
	.d(n24761));
   oa22s01 U23207 (.o(n25673),
	.a(n25881),
	.b(dataIn_E_9_),
	.c(east_input_NIB_storage_data_f_1__9_),
	.d(n24761));
   oa22s01 U23208 (.o(n25674),
	.a(n25881),
	.b(dataIn_E_8_),
	.c(east_input_NIB_storage_data_f_1__8_),
	.d(FE_OFN556_n24761));
   oa22s01 U23209 (.o(n25675),
	.a(n25881),
	.b(dataIn_E_7_),
	.c(east_input_NIB_storage_data_f_1__7_),
	.d(n24761));
   oa22s01 U23210 (.o(n25676),
	.a(n25881),
	.b(dataIn_E_6_),
	.c(east_input_NIB_storage_data_f_1__6_),
	.d(n24761));
   oa22s01 U23211 (.o(n25677),
	.a(n25881),
	.b(dataIn_E_4_),
	.c(east_input_NIB_storage_data_f_1__4_),
	.d(n24761));
   oa22s01 U23212 (.o(n25678),
	.a(n25881),
	.b(dataIn_E_1_),
	.c(east_input_NIB_storage_data_f_1__1_),
	.d(FE_OFN556_n24761));
   na02s01 U23213 (.o(n25209),
	.a(east_input_NIB_storage_data_f_3__54_),
	.b(n24921));
   oa12s01 U23214 (.o(n11843),
	.a(n24934),
	.b(n24921),
	.c(n24935));
   oa12s01 U23215 (.o(n11848),
	.a(n24926),
	.b(n24921),
	.c(n24927));
   oa12s01 U23216 (.o(n11853),
	.a(n24948),
	.b(n24921),
	.c(n24949));
   oa12s01 U23217 (.o(n11858),
	.a(n24950),
	.b(n24921),
	.c(n24951));
   oa12s01 U23218 (.o(n11863),
	.a(n24944),
	.b(n24921),
	.c(n24945));
   oa12s01 U23219 (.o(n11868),
	.a(n24946),
	.b(n24921),
	.c(n24947));
   oa12s01 U23220 (.o(n11873),
	.a(n24922),
	.b(n24921),
	.c(n24923));
   oa12s01 U23221 (.o(n11878),
	.a(n24936),
	.b(n24921),
	.c(n24937));
   oa12s01 U23222 (.o(n11888),
	.a(n24930),
	.b(n24921),
	.c(n24931));
   oa12s01 U23223 (.o(n11898),
	.a(n24928),
	.b(n24921),
	.c(n24929));
   oa12s01 U23224 (.o(n11903),
	.a(n24940),
	.b(n24921),
	.c(n24941));
   oa12s01 U23225 (.o(n11908),
	.a(n24942),
	.b(n24921),
	.c(n24943));
   oa12s01 U23226 (.o(n11913),
	.a(n24938),
	.b(n24921),
	.c(n24939));
   oa12s01 U23227 (.o(n11918),
	.a(n24924),
	.b(n24921),
	.c(n24925));
   oa22s01 U23228 (.o(n25696),
	.a(FE_OFN24818_n24921),
	.b(dataIn_E_33_),
	.c(east_input_NIB_storage_data_f_3__33_),
	.d(FE_OFN940_n24921));
   oa22s01 U23229 (.o(n25697),
	.a(FE_OFN24824_n24921),
	.b(dataIn_E_21_),
	.c(east_input_NIB_storage_data_f_3__21_),
	.d(FE_OFN940_n24921));
   oa22s01 U23230 (.o(n25698),
	.a(FE_OFN942_n24921),
	.b(dataIn_E_20_),
	.c(east_input_NIB_storage_data_f_3__20_),
	.d(FE_OFN940_n24921));
   oa22s01 U23231 (.o(n25699),
	.a(FE_OFN24823_n24921),
	.b(dataIn_E_19_),
	.c(east_input_NIB_storage_data_f_3__19_),
	.d(FE_OFN940_n24921));
   oa22s01 U23232 (.o(n25700),
	.a(FE_OFN24823_n24921),
	.b(dataIn_E_18_),
	.c(east_input_NIB_storage_data_f_3__18_),
	.d(FE_OFN940_n24921));
   oa22s01 U23233 (.o(n25701),
	.a(FE_OFN24818_n24921),
	.b(dataIn_E_17_),
	.c(east_input_NIB_storage_data_f_3__17_),
	.d(FE_OFN940_n24921));
   oa22s01 U23234 (.o(n25702),
	.a(n25869),
	.b(dataIn_E_15_),
	.c(east_input_NIB_storage_data_f_3__15_),
	.d(FE_OFN940_n24921));
   oa22s01 U23235 (.o(n25703),
	.a(FE_OFN24818_n24921),
	.b(dataIn_E_13_),
	.c(east_input_NIB_storage_data_f_3__13_),
	.d(FE_OFN940_n24921));
   oa22s01 U23236 (.o(n25704),
	.a(FE_OFN942_n24921),
	.b(dataIn_E_12_),
	.c(east_input_NIB_storage_data_f_3__12_),
	.d(FE_OFN940_n24921));
   oa22s01 U23237 (.o(n25705),
	.a(FE_OFN24821_n24921),
	.b(dataIn_E_11_),
	.c(east_input_NIB_storage_data_f_3__11_),
	.d(FE_OFN940_n24921));
   oa22s01 U23238 (.o(n25706),
	.a(FE_OFN24816_n24921),
	.b(dataIn_E_10_),
	.c(east_input_NIB_storage_data_f_3__10_),
	.d(FE_OFN940_n24921));
   oa22s01 U23239 (.o(n25707),
	.a(FE_OFN24824_n24921),
	.b(dataIn_E_9_),
	.c(east_input_NIB_storage_data_f_3__9_),
	.d(FE_OFN940_n24921));
   oa22s01 U23240 (.o(n25708),
	.a(FE_OFN24824_n24921),
	.b(dataIn_E_8_),
	.c(east_input_NIB_storage_data_f_3__8_),
	.d(FE_OFN940_n24921));
   oa22s01 U23241 (.o(n25709),
	.a(FE_OFN24824_n24921),
	.b(dataIn_E_7_),
	.c(east_input_NIB_storage_data_f_3__7_),
	.d(FE_OFN940_n24921));
   oa22s01 U23242 (.o(n25710),
	.a(FE_OFN24822_n24921),
	.b(dataIn_E_6_),
	.c(east_input_NIB_storage_data_f_3__6_),
	.d(FE_OFN940_n24921));
   oa22s01 U23243 (.o(n25711),
	.a(FE_OFN24819_n24921),
	.b(dataIn_E_4_),
	.c(east_input_NIB_storage_data_f_3__4_),
	.d(FE_OFN940_n24921));
   oa22s01 U23244 (.o(n25712),
	.a(FE_OFN24824_n24921),
	.b(dataIn_E_1_),
	.c(east_input_NIB_storage_data_f_3__1_),
	.d(FE_OFN940_n24921));
   oa22s01 U23245 (.o(n24833),
	.a(n17771),
	.b(dataIn_N_33_),
	.c(north_input_NIB_storage_data_f_0__33_),
	.d(FE_OFN1092_n20934));
   ao22s01 U23246 (.o(n12313),
	.a(FE_OFN1092_n20934),
	.b(n25859),
	.c(n25858),
	.d(n17771));
   oa22s01 U23247 (.o(n24835),
	.a(n20934),
	.b(dataIn_N_20_),
	.c(north_input_NIB_storage_data_f_0__20_),
	.d(FE_OFN1092_n20934));
   ao22s01 U23248 (.o(n12323),
	.a(FE_OFN1092_n20934),
	.b(n25857),
	.c(n25856),
	.d(n17771));
   ao22s01 U23249 (.o(n12328),
	.a(FE_OFN1092_n20934),
	.b(n25855),
	.c(n25854),
	.d(n17771));
   oa22s01 U23250 (.o(n24830),
	.a(n17771),
	.b(dataIn_N_16_),
	.c(north_input_NIB_storage_data_f_0__16_),
	.d(FE_OFN1092_n20934));
   oa22s01 U23251 (.o(n24832),
	.a(n20934),
	.b(dataIn_N_15_),
	.c(north_input_NIB_storage_data_f_0__15_),
	.d(FE_OFN1092_n20934));
   oa22s01 U23252 (.o(n24831),
	.a(n17771),
	.b(dataIn_N_14_),
	.c(north_input_NIB_storage_data_f_0__14_),
	.d(FE_OFN1092_n20934));
   ao22s01 U23253 (.o(n12353),
	.a(FE_OFN1092_n20934),
	.b(n25853),
	.c(n25852),
	.d(n17771));
   oa22s01 U23254 (.o(n24829),
	.a(n20934),
	.b(dataIn_N_12_),
	.c(north_input_NIB_storage_data_f_0__12_),
	.d(FE_OFN1092_n20934));
   oa22s01 U23255 (.o(n25188),
	.a(n17771),
	.b(dataIn_N_11_),
	.c(north_input_NIB_storage_data_f_0__11_),
	.d(FE_OFN1092_n20934));
   oa22s01 U23256 (.o(n22339),
	.a(n17771),
	.b(dataIn_N_10_),
	.c(north_input_NIB_storage_data_f_0__10_),
	.d(FE_OFN1092_n20934));
   oa22s01 U23257 (.o(n22341),
	.a(n17771),
	.b(dataIn_N_9_),
	.c(north_input_NIB_storage_data_f_0__9_),
	.d(FE_OFN1092_n20934));
   oa22s01 U23258 (.o(n22337),
	.a(n17771),
	.b(dataIn_N_8_),
	.c(north_input_NIB_storage_data_f_0__8_),
	.d(FE_OFN1092_n20934));
   oa22s01 U23259 (.o(n22335),
	.a(n17771),
	.b(dataIn_N_7_),
	.c(north_input_NIB_storage_data_f_0__7_),
	.d(FE_OFN1092_n20934));
   ao22s01 U23260 (.o(n12388),
	.a(FE_OFN1092_n20934),
	.b(n25851),
	.c(n25850),
	.d(n17771));
   oa22s01 U23261 (.o(n22340),
	.a(n17771),
	.b(dataIn_N_4_),
	.c(north_input_NIB_storage_data_f_0__4_),
	.d(FE_OFN1092_n20934));
   oa22s01 U23262 (.o(n22333),
	.a(n17771),
	.b(dataIn_N_3_),
	.c(north_input_NIB_storage_data_f_0__3_),
	.d(FE_OFN1092_n20934));
   oa22s01 U23263 (.o(n22338),
	.a(n17771),
	.b(dataIn_N_2_),
	.c(north_input_NIB_storage_data_f_0__2_),
	.d(FE_OFN1092_n20934));
   oa22s01 U23264 (.o(n22334),
	.a(n17771),
	.b(dataIn_N_1_),
	.c(north_input_NIB_storage_data_f_0__1_),
	.d(FE_OFN1092_n20934));
   oa22s01 U23265 (.o(n22336),
	.a(n17771),
	.b(dataIn_N_0_),
	.c(north_input_NIB_storage_data_f_0__0_),
	.d(FE_OFN1092_n20934));
   no02f02 U23266 (.o(n18606),
	.a(n18607),
	.b(n18399));
   ao12m06 U23267 (.o(n25019),
	.a(n18647),
	.b(proc_output_space_is_one_f),
	.c(n22061));
   in01s01 U23268 (.o(n18405),
	.a(n18406));
   no02s01 U23269 (.o(n18406),
	.a(n18408),
	.b(n18407));
   na02s01 U23271 (.o(n19468),
	.a(n25979),
	.b(n25112));
   in01s01 U23272 (.o(n18408),
	.a(n19468));
   no02s01 U23273 (.o(n25377),
	.a(n25234),
	.b(n25929));
   no02s01 U23274 (.o(n20524),
	.a(east_input_NIB_elements_in_array_f_0_),
	.b(east_input_NIB_elements_in_array_f_1_));
   no02s01 U23275 (.o(n25343),
	.a(n25268),
	.b(n25897));
   na02s01 U23276 (.o(n18600),
	.a(east_input_NIB_elements_in_array_f_1_),
	.b(east_input_NIB_elements_in_array_f_0_));
   in01f03 U23277 (.o(n25129),
	.a(north_output_current_route_connection_2_));
   na03f20 U23278 (.o(n18064),
	.a(n18384),
	.b(n18383),
	.c(n19586));
   na04f20 U23279 (.o(n19627),
	.a(n18070),
	.b(n18069),
	.c(n18068),
	.d(n18065));
   ao22f08 U23280 (.o(n18067),
	.a(proc_input_NIB_storage_data_f_0__58_),
	.b(FE_OCPN25830_n),
	.c(proc_input_NIB_storage_data_f_13__58_),
	.d(n24454));
   ao22f08 U23281 (.o(n19583),
	.a(FE_OCPN25947_n19595),
	.b(proc_input_NIB_storage_data_f_15__61_),
	.c(proc_input_NIB_storage_data_f_5__61_),
	.d(FE_RN_49));
   ao22f06 U23282 (.o(n18417),
	.a(proc_input_NIB_storage_data_f_10__57_),
	.b(FE_OCPN25958_n18039),
	.c(proc_input_NIB_storage_data_f_5__57_),
	.d(FE_RN_49));
   ao22f02 U23283 (.o(n20066),
	.a(proc_input_NIB_storage_data_f_7__28_),
	.b(FE_OFN20_n17779),
	.c(proc_input_NIB_storage_data_f_5__28_),
	.d(FE_RN_49));
   no02f10 U23285 (.o(n20325),
	.a(east_output_control_planned_f),
	.b(validOut_E));
   no02f10 U23286 (.o(validOut_E),
	.a(n23400),
	.b(n20212));
   no03f08 U23287 (.o(n22865),
	.a(n19724),
	.b(n19723),
	.c(n18075));
   no04f08 U23288 (.o(n19731),
	.a(n19725),
	.b(n19724),
	.c(n19723),
	.d(n18075));
   na04f10 U23289 (.o(n18075),
	.a(n19687),
	.b(n19686),
	.c(n19684),
	.d(n19685));
   no02f10 U23290 (.o(n18225),
	.a(n19600),
	.b(n18076));
   na02f10 U23291 (.o(n18076),
	.a(n19598),
	.b(n19599));
   no02f08 U23292 (.o(n26020),
	.a(n20529),
	.b(n18392));
   ao22m02 U23293 (.o(n19745),
	.a(proc_input_NIB_storage_data_f_7__32_),
	.b(n17779),
	.c(proc_input_NIB_storage_data_f_5__32_),
	.d(FE_RN_49));
   ao22f02 U23294 (.o(n19771),
	.a(proc_input_NIB_storage_data_f_7__30_),
	.b(n17779),
	.c(proc_input_NIB_storage_data_f_5__30_),
	.d(FE_RN_49));
   ao22f08 U23295 (.o(n18081),
	.a(proc_input_NIB_storage_data_f_12__50_),
	.b(FE_OFN24803_n19500),
	.c(proc_input_NIB_storage_data_f_2__50_),
	.d(FE_OCPN25814_FE_OFN186_n24453));
   no04f20 U23296 (.o(n23184),
	.a(n18091),
	.b(n18090),
	.c(n18993),
	.d(n18089));
   in01f08 U23297 (.o(n18089),
	.a(n18991));
   no02f10 U23298 (.o(n18090),
	.a(n18995),
	.b(n18989));
   no02f08 U23299 (.o(n18091),
	.a(n24465),
	.b(n18992));
   na02f06 U23300 (.o(n18380),
	.a(n19737),
	.b(n20364));
   na03f04 U23301 (.o(n2843),
	.a(n25048),
	.b(n25047),
	.c(n25046));
   na02f10 U23302 (.o(n18093),
	.a(n19621),
	.b(n19620));
   no02f06 U23303 (.o(n20351),
	.a(n19475),
	.b(n19474));
   ao22f06 U23304 (.o(n19660),
	.a(FE_OCPN25959_n18039),
	.b(proc_input_NIB_storage_data_f_10__53_),
	.c(FE_OCPN25839_n24342),
	.d(proc_input_NIB_storage_data_f_0__53_));
   no02f04 U23305 (.o(n18095),
	.a(n18628),
	.b(n18059));
   oa12f08 U23306 (.o(n19464),
	.a(n19462),
	.b(n20147),
	.c(n19463));
   in01m01 U23307 (.o(n25070),
	.a(south_input_NIB_head_ptr_f_0_));
   na02f10 U23308 (.o(n19634),
	.a(n18160),
	.b(n18155));
   na03f40 U23309 (.o(n25516),
	.a(n18180),
	.b(n18179),
	.c(n18178));
   na04f04 U23310 (.o(n24962),
	.a(n24960),
	.b(n24959),
	.c(n24958),
	.d(n24957));
   in01f04 U23312 (.o(n18098),
	.a(n18059));
   in01f04 U23313 (.o(n18099),
	.a(n18098));
   ao22f10 U23314 (.o(n19525),
	.a(n19705),
	.b(proc_input_NIB_storage_data_f_9__39_),
	.c(FE_OCPN25950_n18039),
	.d(proc_input_NIB_storage_data_f_10__39_));
   ao22f04 U23315 (.o(n19684),
	.a(n20012),
	.b(proc_input_NIB_storage_data_f_9__48_),
	.c(FE_OCPN25949_n18039),
	.d(proc_input_NIB_storage_data_f_10__48_));
   no02f10 U23316 (.o(n18102),
	.a(n19616),
	.b(n19615));
   no02f10 U23317 (.o(n23548),
	.a(n19616),
	.b(n19615));
   no02f20 U23318 (.o(n20222),
	.a(n18382),
	.b(n18381));
   na02f20 U23319 (.o(n19632),
	.a(n18237),
	.b(n18234));
   in01s01 U23320 (.o(n18105),
	.a(FE_OCPN25965_proc_input_NIB_head_ptr_f_2));
   no02f10 U23321 (.o(n18155),
	.a(n18157),
	.b(n18156));
   na02f02 U23322 (.o(n2693),
	.a(n25426),
	.b(n25425));
   in01s01 U23323 (.o(n18106),
	.a(n25042));
   in01s01 U23324 (.o(n18107),
	.a(n18106));
   no04f03 U23325 (.o(n18275),
	.a(n18276),
	.b(n25132),
	.c(n25133),
	.d(n25131));
   no02f01 U23326 (.o(n21487),
	.a(n18258),
	.b(n18256));
   no02f01 U23327 (.o(n21490),
	.a(n18261),
	.b(n18259));
   no02s01 U23328 (.o(n22316),
	.a(n18267),
	.b(n18265));
   no02f01 U23329 (.o(n23320),
	.a(n18270),
	.b(n18268));
   in01s01 U23330 (.o(n18108),
	.a(n19910));
   in01f02 U23331 (.o(n18109),
	.a(n18108));
   ao12m02 U23332 (.o(n24158),
	.a(n18559),
	.b(FE_OCPN25834_n),
	.c(proc_input_NIB_storage_data_f_0__17_));
   no02s01 U23333 (.o(n25381),
	.a(west_input_NIB_elements_in_array_f_0_),
	.b(validIn_W));
   no02f01 U23334 (.o(n21713),
	.a(n18264),
	.b(n18262));
   no02f02 U23335 (.o(n20411),
	.a(n20409),
	.b(n23480));
   in01s01 U23336 (.o(n18616),
	.a(n25343));
   oa22m03 U23338 (.o(n20106),
	.a(proc_input_control_thanks_all_f),
	.b(proc_input_control_tail_last_f),
	.c(proc_input_control_count_one_f),
	.d(n21688));
   ao12f01 U23339 (.o(n21742),
	.a(n18561),
	.b(FE_OFN25644_n19504),
	.c(proc_input_NIB_storage_data_f_14__8_));
   ao12f01 U23341 (.o(n21317),
	.a(n18335),
	.b(FE_RN_13),
	.c(south_input_NIB_storage_data_f_3__5_));
   ao12f01 U23342 (.o(n24052),
	.a(n18345),
	.b(FE_OFN24741_n18683),
	.c(south_input_NIB_storage_data_f_1__3_));
   ao12f01 U23343 (.o(n24144),
	.a(n18337),
	.b(FE_RN_13),
	.c(south_input_NIB_storage_data_f_3__2_));
   in01s01 U23344 (.o(n18641),
	.a(n25377));
   in01s01 U23345 (.o(n18407),
	.a(n25044));
   ao12f02 U23346 (.o(n20319),
	.a(n19025),
	.b(n25506),
	.c(proc_input_valid));
   na02s01 U23347 (.o(n18599),
	.a(n20524),
	.b(validIn_E));
   in01s01 U23348 (.o(n18543),
	.a(n25019));
   na02f20 U23349 (.o(n25411),
	.a(n25050),
	.b(n25422));
   ao22f08 U23350 (.o(n19597),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__63_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__63_));
   na02f08 U23352 (.o(n25048),
	.a(n18107),
	.b(n18113));
   na02f10 U23353 (.o(n18113),
	.a(n25470),
	.b(n25469));
   oa22f02 U23354 (.o(n2853),
	.a(proc_input_NIB_elements_in_array_f_0_),
	.b(n25113),
	.c(n25112),
	.d(n18113));
   na02f10 U23355 (.o(n18847),
	.a(n18114),
	.b(n18846));
   oa22f06 U23356 (.o(n20439),
	.a(n18114),
	.b(n18870),
	.c(n18872),
	.d(n18871));
   ao22f08 U23357 (.o(n18114),
	.a(n18840),
	.b(n18845),
	.c(n18841),
	.d(n18842));
   in01f08 U23358 (.o(n18115),
	.a(n19742));
   na02f10 U23359 (.o(n18124),
	.a(n18115),
	.b(n18434));
   ao22f10 U23360 (.o(n18413),
	.a(proc_input_NIB_storage_data_f_14__57_),
	.b(n19769),
	.c(FE_OFN24803_n19500),
	.d(proc_input_NIB_storage_data_f_12__57_));
   na03f10 U23362 (.o(n18436),
	.a(n18422),
	.b(n19738),
	.c(n19549));
   na02f10 U23364 (.o(n18116),
	.a(n19043),
	.b(n18713));
   no02f10 U23365 (.o(n20227),
	.a(n18885),
	.b(n18118));
   in01f20 U23366 (.o(n18762),
	.a(n18714));
   no02f40 U23369 (.o(n19306),
	.a(east_input_NIB_head_ptr_f_1_),
	.b(n18391));
   na02f04 U23371 (.o(n19080),
	.a(FE_OFN24769_n19075),
	.b(north_input_NIB_storage_data_f_0__40_));
   no02f40 U23372 (.o(n19914),
	.a(east_input_NIB_head_ptr_f_0_),
	.b(n18442));
   na02f08 U23373 (.o(n18374),
	.a(FE_OFN65_n19542),
	.b(n23189));
   no03f04 U23374 (.o(n19858),
	.a(FE_OFN93_n21667),
	.b(n19860),
	.c(n19857));
   na02f10 U23375 (.o(n25009),
	.a(n20411),
	.b(n20410));
   oa22f02 U23376 (.o(proc_output_control_N467),
	.a(n18496),
	.b(n25423),
	.c(n25422),
	.d(n25421));
   ao22f20 U23377 (.o(n19590),
	.a(proc_input_NIB_storage_data_f_5__51_),
	.b(FE_RN_49),
	.c(proc_input_NIB_storage_data_f_15__51_),
	.d(FE_OCPN25947_n19595));
   ao22f10 U23378 (.o(n19667),
	.a(myChipID_f_4_),
	.b(n18120),
	.c(n21660),
	.d(FE_OFN53_n19355));
   na02f40 U23379 (.o(n19547),
	.a(n17789),
	.b(n17788));
   na02f08 U23380 (.o(n18173),
	.a(FE_RN_5),
	.b(west_input_NIB_storage_data_f_3__58_));
   oa22f04 U23381 (.o(n20180),
	.a(n20379),
	.b(n20165),
	.c(n20297),
	.d(n20164));
   na02f20 U23383 (.o(n19530),
	.a(FE_RN_24),
	.b(n18121));
   no04f20 U23384 (.o(n18558),
	.a(n18433),
	.b(n20215),
	.c(n18124),
	.d(n18122));
   na02f10 U23385 (.o(n18122),
	.a(n18435),
	.b(n18123));
   no02f04 U23386 (.o(n19860),
	.a(n22517),
	.b(n24968));
   in01f06 U23387 (.o(n20155),
	.a(n19121));
   oa22f10 U23388 (.o(n18734),
	.a(myLocY_f_6_),
	.b(n23186),
	.c(myLocY_f_5_),
	.d(n17751));
   oa12m02 U23389 (.o(n19852),
	.a(n19849),
	.b(n19851),
	.c(n19850));
   oa22f10 U23390 (.o(n18924),
	.a(n18923),
	.b(n24465),
	.c(FE_OFN30_n18974),
	.d(n18125));
   oa22f10 U23391 (.o(n18896),
	.a(n18895),
	.b(n24465),
	.c(FE_OFN30_n18974),
	.d(n18126));
   na04f20 U23393 (.o(n19408),
	.a(n19407),
	.b(n19406),
	.c(n19405),
	.d(n19404));
   no03f40 U23394 (.o(n20147),
	.a(n19410),
	.b(n19409),
	.c(FE_RN_20));
   no02f20 U23395 (.o(n19504),
	.a(n19505),
	.b(n25140));
   na02f20 U23396 (.o(n23508),
	.a(n18912),
	.b(n18911));
   na02f08 U23398 (.o(n18174),
	.a(n18960),
	.b(west_input_NIB_storage_data_f_2__58_));
   no02f80 U23399 (.o(n18960),
	.a(FE_OCPN25902_west_input_NIB_head_ptr_f_0),
	.b(FE_OCPN25820_west_input_NIB_head_ptr_f_1));
   na02f10 U23400 (.o(n18245),
	.a(n18247),
	.b(n18246));
   oa22f10 U23401 (.o(n19187),
	.a(n21408),
	.b(n19347),
	.c(myChipID_f_5_),
	.d(n21485));
   in01f10 U23402 (.o(n19200),
	.a(n19187));
   no02f40 U23404 (.o(n18131),
	.a(FE_RN_29),
	.b(n18533));
   no04f08 U23405 (.o(n20357),
	.a(n20356),
	.b(n20355),
	.c(n20528),
	.d(n20354));
   ao22f10 U23406 (.o(n19152),
	.a(n21865),
	.b(north_input_NIB_storage_data_f_2__51_),
	.c(FE_OFN25610_n19071),
	.d(north_input_NIB_storage_data_f_1__51_));
   no02f10 U23407 (.o(n19196),
	.a(n19387),
	.b(n23542));
   ao22f08 U23408 (.o(n19598),
	.a(n20056),
	.b(proc_input_NIB_storage_data_f_9__63_),
	.c(n17742),
	.d(proc_input_NIB_storage_data_f_4__63_));
   no02f10 U23409 (.o(n19035),
	.a(FE_RN_4),
	.b(n18132));
   ao22f02 U23410 (.o(n24991),
	.a(n24987),
	.b(n24986),
	.c(n24985),
	.d(n24984));
   na02f20 U23412 (.o(n21160),
	.a(n18685),
	.b(n18684));
   na02f20 U23413 (.o(n18532),
	.a(n19587),
	.b(n19589));
   na02f20 U23414 (.o(n18507),
	.a(n20127),
	.b(n18134));
   no02f20 U23415 (.o(n18134),
	.a(n25987),
	.b(n26017));
   na02f20 U23416 (.o(n18870),
	.a(n18830),
	.b(n18829));
   in01f20 U23417 (.o(n21315),
	.a(n18754));
   no02f10 U23418 (.o(n19170),
	.a(myChipID_f_6_),
	.b(n19168));
   in01f08 U23419 (.o(n18966),
	.a(n18964));
   no03f40 U23420 (.o(n23993),
	.a(n18898),
	.b(n18897),
	.c(n18896));
   na02f20 U23421 (.o(n23613),
	.a(n19167),
	.b(n19166));
   na02f20 U23422 (.o(n23612),
	.a(n18940),
	.b(n18939));
   na02f20 U23423 (.o(n24003),
	.a(n19175),
	.b(n19174));
   na02f40 U23425 (.o(n21748),
	.a(FE_OFN24743_n19499),
	.b(FE_OFN25607_n18151));
   no02f20 U23426 (.o(n19595),
	.a(n19505),
	.b(n25072));
   na02f20 U23427 (.o(n21332),
	.a(n18676),
	.b(n18675));
   ao22f04 U23428 (.o(n19512),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__40_),
	.c(n21768),
	.d(proc_input_NIB_storage_data_f_3__40_));
   oa22f02 U23429 (.o(north_output_control_N469),
	.a(n18454),
	.b(n18451),
	.c(n25137),
	.d(n25129));
   no02f10 U23430 (.o(n18411),
	.a(n18137),
	.b(n18136));
   na02f10 U23431 (.o(n18136),
	.a(n19027),
	.b(n19833));
   na02f20 U23433 (.o(n23994),
	.a(n19172),
	.b(n19171));
   na02f20 U23435 (.o(n18528),
	.a(n19585),
	.b(n19588));
   ao22f10 U23436 (.o(n19618),
	.a(n23548),
	.b(myChipID_f_10_),
	.c(n19617),
	.d(n23512));
   na03f08 U23437 (.o(n20146),
	.a(n19823),
	.b(FE_RN_6),
	.c(n18140));
   oa22f20 U23438 (.o(n19357),
	.a(myChipID_f_4_),
	.b(n23992),
	.c(n19635),
	.d(n23611));
   in01f10 U23439 (.o(n18888),
	.a(n21465));
   no02f20 U23440 (.o(n18892),
	.a(myChipID_f_3_),
	.b(n18888));
   ao12f10 U23441 (.o(n19197),
	.a(n19196),
	.b(n19387),
	.c(n23542));
   oa12f08 U23442 (.o(n25084),
	.a(n20473),
	.b(n20475),
	.c(FE_RN_2));
   na02f40 U23443 (.o(n21747),
	.a(FE_OFN24793_n17934),
	.b(FE_OCPN25946_n19501));
   ao22f20 U23445 (.o(n18582),
	.a(n24473),
	.b(south_input_NIB_storage_data_f_3__62_),
	.c(south_input_NIB_storage_data_f_0__62_),
	.d(FE_OFN24744_n18648));
   na02f20 U23447 (.o(n21745),
	.a(FE_RN_28),
	.b(FE_OCPN25932_n19501));
   no04f20 U23449 (.o(n19379),
	.a(n18148),
	.b(n19377),
	.c(n19376),
	.d(n18147));
   in01f10 U23450 (.o(n18147),
	.a(n19374));
   no04f40 U23451 (.o(n22889),
	.a(n18150),
	.b(n19341),
	.c(n19340),
	.d(n18149));
   ao12f08 U23452 (.o(n19295),
	.a(n19282),
	.b(n19825),
	.c(n19283));
   ao22f10 U23453 (.o(n18917),
	.a(myChipID_f_12_),
	.b(FE_OCPN25904_n18927),
	.c(n19617),
	.d(n23508));
   na02f20 U23454 (.o(n18151),
	.a(FE_OCPN25966_proc_input_NIB_head_ptr_f_2),
	.b(proc_input_NIB_head_ptr_f_3_));
   na02f08 U23455 (.o(n18157),
	.a(n18159),
	.b(n18158));
   ao22f06 U23456 (.o(n18159),
	.a(proc_input_NIB_storage_data_f_11__56_),
	.b(FE_OCPN25921_n19547),
	.c(proc_input_NIB_storage_data_f_9__56_),
	.d(FE_OFN25681_n17814));
   ao22f06 U23457 (.o(n18163),
	.a(proc_input_NIB_storage_data_f_3__56_),
	.b(FE_RN_33),
	.c(proc_input_NIB_storage_data_f_0__56_),
	.d(FE_OCPN25839_n24342));
   in01f04 U23458 (.o(n18170),
	.a(n19085));
   no02f20 U23459 (.o(n26025),
	.a(n23400),
	.b(n19026));
   no03f20 U23460 (.o(n18902),
	.a(n18181),
	.b(n18176),
	.c(n18172));
   oa22f10 U23461 (.o(n18172),
	.a(n19622),
	.b(n25516),
	.c(n19575),
	.d(n23587));
   na03f20 U23462 (.o(n23587),
	.a(n18175),
	.b(n18174),
	.c(n18173));
   na02f10 U23463 (.o(n18179),
	.a(FE_RN_5),
	.b(west_input_NIB_storage_data_f_3__59_));
   ao22f20 U23464 (.o(n18180),
	.a(n18828),
	.b(west_input_NIB_storage_data_f_1__59_),
	.c(FE_RN_66),
	.d(west_input_NIB_storage_data_f_0__59_));
   no02f20 U23465 (.o(n18181),
	.a(n19633),
	.b(n23317));
   na03f20 U23466 (.o(n23317),
	.a(n18184),
	.b(n18183),
	.c(n18182));
   na02f08 U23467 (.o(n18182),
	.a(west_input_NIB_storage_data_f_3__55_),
	.b(FE_RN_5));
   no03f04 U23468 (.o(n20348),
	.a(n18624),
	.b(n18623),
	.c(n20341));
   no03f06 U23469 (.o(n18279),
	.a(n18283),
	.b(n18280),
	.c(n20468));
   no02f20 U23470 (.o(n19508),
	.a(n19507),
	.b(n19506));
   ao12f02 U23471 (.o(n19566),
	.a(n20199),
	.b(n19565),
	.c(n19564));
   oa12f02 U23472 (.o(n20195),
	.a(n20193),
	.b(n20194),
	.c(n20231));
   oa22f02 U23473 (.o(north_output_control_N468),
	.a(n25130),
	.b(n25137),
	.c(n18279),
	.d(n18277));
   no02f01 U23474 (.o(north_output_control_N72),
	.a(FE_RN_67),
	.b(n18594));
   no02f08 U23475 (.o(n26024),
	.a(FE_RN_67),
	.b(n19471));
   na02f08 U23476 (.o(n18219),
	.a(n18273),
	.b(n20475));
   ao12f10 U23477 (.o(n18221),
	.a(n25087),
	.b(FE_RN_2),
	.c(n18273));
   ao22f08 U23478 (.o(n18229),
	.a(proc_input_NIB_storage_data_f_3__62_),
	.b(n17754),
	.c(proc_input_NIB_storage_data_f_8__62_),
	.d(FE_OFN25645_n21748));
   no02f10 U23479 (.o(n18234),
	.a(n18236),
	.b(n18235));
   no02f10 U23480 (.o(n18237),
	.a(n18239),
	.b(n18238));
   na02f08 U23481 (.o(n18238),
	.a(n18417),
	.b(n18420));
   na02f10 U23482 (.o(n18248),
	.a(n18242),
	.b(n18241));
   na02f10 U23483 (.o(n18241),
	.a(n19622),
	.b(n25518));
   na03f20 U23484 (.o(n25518),
	.a(n18254),
	.b(n18255),
	.c(n18253));
   no02f10 U23485 (.o(n18242),
	.a(n18244),
	.b(n18243));
   no02f08 U23486 (.o(n18243),
	.a(myChipID_f_1_),
	.b(n19151));
   no02f10 U23487 (.o(n18244),
	.a(myChipID_f_1_),
	.b(n19152));
   no03f20 U23488 (.o(n18304),
	.a(n18249),
	.b(n18248),
	.c(n18245));
   na04f10 U23489 (.o(n18246),
	.a(n18253),
	.b(n18255),
	.c(n18254),
	.d(myChipID_f_9_));
   na03f10 U23490 (.o(n18247),
	.a(n19151),
	.b(n19152),
	.c(myChipID_f_1_));
   no02f10 U23491 (.o(n18249),
	.a(n18251),
	.b(n18250));
   in01f08 U23492 (.o(n18250),
	.a(n18252));
   na02f10 U23493 (.o(n18254),
	.a(FE_OFN25610_n19071),
	.b(north_input_NIB_storage_data_f_1__59_));
   no02f20 U23494 (.o(n21485),
	.a(n18272),
	.b(n18271));
   in01f10 U23495 (.o(n18271),
	.a(n19186));
   in01f10 U23496 (.o(n18272),
	.a(n19185));
   no02f04 U23497 (.o(n18293),
	.a(n25091),
	.b(n19059));
   na03f20 U23498 (.o(n19203),
	.a(n18304),
	.b(n18302),
	.c(n18299));
   no02f10 U23499 (.o(n18299),
	.a(n18301),
	.b(n18300));
   oa22f10 U23500 (.o(n18300),
	.a(n18461),
	.b(n18460),
	.c(myChipID_f_3_),
	.d(n19150));
   oa22f08 U23501 (.o(n18301),
	.a(n19666),
	.b(n23331),
	.c(myChipID_f_0_),
	.d(n19165));
   ao12f10 U23502 (.o(n18302),
	.a(n18303),
	.b(n19575),
	.c(n18459));
   no02f10 U23503 (.o(n18303),
	.a(n19657),
	.b(n23342));
   na02f40 U23504 (.o(n20109),
	.a(n20343),
	.b(n18305));
   na02f40 U23505 (.o(n18305),
	.a(n20403),
	.b(n19248));
   na03f20 U23506 (.o(n23333),
	.a(n18311),
	.b(n18309),
	.c(n18306));
   no02f10 U23507 (.o(n18306),
	.a(n18308),
	.b(n18307));
   no02f20 U23508 (.o(n18309),
	.a(n18094),
	.b(n18310));
   no02f20 U23509 (.o(n18311),
	.a(n18313),
	.b(n18312));
   in01f08 U23510 (.o(n18313),
	.a(n19665));
   na02f04 U23511 (.o(n18314),
	.a(proc_input_NIB_storage_data_f_3__41_),
	.b(n19709));
   na03f20 U23512 (.o(n20286),
	.a(n20279),
	.b(n20284),
	.c(n18324));
   no02f10 U23513 (.o(n18324),
	.a(n18325),
	.b(n20278));
   no02f10 U23514 (.o(n18325),
	.a(myLocX_f_0_),
	.b(n20926));
   na02f20 U23515 (.o(n19830),
	.a(n20274),
	.b(n20282));
   no02f10 U23516 (.o(n20282),
	.a(n20273),
	.b(n18328));
   no02f10 U23517 (.o(n20274),
	.a(n20277),
	.b(n18777));
   no02f10 U23518 (.o(n20277),
	.a(myLocX_f_7_),
	.b(n22822));
   ao22f10 U23519 (.o(n18674),
	.a(n24473),
	.b(south_input_NIB_storage_data_f_3__51_),
	.c(south_input_NIB_storage_data_f_0__51_),
	.d(FE_RN_62));
   na02f10 U23520 (.o(n18587),
	.a(south_input_NIB_storage_data_f_0__60_),
	.b(FE_OFN24744_n18648));
   ao22f20 U23521 (.o(n18653),
	.a(n24473),
	.b(south_input_NIB_storage_data_f_3__59_),
	.c(south_input_NIB_storage_data_f_0__59_),
	.d(FE_RN_62));
   no02f10 U23522 (.o(n18343),
	.a(n18344),
	.b(FE_OFN24745_n18648));
   ao22f20 U23523 (.o(n18662),
	.a(n24473),
	.b(south_input_NIB_storage_data_f_3__61_),
	.c(south_input_NIB_storage_data_f_0__61_),
	.d(FE_RN_62));
   in01f10 U23524 (.o(n18583),
	.a(n18333));
   ao12f08 U23525 (.o(n18710),
	.a(n18343),
	.b(FE_OCPN25945_n24965),
	.c(south_input_NIB_storage_data_f_3__38_));
   no02f10 U23526 (.o(n20467),
	.a(n20271),
	.b(n19832));
   na02f08 U23527 (.o(n20372),
	.a(n18095),
	.b(n20217));
   na02f10 U23528 (.o(n23496),
	.a(n18367),
	.b(n18358));
   na02f04 U23529 (.o(n18364),
	.a(n18366),
	.b(n18365));
   in01f08 U23530 (.o(n18381),
	.a(n20362));
   in01f08 U23531 (.o(n18382),
	.a(n20361));
   na02f40 U23532 (.o(n19550),
	.a(n18145),
	.b(n18385));
   no04f10 U23534 (.o(n22850),
	.a(n18390),
	.b(n18388),
	.c(n18387),
	.d(n18389));
   no04f08 U23535 (.o(n18628),
	.a(n18390),
	.b(n18388),
	.c(n18387),
	.d(n18386));
   na03f10 U23536 (.o(n18387),
	.a(n19710),
	.b(n19713),
	.c(n19714));
   na02f08 U23537 (.o(n19474),
	.a(n20252),
	.b(n20147));
   no02f10 U23538 (.o(n19475),
	.a(n19295),
	.b(n20251));
   na02f10 U23540 (.o(n18394),
	.a(n18395),
	.b(n18396));
   ao12f10 U23541 (.o(n18396),
	.a(west_output_control_planned_f),
	.b(n19475),
	.c(n20377));
   oa12f10 U23542 (.o(n20512),
	.a(n19480),
	.b(FE_RN_6),
	.c(n17774));
   na02f04 U23543 (.o(n19487),
	.a(n19486),
	.b(n18399));
   na02f04 U23544 (.o(n19485),
	.a(n25347),
	.b(n18399));
   na02f10 U23545 (.o(n18614),
	.a(n25433),
	.b(n18399));
   no02f10 U23546 (.o(n22943),
	.a(n18411),
	.b(n18814));
   no03f20 U23547 (.o(n19027),
	.a(n19830),
	.b(n20286),
	.c(n18778));
   ao22f04 U23548 (.o(n18420),
	.a(proc_input_NIB_storage_data_f_9__57_),
	.b(FE_OFN25682_n17814),
	.c(proc_input_NIB_storage_data_f_13__57_),
	.d(FE_OFN25602_n19530));
   na02f10 U23549 (.o(n19738),
	.a(n22842),
	.b(myLocY_f_1_));
   no02f04 U23550 (.o(n18423),
	.a(FE_RN_34),
	.b(n18424));
   no02f10 U23551 (.o(n25170),
	.a(n20452),
	.b(n20451));
   na02f10 U23552 (.o(n20215),
	.a(n20364),
	.b(n19737));
   na02f10 U23553 (.o(n19742),
	.a(n18467),
	.b(n19564));
   no02f10 U23554 (.o(n18435),
	.a(n20199),
	.b(n18436));
   na02f10 U23555 (.o(n20199),
	.a(n19562),
	.b(n19563));
   in01f08 U23556 (.o(n19733),
	.a(n23504));
   na02f10 U23559 (.o(n19668),
	.a(n18463),
	.b(n18462));
   na02f10 U23560 (.o(n18462),
	.a(n19666),
	.b(n23333));
   no02f10 U23561 (.o(n18467),
	.a(n20201),
	.b(n18468));
   no02f10 U23562 (.o(n22834),
	.a(n19560),
	.b(n19559));
   no02f10 U23563 (.o(n20201),
	.a(myLocY_f_1_),
	.b(n22842));
   no03f20 U23564 (.o(n22842),
	.a(n18487),
	.b(n18480),
	.c(n18484));
   na02f04 U23565 (.o(n18472),
	.a(n19872),
	.b(n20443));
   no02f06 U23566 (.o(n20448),
	.a(n20437),
	.b(n19871));
   in01m04 U23567 (.o(n18481),
	.a(n18565));
   na04f20 U23568 (.o(n18487),
	.a(n18491),
	.b(n18490),
	.c(n18489),
	.d(n18488));
   no02f20 U23569 (.o(validOut_P),
	.a(n25019),
	.b(n22943));
   na02f04 U23570 (.o(n18512),
	.a(proc_input_NIB_storage_data_f_4__45_),
	.b(n17742));
   na02f08 U23571 (.o(n18518),
	.a(n18520),
	.b(n18519));
   no02f20 U23573 (.o(n19655),
	.a(n25072),
	.b(FE_OCPN25931_n19501));
   na02f02 U23574 (.o(n25989),
	.a(n25236),
	.b(n18541));
   na02m02 U23575 (.o(n18542),
	.a(n18814),
	.b(n18543));
   no02f20 U23576 (.o(n18544),
	.a(n25986),
	.b(n25992));
   no02f20 U23577 (.o(n25986),
	.a(n25029),
	.b(n17759));
   no02f02 U23578 (.o(n18577),
	.a(n25147),
	.b(n18578));
   na02f01 U23579 (.o(n18578),
	.a(east_input_NIB_head_ptr_f_1_),
	.b(FE_OFN25596_reset));
   no02f10 U23580 (.o(n18651),
	.a(n18586),
	.b(n18579));
   na03f10 U23581 (.o(n21407),
	.a(n18582),
	.b(n18581),
	.c(n18580));
   na02f20 U23582 (.o(n18580),
	.a(south_input_NIB_storage_data_f_2__62_),
	.b(FE_RN_17));
   na03f40 U23583 (.o(n23995),
	.a(n18585),
	.b(n18584),
	.c(n18583));
   na02f10 U23584 (.o(n18584),
	.a(south_input_NIB_storage_data_f_2__54_),
	.b(n21806));
   na03f20 U23585 (.o(n20745),
	.a(n18589),
	.b(n18588),
	.c(n18587));
   na02f10 U23586 (.o(n18588),
	.a(south_input_NIB_storage_data_f_2__60_),
	.b(n21806));
   ao22f20 U23587 (.o(n18589),
	.a(south_input_NIB_storage_data_f_1__60_),
	.b(n17756),
	.c(n24473),
	.d(south_input_NIB_storage_data_f_3__60_));
   no02f20 U23588 (.o(n18714),
	.a(south_input_NIB_head_ptr_f_0_),
	.b(FE_RN_30));
   ao22f20 U23591 (.o(n18684),
	.a(n18061),
	.b(south_input_NIB_storage_data_f_1__52_),
	.c(south_input_NIB_storage_data_f_2__52_),
	.d(n21315));
   ao12f02 U23592 (.o(n19963),
	.a(n18602),
	.b(FE_OFN24741_n18683),
	.c(south_input_NIB_storage_data_f_1__29_));
   in01f08 U23593 (.o(n26027),
	.a(n18614));
   na03f20 U23594 (.o(n18733),
	.a(n18619),
	.b(n18618),
	.c(n18617));
   na02f20 U23595 (.o(n18618),
	.a(south_input_NIB_storage_data_f_2__39_),
	.b(n17782));
   no03f20 U23596 (.o(n23186),
	.a(n18729),
	.b(n18620),
	.c(n18728));
   no03f06 U23597 (.o(n18623),
	.a(FE_RN_26),
	.b(n24981),
	.c(FE_RN_18_0));
   no02f08 U23598 (.o(n18629),
	.a(n19708),
	.b(n23496));
   no02f10 U23599 (.o(n19722),
	.a(n19701),
	.b(n23326));
   no02f10 U23600 (.o(n20364),
	.a(n18630),
	.b(n20216));
   no02f10 U23601 (.o(n20216),
	.a(myLocX_f_2_),
	.b(n19733));
   no02f10 U23602 (.o(n18630),
	.a(myLocX_f_1_),
	.b(n19732));
   no02f10 U23603 (.o(n19737),
	.a(n20368),
	.b(n19735));
   na02f20 U23604 (.o(n18683),
	.a(FE_RN_42),
	.b(south_input_NIB_head_ptr_f_0_));
   in01f06 U23605 (.o(n25987),
	.a(n18642));
   na02f10 U23606 (.o(n20410),
	.a(n20294),
	.b(n20178));
   no03f02 U23607 (.o(south_output_control_N470),
	.a(reset),
	.b(n20348),
	.c(n20347));
   ao22f02 U23609 (.o(n2443),
	.a(n25325),
	.b(n25324),
	.c(n25323),
	.d(n25322));
   no02f02 U23610 (.o(n2863),
	.a(n25074),
	.b(n25073));
   na03f03 U23611 (.o(n25069),
	.a(n25067),
	.b(n25066),
	.c(n25065));
   na02f04 U23613 (.o(n2873),
	.a(n20510),
	.b(n20509));
   ao12f02 U23614 (.o(n25113),
	.a(n25111),
	.b(n25974),
	.c(thanksIn_P));
   no03f06 U23615 (.o(n25181),
	.a(n25180),
	.b(n25179),
	.c(n25178));
   oa22f02 U23616 (.o(n26000),
	.a(n20329),
	.b(n20328),
	.c(n25384),
	.d(n20327));
   no02f04 U23617 (.o(n20329),
	.a(n20317),
	.b(n20316));
   na02f02 U23618 (.o(n20460),
	.a(n20539),
	.b(n20457));
   oa22f02 U23619 (.o(n2563),
	.a(north_input_NIB_head_ptr_f_0_),
	.b(n25110),
	.c(n25429),
	.d(n25109));
   ao12f02 U23620 (.o(n24987),
	.a(n17758),
	.b(n24976),
	.c(n24975));
   na02f04 U23621 (.o(n24975),
	.a(n24973),
	.b(n24972));
   na03f02 U23622 (.o(n26003),
	.a(n20562),
	.b(n20561),
	.c(n20560));
   ao12f02 U23623 (.o(west_output_control_N470),
	.a(n20459),
	.b(n20461),
	.c(n20460));
   oa12f04 U23624 (.o(n20459),
	.a(FE_OFN575_n25463),
	.b(n20537),
	.c(n20458));
   ao12f02 U23626 (.o(n2578),
	.a(n25277),
	.b(n25432),
	.c(n25278));
   no03f02 U23627 (.o(west_output_control_N467),
	.a(FE_OFN5_reset),
	.b(n25187),
	.c(n25186));
   ao12f02 U23628 (.o(east_output_control_N469),
	.a(n25068),
	.b(n25384),
	.c(n25069));
   ao12f02 U23629 (.o(west_output_control_N468),
	.a(n20542),
	.b(n20544),
	.c(n20543));
   oa12f04 U23630 (.o(n20542),
	.a(FE_OFN575_n25463),
	.b(n20541),
	.c(n20540));
   oa12f02 U23632 (.o(n20536),
	.a(n21695),
	.b(n20535),
	.c(n25174));
   oa22f02 U23633 (.o(n2833),
	.a(n25490),
	.b(n25489),
	.c(n25488),
	.d(n25487));
   in01f02 U23634 (.o(n25110),
	.a(n26010));
   oa12f02 U23635 (.o(n2423),
	.a(n25146),
	.b(n25148),
	.c(n25147));
   no02f02 U23636 (.o(n2433),
	.a(n25342),
	.b(n25341));
   in01f02 U23637 (.o(n20124),
	.a(n20113));
   oa22f02 U23638 (.o(n20453),
	.a(FE_OFN526_n24731),
	.b(n25169),
	.c(n17786),
	.d(n25170));
   no04f20 U23639 (.o(n19146),
	.a(n19131),
	.b(n20175),
	.c(n19144),
	.d(n19130));
   ao12f02 U23640 (.o(n19888),
	.a(n19887),
	.b(n24976),
	.c(n24982));
   no03f06 U23641 (.o(n20373),
	.a(n20368),
	.b(n20367),
	.c(n20366));
   na03f03 U23643 (.o(n25313),
	.a(n25312),
	.b(n25311),
	.c(n25310));
   oa22f02 U23644 (.o(n2558),
	.a(n25432),
	.b(n25431),
	.c(n25430),
	.d(n25429));
   na02m02 U23645 (.o(n25119),
	.a(n25115),
	.b(n25114));
   ao22f02 U23646 (.o(east_output_control_N468),
	.a(n25403),
	.b(n25402),
	.c(n25401),
	.d(n25400));
   ao12f02 U23647 (.o(proc_output_control_N470),
	.a(FE_OFN5_reset),
	.b(n25314),
	.c(n25313));
   na02f02 U23648 (.o(n25991),
	.a(n25272),
	.b(n25271));
   na02f04 U23649 (.o(n25271),
	.a(n25270),
	.b(n26027));
   na02f04 U23650 (.o(n25349),
	.a(n26027),
	.b(n25348));
   na02f02 U23651 (.o(n25990),
	.a(n25350),
	.b(n25349));
   in01f10 U23652 (.o(n18668),
	.a(n18664));
   no03f40 U23653 (.o(n20437),
	.a(n18947),
	.b(n18946),
	.c(n18945));
   na02s01 U23654 (.o(n25126),
	.a(FE_OFN428_n22902),
	.b(FE_OFN25975_n21666));
   in01f01 U23655 (.o(n25097),
	.a(n25126));
   ao12f02 U23658 (.o(n20396),
	.a(n20392),
	.b(n20394),
	.c(n20393));
   no03f01 U23659 (.o(n25720),
	.a(ec_thanks_n_to_p_reg),
	.b(ec_thanks_p_to_p_reg),
	.c(ec_thanks_s_to_p_reg));
   in01s01 U23660 (.o(n25721),
	.a(n25720));
   no02f02 U23661 (.o(n20193),
	.a(n20192),
	.b(n20191));
   no02s01 U23662 (.o(n25784),
	.a(n25783),
	.b(n25785));
   ao22s01 U23663 (.o(n25725),
	.a(n25724),
	.b(ec_cfg_0_),
	.c(n25723),
	.d(n25722));
   no04f20 U23664 (.o(n20175),
	.a(n20155),
	.b(n19126),
	.c(n20154),
	.d(n19125));
   in01s01 U23665 (.o(n25756),
	.a(ec_south_input_valid_reg));
   ao22f04 U23666 (.o(n19097),
	.a(FE_RN_11),
	.b(north_input_NIB_storage_data_f_2__37_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__37_));
   in01s01 U23668 (.o(n25727),
	.a(n25726));
   in01s01 U23669 (.o(n25765),
	.a(n25764));
   no02f08 U23670 (.o(n18963),
	.a(n19871),
	.b(n20263));
   na02f02 U23671 (.o(n24664),
	.a(n24100),
	.b(n24099));
   na02f02 U23672 (.o(n24703),
	.a(n24075),
	.b(n24074));
   na02f02 U23673 (.o(n23560),
	.a(n21828),
	.b(n21827));
   na02f03 U23674 (.o(n23579),
	.a(n21786),
	.b(n21785));
   na02f02 U23675 (.o(n24601),
	.a(n24282),
	.b(n24281));
   na02f02 U23676 (.o(n24631),
	.a(n24475),
	.b(n24474));
   na02f04 U23677 (.o(n24741),
	.a(n24212),
	.b(n24211));
   na02f02 U23679 (.o(n24019),
	.a(n21860),
	.b(n21859));
   in01f03 U23680 (.o(n18833),
	.a(n18832));
   in01f01 U23681 (.o(n23630),
	.a(n18910));
   in01s01 U23682 (.o(n25436),
	.a(west_output_space_yummy_f));
   in01s01 U23684 (.o(n20768),
	.a(n21156));
   no03f20 U23685 (.o(n19244),
	.a(n19147),
	.b(n19146),
	.c(n19145));
   in01s01 U23686 (.o(n20648),
	.a(north_input_control_thanks_all_f));
   na04f04 U23687 (.o(n25388),
	.a(n19022),
	.b(n25387),
	.c(FE_OFN25598_reset),
	.d(n25392));
   in01s01 U23688 (.o(n20726),
	.a(west_input_control_count_f_4_));
   in01s01 U23689 (.o(n22388),
	.a(east_output_space_count_f_0_));
   no02s01 U23690 (.o(n21650),
	.a(proc_input_control_count_f_5_),
	.b(proc_input_control_count_f_6_));
   ao22f04 U23691 (.o(n19060),
	.a(n19054),
	.b(east_input_valid),
	.c(n19056),
	.d(north_input_valid));
   in01s01 U23692 (.o(n22066),
	.a(n22076));
   in01s01 U23693 (.o(n25729),
	.a(ec_cfg_2_));
   in01s01 U23694 (.o(n25714),
	.a(ec_thanks_s_to_p_reg));
   no02s01 U23695 (.o(n25753),
	.a(ec_cfg_6_),
	.b(ec_wants_to_send_but_cannot_S));
   no02s01 U23696 (.o(n25806),
	.a(ec_cfg_12_),
	.b(n25808));
   ao22f01 U23697 (.o(n22363),
	.a(FE_OFN94_n21695),
	.b(n23976),
	.c(n17755),
	.d(n23977));
   ao22f01 U23698 (.o(n24521),
	.a(FE_OFN105_n22517),
	.b(n24703),
	.c(FE_OFN93_n21667),
	.d(FE_OFN515_n24702));
   ao12f04 U23699 (.o(n25182),
	.a(n25172),
	.b(n25174),
	.c(n25173));
   no02f04 U23700 (.o(n20122),
	.a(reset),
	.b(n20121));
   na02f02 U23701 (.o(n19936),
	.a(n19935),
	.b(n19934));
   in01s01 U23702 (.o(n20736),
	.a(n20735));
   in01s01 U23703 (.o(n22381),
	.a(n22377));
   na02s01 U23704 (.o(n25467),
	.a(n25466),
	.b(n25465));
   no02f01 U23705 (.o(n25731),
	.a(n25730),
	.b(n25729));
   ao22s01 U23706 (.o(n25750),
	.a(ec_cfg_4_),
	.b(n25742),
	.c(n25741),
	.d(n25746));
   ao22s01 U23707 (.o(n25812),
	.a(ec_cfg_13_),
	.b(n25803),
	.c(n25802),
	.d(n25808));
   na02f02 U23708 (.o(n24582),
	.a(n24581),
	.b(n24580));
   na02f02 U23709 (.o(n23954),
	.a(n23953),
	.b(n23952));
   na02f02 U23710 (.o(n23635),
	.a(n23634),
	.b(n23633));
   na02f02 U23711 (.o(n22345),
	.a(n22344),
	.b(n22343));
   oa22f01 U23712 (.o(n21546),
	.a(FE_OFN483_n23987),
	.b(n22772),
	.c(n23986),
	.d(n22773));
   na02f02 U23713 (.o(n22235),
	.a(n22234),
	.b(n22233));
   na02f02 U23714 (.o(n22600),
	.a(n22599),
	.b(n22598));
   na02f02 U23715 (.o(n24534),
	.a(n24533),
	.b(n24532));
   na02f02 U23716 (.o(n21374),
	.a(n21373),
	.b(n21372));
   na02f01 U23717 (.o(n24332),
	.a(n24331),
	.b(n24330));
   na02f02 U23719 (.o(n20963),
	.a(n20962),
	.b(n20961));
   in01s01 U23721 (.o(n21589),
	.a(n24030));
   ao22f02 U23722 (.o(n25342),
	.a(n25330),
	.b(n25329),
	.c(n25340),
	.d(FE_OFN25596_reset));
   in01s01 U23723 (.o(n20483),
	.a(n20481));
   na02s01 U23724 (.o(n20711),
	.a(n25433),
	.b(n20737));
   na02s01 U23725 (.o(n22911),
	.a(n23550),
	.b(n22495));
   na02s01 U23727 (.o(n23828),
	.a(proc_input_NIB_storage_data_f_0__61_),
	.b(FE_OFN25618_n23789));
   na02f01 U23728 (.o(n23891),
	.a(proc_input_NIB_storage_data_f_0__46_),
	.b(n25547));
   na02f01 U23729 (.o(n23790),
	.a(proc_input_NIB_storage_data_f_0__31_),
	.b(FE_OFN25622_n23789));
   oa22f01 U23730 (.o(n25529),
	.a(FE_OFN25620_n23789),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_0__18_),
	.d(FE_OFN580_n25547));
   oa22s01 U23731 (.o(n25544),
	.a(FE_OFN25621_n23789),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_0__3_),
	.d(FE_OFN580_n25547));
   na02s01 U23732 (.o(n23831),
	.a(proc_input_NIB_storage_data_f_1__52_),
	.b(FE_OFN374_n17762));
   na02f01 U23733 (.o(n23775),
	.a(proc_input_NIB_storage_data_f_1__37_),
	.b(FE_OFN373_n17762));
   na02f01 U23734 (.o(n23763),
	.a(proc_input_NIB_storage_data_f_1__23_),
	.b(FE_OFN373_n17762));
   oa22f01 U23735 (.o(n25562),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_1__9_),
	.d(n25571));
   na02s01 U23736 (.o(n23899),
	.a(proc_input_NIB_storage_data_f_2__58_),
	.b(FE_OFN272_n25595));
   na02s01 U23737 (.o(n23774),
	.a(proc_input_NIB_storage_data_f_2__43_),
	.b(n17764));
   na02s01 U23738 (.o(n23758),
	.a(proc_input_NIB_storage_data_f_2__28_),
	.b(n17764));
   oa22f01 U23739 (.o(n25580),
	.a(n17764),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_2__15_),
	.d(n25595));
   oa22f01 U23740 (.o(n25596),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_2__0_),
	.d(n25595));
   na02s01 U23741 (.o(n23867),
	.a(proc_input_NIB_storage_data_f_3__49_),
	.b(FE_OFN25778_FE_OFN582_n25619));
   na02s01 U23742 (.o(n23748),
	.a(proc_input_NIB_storage_data_f_3__34_),
	.b(FE_OFN25777_FE_OFN582_n25619));
   oa22s01 U23743 (.o(n25598),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_3__21_),
	.d(n25619));
   oa22s01 U23744 (.o(n25613),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_3__6_),
	.d(n25619));
   na02s01 U23745 (.o(n23723),
	.a(proc_input_NIB_storage_data_f_4__55_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02s01 U23746 (.o(n23165),
	.a(proc_input_NIB_storage_data_f_4__41_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02f02 U23747 (.o(n23638),
	.a(proc_input_NIB_storage_data_f_4__26_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   oa22m01 U23748 (.o(n23123),
	.a(FE_OFN25761_FE_OFN1077_n17766),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_4__13_),
	.d(n23090));
   na02s01 U23749 (.o(n23648),
	.a(proc_input_NIB_storage_data_f_5__62_),
	.b(FE_OFN368_n17761));
   na02s01 U23750 (.o(n23167),
	.a(proc_input_NIB_storage_data_f_5__47_),
	.b(FE_OFN369_n17761));
   oa22m01 U23751 (.o(n23133),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_5__33_),
	.d(n23102));
   oa22m01 U23752 (.o(n23131),
	.a(FE_OFN368_n17761),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_5__20_),
	.d(n23102));
   oa22m01 U23753 (.o(n23109),
	.a(FE_OFN369_n17761),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_5__5_),
	.d(n23102));
   na02s01 U23754 (.o(n23362),
	.a(proc_input_NIB_storage_data_f_6__40_),
	.b(FE_OFN25798_n23051));
   na02s01 U23755 (.o(n23707),
	.a(proc_input_NIB_storage_data_f_6__25_),
	.b(FE_OFN25801_n23051));
   oa22f01 U23756 (.o(n23065),
	.a(n23051),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_6__12_),
	.d(FE_OFN440_n23051));
   na02s01 U23757 (.o(n23709),
	.a(proc_input_NIB_storage_data_f_7__61_),
	.b(n17767));
   na02s01 U23758 (.o(n23728),
	.a(proc_input_NIB_storage_data_f_7__46_),
	.b(n17767));
   oa22s01 U23759 (.o(n23079),
	.a(FE_OFN1081_n17767),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_7__18_),
	.d(n23046));
   oa22s01 U23760 (.o(n23062),
	.a(n17767),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_7__3_),
	.d(n23046));
   na02s01 U23761 (.o(n23380),
	.a(proc_input_NIB_storage_data_f_11__52_),
	.b(FE_OFN1085_n22923));
   na02s01 U23762 (.o(n22921),
	.a(proc_input_NIB_storage_data_f_11__38_),
	.b(FE_OFN1086_n22923));
   na02s01 U23763 (.o(n23384),
	.a(proc_input_NIB_storage_data_f_11__23_),
	.b(FE_OFN1086_n22923));
   oa22s01 U23764 (.o(n22784),
	.a(FE_OFN1085_n22923),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_11__10_),
	.d(n22779));
   na02s01 U23765 (.o(n23284),
	.a(proc_input_NIB_storage_data_f_15__61_),
	.b(n17768));
   na02s01 U23766 (.o(n23270),
	.a(proc_input_NIB_storage_data_f_15__46_),
	.b(n17768));
   oa22s01 U23767 (.o(n25631),
	.a(FE_OFN585_n25643),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_15__12_),
	.d(n25643));
   ao12s01 U23768 (.o(n25981),
	.a(proc_input_NIB_tail_ptr_f_2_),
	.b(n25980),
	.c(n25979));
   na02s01 U23769 (.o(n22561),
	.a(west_input_NIB_storage_data_f_0__25_),
	.b(FE_OFN24796_n20854));
   in01s01 U23770 (.o(n25966),
	.a(west_input_NIB_storage_data_f_0__11_));
   na02f01 U23771 (.o(n22585),
	.a(west_input_NIB_storage_data_f_1__32_),
	.b(FE_OFN381_n17772));
   in01s01 U23772 (.o(n25954),
	.a(west_input_NIB_storage_data_f_1__17_));
   oa22s01 U23773 (.o(n22266),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_3_),
	.c(west_input_NIB_storage_data_f_1__3_),
	.d(FE_OFN380_n17772));
   in01s01 U23774 (.o(n25943),
	.a(west_input_NIB_storage_data_f_2__9_));
   in01s01 U23775 (.o(n21093),
	.a(dataIn_W_62_));
   in01s01 U23776 (.o(n21125),
	.a(dataIn_W_47_));
   in01s01 U23777 (.o(n22736),
	.a(dataIn_W_24_));
   na02s01 U23778 (.o(n20829),
	.a(south_input_NIB_storage_data_f_0__29_),
	.b(FE_OFN952_n25916));
   oa22s01 U23779 (.o(n24800),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_14_),
	.c(south_input_NIB_storage_data_f_0__14_),
	.d(FE_OFN83_n20814));
   oa22s01 U23780 (.o(n22254),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_2_),
	.c(south_input_NIB_storage_data_f_0__2_),
	.d(FE_OFN83_n20814));
   oa22f01 U23781 (.o(n24815),
	.a(FE_OFN25787_n17770),
	.b(dataIn_S_21_),
	.c(south_input_NIB_storage_data_f_1__21_),
	.d(n20797));
   in01s01 U23782 (.o(n20998),
	.a(dataIn_S_49_));
   in01s01 U23783 (.o(n22667),
	.a(dataIn_S_34_));
   na02s01 U23784 (.o(n21031),
	.a(south_input_NIB_storage_data_f_3__26_),
	.b(n17769));
   oa22s01 U23785 (.o(n24842),
	.a(n17769),
	.b(dataIn_S_17_),
	.c(south_input_NIB_storage_data_f_3__17_),
	.d(n20996));
   in01s01 U23786 (.o(n25893),
	.a(east_input_NIB_storage_data_f_0__16_));
   in01s01 U23787 (.o(n24771),
	.a(east_input_NIB_storage_data_f_1__58_));
   na02s01 U23788 (.o(n24790),
	.a(dataIn_E_50_),
	.b(FE_OFN555_n24761));
   na02s01 U23789 (.o(n24898),
	.a(dataIn_E_35_),
	.b(n24761));
   na02s01 U23790 (.o(n24882),
	.a(dataIn_E_27_),
	.b(FE_OFN555_n24761));
   in01s01 U23791 (.o(n25879),
	.a(east_input_NIB_storage_data_f_1__5_));
   in01s01 U23792 (.o(n25196),
	.a(dataIn_E_55_));
   in01s01 U23793 (.o(n24931),
	.a(dataIn_E_40_));
   in01s01 U23794 (.o(n25222),
	.a(dataIn_E_32_));
   in01s01 U23795 (.o(n25865),
	.a(east_input_NIB_storage_data_f_3__3_));
   na02s01 U23796 (.o(n20953),
	.a(north_input_NIB_storage_data_f_0__62_),
	.b(n17771));
   na02s01 U23797 (.o(n20943),
	.a(north_input_NIB_storage_data_f_0__47_),
	.b(n20934));
   na02s01 U23798 (.o(n22639),
	.a(north_input_NIB_storage_data_f_0__32_),
	.b(n20934));
   oa22s01 U23799 (.o(n24834),
	.a(n20934),
	.b(dataIn_N_17_),
	.c(north_input_NIB_storage_data_f_0__17_),
	.d(FE_OFN1092_n20934));
   oa22s01 U23800 (.o(n22342),
	.a(n17771),
	.b(dataIn_N_5_),
	.c(north_input_NIB_storage_data_f_0__5_),
	.d(FE_OFN1092_n20934));
   in01s01 U23801 (.o(n22634),
	.a(dataIn_N_49_));
   in01s01 U23802 (.o(n22648),
	.a(dataIn_N_34_));
   in01s01 U23803 (.o(n21266),
	.a(dataIn_N_26_));
   in01s01 U23804 (.o(n25855),
	.a(dataIn_N_18_));
   in01s01 U23805 (.o(n25851),
	.a(dataIn_N_6_));
   in01s01 U23806 (.o(n20608),
	.a(myLocY_6_));
   in01s01 U23807 (.o(n20605),
	.a(myChipID_13_));
   ao12f01 U23808 (.o(n25733),
	.a(n25731),
	.b(ec_thanks_w_to_p_reg),
	.c(n25732));
   in01s01 U23810 (.o(n24026),
	.a(n24025));
   no02f01 U23813 (.o(n22532),
	.a(n22531),
	.b(n22530));
   no02m01 U23815 (.o(n22756),
	.a(n22755),
	.b(n22754));
   in01s01 U23816 (.o(n22613),
	.a(n22612));
   in01s01 U23817 (.o(n22438),
	.a(n22437));
   no02f02 U23818 (.o(n21605),
	.a(n21604),
	.b(n21603));
   no02f02 U23819 (.o(n21602),
	.a(n21601),
	.b(n21600));
   in01f01 U23820 (.o(n24371),
	.a(n24370));
   in01s01 U23821 (.o(n24415),
	.a(n24414));
   no02f01 U23822 (.o(n20915),
	.a(n20914),
	.b(n20913));
   no02f02 U23825 (.o(n21483),
	.a(n21482),
	.b(n21481));
   no02f01 U23826 (.o(n21144),
	.a(n21143),
	.b(n21142));
   oa12f02 U23828 (.o(n2573),
	.a(n25291),
	.b(n25293),
	.c(n25292));
   oa22f01 U23829 (.o(proc_input_control_N44),
	.a(FE_OFN127_n23536),
	.b(n21694),
	.c(n21645),
	.d(n21689));
   in01s01 U23830 (.o(n3343),
	.a(n25534));
   in01s01 U23831 (.o(n3643),
	.a(n25554));
   in01s01 U23832 (.o(n3718),
	.a(n25569));
   in01s01 U23833 (.o(n3943),
	.a(n25574));
   in01s01 U23834 (.o(n4018),
	.a(n25589));
   in01s01 U23835 (.o(n4318),
	.a(n25609));
   in01s01 U23836 (.o(n4618),
	.a(n23121));
   in01s01 U23837 (.o(n4843),
	.a(n23133));
   in01s01 U23838 (.o(n4918),
	.a(n23127));
   in01s01 U23839 (.o(n4993),
	.a(n23107));
   in01s01 U23840 (.o(n5293),
	.a(n23068));
   in01s01 U23841 (.o(n5593),
	.a(n23056));
   in01s01 U23842 (.o(n5893),
	.a(n23463));
   in01s01 U23843 (.o(n5968),
	.a(n23446));
   in01s01 U23844 (.o(n6193),
	.a(n23442));
   in01s01 U23845 (.o(n6268),
	.a(n23421));
   in01s01 U23846 (.o(n6568),
	.a(n23437));
   in01s01 U23847 (.o(n6868),
	.a(n22793));
   in01s01 U23848 (.o(n7168),
	.a(n23205));
   in01s01 U23849 (.o(n7243),
	.a(n23220));
   in01s01 U23850 (.o(n7468),
	.a(n23208));
   in01s01 U23851 (.o(n7543),
	.a(n23230));
   in01s01 U23852 (.o(n7843),
	.a(n23254));
   in01s01 U23853 (.o(n8143),
	.a(n25630));
   no02s01 U23854 (.o(n8218),
	.a(n25983),
	.b(n25981));
   oa12s01 U23855 (.o(n8293),
	.a(n20864),
	.b(FE_OFN25750_FE_OFN24796_n20854),
	.c(n21084));
   oa12f01 U23856 (.o(n8368),
	.a(n20878),
	.b(FE_OFN25751_FE_OFN24796_n20854),
	.c(n21117));
   in01s01 U23857 (.o(n8443),
	.a(n24809));
   in01s01 U23858 (.o(n8518),
	.a(n22260));
   oa12f01 U23859 (.o(n8593),
	.a(n22586),
	.b(FE_OFN381_n17772),
	.c(n22724));
   oa12f01 U23860 (.o(n8668),
	.a(n20906),
	.b(FE_OFN381_n17772),
	.c(n21109));
   oa12s01 U23861 (.o(n8743),
	.a(n20898),
	.b(FE_OFN381_n17772),
	.c(n22726));
   ao22s01 U23862 (.o(n8818),
	.a(FE_OFN380_n17772),
	.b(n25964),
	.c(n25952),
	.d(FE_OFN382_n17772));
   in01s01 U23863 (.o(n9118),
	.a(n24853));
   in01s01 U23864 (.o(n9343),
	.a(n24868));
   in01s01 U23865 (.o(n9418),
	.a(n24867));
   in01s01 U23866 (.o(n9493),
	.a(n22419));
   oa12s01 U23867 (.o(n9568),
	.a(n20843),
	.b(FE_OFN403_n20815),
	.c(n21040));
   oa12s01 U23868 (.o(n9643),
	.a(n22547),
	.b(FE_OFN952_n25916),
	.c(n22582));
   oa12s01 U23869 (.o(n9718),
	.a(n20823),
	.b(FE_OFN952_n25916),
	.c(n21044));
   in01s01 U23870 (.o(n9793),
	.a(n22255));
   oa12s01 U23871 (.o(n9868),
	.a(n20842),
	.b(FE_OFN25857_FE_OFN899_n17770),
	.c(n21022));
   oa12f01 U23872 (.o(n9943),
	.a(n22576),
	.b(FE_OFN25785_n17770),
	.c(n22692));
   oa12s01 U23873 (.o(n10018),
	.a(n20800),
	.b(FE_OFN25785_n17770),
	.c(n21030));
   in01s01 U23874 (.o(n10093),
	.a(n24813));
   in01s01 U23875 (.o(n10393),
	.a(n24836));
   in01s01 U23876 (.o(n10468),
	.a(n22397));
   oa12s01 U23877 (.o(n10543),
	.a(n22483),
	.b(n22484),
	.c(FE_OFN896_n17769));
   oa12s01 U23878 (.o(n10618),
	.a(n22669),
	.b(n22706),
	.c(n17769));
   in01s01 U23879 (.o(n10693),
	.a(n24847));
   in01s01 U23880 (.o(n10768),
	.a(n22403));
   in01s01 U23881 (.o(n11068),
	.a(n25653));
   in01s01 U23882 (.o(n11443),
	.a(n25678));
   in01s01 U23883 (.o(n11668),
	.a(n25681));
   in01s01 U23884 (.o(n12043),
	.a(n25707));
   oa12s01 U23885 (.o(n12118),
	.a(n20952),
	.b(n17771),
	.c(n21287));
   oa12s01 U23886 (.o(n12193),
	.a(n22631),
	.b(n20934),
	.c(n22632));
   oa12s01 U23887 (.o(n12268),
	.a(n20941),
	.b(n20934),
	.c(n21259));
   in01s01 U23888 (.o(n12343),
	.a(n24832));
   in01s01 U23889 (.o(n12418),
	.a(n22336));
   in01s01 U23890 (.o(n12718),
	.a(n22468));
   in01s01 U23891 (.o(n13018),
	.a(n22058));
   in01s01 U23892 (.o(n13318),
	.a(n22458));
   oa12f01 U23893 (.o(FE_OFN1066_dataOut_P_5),
	.a(n23981),
	.b(n23982),
	.c(FE_OFN524_n24728));
   oa12f02 U23894 (.o(dataOut_W_61_),
	.a(n22756),
	.b(n24009),
	.c(FE_OFN25878_n19446));
   oa12f01 U23895 (.o(FE_OFN25733_dataOut_E_8),
	.a(n21767),
	.b(n23154),
	.c(FE_OFN25895_n25395));
   no02f01 U23896 (.o(n18646),
	.a(proc_output_space_is_two_or_more_f),
	.b(proc_output_space_yummy_f));
   na02f80 U23897 (.o(n24965),
	.a(south_input_NIB_head_ptr_f_0_),
	.b(south_input_NIB_head_ptr_f_1_));
   no02f40 U23899 (.o(n18648),
	.a(south_input_NIB_head_ptr_f_1_),
	.b(south_input_NIB_head_ptr_f_0_));
   in01f10 U23903 (.o(n18701),
	.a(n18651));
   in01f40 U23904 (.o(n19973),
	.a(n18754));
   na02f10 U23905 (.o(n18654),
	.a(n18060),
	.b(south_input_NIB_storage_data_f_1__58_));
   oa22f10 U23906 (.o(n18657),
	.a(n24965),
	.b(n18656),
	.c(FE_OFN24745_n18648),
	.d(n18655));
   no03f20 U23907 (.o(n23590),
	.a(n18659),
	.b(n18658),
	.c(n18657));
   in01f10 U23908 (.o(n18660),
	.a(FE_RN_43));
   ao22f20 U23909 (.o(n18682),
	.a(n19622),
	.b(n18028),
	.c(n19575),
	.d(n18660));
   ao22f10 U23910 (.o(n18661),
	.a(n21806),
	.b(south_input_NIB_storage_data_f_2__61_),
	.c(FE_RN_55),
	.d(south_input_NIB_storage_data_f_1__61_));
   na02f20 U23911 (.o(n24004),
	.a(n18662),
	.b(n18661));
   oa22f10 U23912 (.o(n18667),
	.a(n24965),
	.b(n18666),
	.c(n24964),
	.d(n18665));
   no03f20 U23913 (.o(n21484),
	.a(n18669),
	.b(n18668),
	.c(n18667));
   in01f10 U23914 (.o(n18670),
	.a(n21484));
   ao22f20 U23915 (.o(n18681),
	.a(n19584),
	.b(n24004),
	.c(n19633),
	.d(n18670));
   na02f20 U23916 (.o(n23332),
	.a(n18672),
	.b(n18671));
   na02f20 U23917 (.o(n25510),
	.a(n18674),
	.b(n18673));
   ao22f20 U23918 (.o(n18680),
	.a(n19666),
	.b(n23332),
	.c(n19594),
	.d(n25510));
   ao22f20 U23919 (.o(n18676),
	.a(n24473),
	.b(south_input_NIB_storage_data_f_3__56_),
	.c(FE_OFN24744_n18648),
	.d(south_input_NIB_storage_data_f_0__56_));
   ao22f20 U23920 (.o(n18675),
	.a(n21315),
	.b(south_input_NIB_storage_data_f_2__56_),
	.c(n18061),
	.d(south_input_NIB_storage_data_f_1__56_));
   ao22f20 U23921 (.o(n18678),
	.a(n24473),
	.b(south_input_NIB_storage_data_f_3__57_),
	.c(FE_RN_62),
	.d(south_input_NIB_storage_data_f_0__57_));
   ao22f20 U23922 (.o(n18677),
	.a(FE_RN_17),
	.b(south_input_NIB_storage_data_f_2__57_),
	.c(n18061),
	.d(south_input_NIB_storage_data_f_1__57_));
   na02f20 U23923 (.o(n20641),
	.a(n18678),
	.b(n18677));
   ao22f20 U23924 (.o(n18679),
	.a(n19635),
	.b(FE_RN_68),
	.c(FE_OFN73_n19631),
	.d(n20641));
   na04f40 U23925 (.o(n18700),
	.a(n18682),
	.b(n18681),
	.c(n18680),
	.d(n18679));
   ao22f10 U23926 (.o(n18685),
	.a(n24473),
	.b(south_input_NIB_storage_data_f_3__52_),
	.c(FE_OFN24744_n18648),
	.d(south_input_NIB_storage_data_f_0__52_));
   ao22f20 U23927 (.o(n18687),
	.a(n24473),
	.b(south_input_NIB_storage_data_f_3__50_),
	.c(FE_RN_62),
	.d(south_input_NIB_storage_data_f_0__50_));
   na02f20 U23928 (.o(n23341),
	.a(n18687),
	.b(n18686));
   ao22f10 U23929 (.o(n18691),
	.a(n19647),
	.b(n21160),
	.c(n19657),
	.d(n23341));
   ao22f20 U23930 (.o(n18690),
	.a(n19347),
	.b(FE_RN_60),
	.c(n19387),
	.d(n20745));
   ao22f20 U23931 (.o(n18689),
	.a(FE_OFN53_n19355),
	.b(n23995),
	.c(n19617),
	.d(n23509));
   ao22f10 U23932 (.o(n18688),
	.a(myChipID_f_8_),
	.b(n23590),
	.c(myChipID_f_5_),
	.d(n21484));
   oa22f10 U23933 (.o(n18693),
	.a(n19622),
	.b(n25517),
	.c(n19584),
	.d(FE_RN_56));
   oa22f10 U23934 (.o(n18692),
	.a(n19666),
	.b(n23332),
	.c(n19594),
	.d(n25510));
   no02f10 U23935 (.o(n18697),
	.a(n18693),
	.b(n18692));
   oa22f10 U23936 (.o(n18695),
	.a(n19647),
	.b(n21160),
	.c(n19635),
	.d(n21332));
   oa22f10 U23937 (.o(n18694),
	.a(n19657),
	.b(n23341),
	.c(FE_OFN73_n19631),
	.d(FE_RN_44));
   no02f10 U23938 (.o(n18696),
	.a(n18695),
	.b(n18694));
   na02f20 U23939 (.o(n18698),
	.a(n18697),
	.b(n18696));
   ao22f08 U23940 (.o(n18702),
	.a(n17782),
	.b(south_input_NIB_storage_data_f_2__37_),
	.c(FE_OFN24742_n18683),
	.d(south_input_NIB_storage_data_f_1__37_));
   no02f10 U23941 (.o(n19038),
	.a(n19837),
	.b(n19839));
   no02f20 U23942 (.o(n19838),
	.a(myLocY_f_3_),
	.b(n22877));
   no02f20 U23943 (.o(n19848),
	.a(myLocY_f_4_),
	.b(n22884));
   no02f10 U23944 (.o(n19041),
	.a(n19851),
	.b(n18717));
   in01f08 U23945 (.o(n18724),
	.a(n18718));
   no03f20 U23946 (.o(n22928),
	.a(n18724),
	.b(n18723),
	.c(n18722));
   in01f10 U23947 (.o(n18731),
	.a(n22928));
   oa22f10 U23948 (.o(n19046),
	.a(n19518),
	.b(n18731),
	.c(FE_OFN65_n19542),
	.d(n18730));
   in01f08 U23949 (.o(n18732),
	.a(n19046));
   na02f10 U23950 (.o(n19836),
	.a(n19041),
	.b(n18732));
   no02f10 U23951 (.o(n19044),
	.a(myLocY_f_7_),
	.b(n22928));
   no02f10 U23952 (.o(n19849),
	.a(n19044),
	.b(n18734));
   no02f10 U23953 (.o(n19037),
	.a(n18735),
	.b(n19842));
   na02f10 U23954 (.o(n18736),
	.a(n19849),
	.b(n19037));
   na02f08 U23955 (.o(n18743),
	.a(n17782),
	.b(south_input_NIB_storage_data_f_2__44_));
   na02f10 U23956 (.o(n23493),
	.a(n18742),
	.b(n18741));
   no02f10 U23957 (.o(n18776),
	.a(n18775),
	.b(n18774));
   oa22f08 U23958 (.o(n18777),
	.a(myLocX_f_5_),
	.b(n18776),
	.c(myLocX_f_6_),
	.d(n22861));
   no02f10 U23959 (.o(n25050),
	.a(proc_output_current_route_connection_2_),
	.b(n25038));
   na02f10 U23960 (.o(n20501),
	.a(proc_output_current_route_connection_0_),
	.b(n25050));
   in01f02 U23961 (.o(n25486),
	.a(proc_input_NIB_elements_in_array_f_4_));
   na02f06 U23962 (.o(n18796),
	.a(n17782),
	.b(south_input_NIB_storage_data_f_2__30_));
   no02f40 U23965 (.o(n18959),
	.a(n18827),
	.b(FE_OCPN25899_west_input_NIB_head_ptr_f_0));
   no02f40 U23968 (.o(n18815),
	.a(west_input_NIB_head_ptr_f_1_),
	.b(west_input_NIB_head_ptr_f_0_));
   na02f08 U23970 (.o(n18816),
	.a(west_input_NIB_head_ptr_f_0_),
	.b(west_input_NIB_storage_data_f_1__44_));
   oa22f04 U23971 (.o(n18825),
	.a(west_input_NIB_head_ptr_f_1_),
	.b(n18821),
	.c(n18820),
	.d(FE_OCPN25820_west_input_NIB_head_ptr_f_1));
   oa22f04 U23972 (.o(n18824),
	.a(west_input_NIB_head_ptr_f_1_),
	.b(n18823),
	.c(n18822),
	.d(FE_OCPN25820_west_input_NIB_head_ptr_f_1));
   no02f10 U23974 (.o(n18872),
	.a(myLocX_f_3_),
	.b(n21342));
   no02f10 U23975 (.o(n18830),
	.a(n18826),
	.b(n18872));
   ao22f04 U23977 (.o(n18835),
	.a(FE_RN_5),
	.b(west_input_NIB_storage_data_f_3__43_),
	.c(FE_OFN27_n18974),
	.d(west_input_NIB_storage_data_f_0__43_));
   no02f40 U23979 (.o(n18828),
	.a(west_input_NIB_head_ptr_f_1_),
	.b(FE_OCPN25900_west_input_NIB_head_ptr_f_0));
   in01f06 U23982 (.o(n18834),
	.a(n18831));
   no02f10 U23983 (.o(n21403),
	.a(n18834),
	.b(n18833));
   ao22f10 U23984 (.o(n18871),
	.a(myLocX_f_2_),
	.b(n21403),
	.c(myLocX_f_3_),
	.d(n21342));
   in01f10 U23985 (.o(n18848),
	.a(n18871));
   no02f08 U23986 (.o(n18841),
	.a(n19708),
	.b(n18836));
   ao22f04 U23988 (.o(n18845),
	.a(FE_OFN27_n18974),
	.b(west_input_NIB_storage_data_f_0__42_),
	.c(n18960),
	.d(west_input_NIB_storage_data_f_2__42_));
   oa22f06 U23989 (.o(n18843),
	.a(FE_RN_47),
	.b(n18839),
	.c(FE_OCPN25926_n18828),
	.d(n18838));
   no03f20 U23990 (.o(n18964),
	.a(n18870),
	.b(n18848),
	.c(n18847));
   na02f10 U23991 (.o(n18851),
	.a(n18127),
	.b(west_input_NIB_storage_data_f_0__48_));
   oa12f10 U23992 (.o(n18853),
	.a(n18851),
	.b(n18852),
	.c(FE_RN_47));
   no03f20 U23993 (.o(n22859),
	.a(n18855),
	.b(n18854),
	.c(n18853));
   na02f08 U23994 (.o(n18858),
	.a(n18127),
	.b(west_input_NIB_storage_data_f_0__49_));
   oa12f08 U23995 (.o(n18860),
	.a(n18858),
	.b(n18859),
	.c(FE_RN_47));
   ao22f08 U23996 (.o(n18873),
	.a(myLocX_f_6_),
	.b(n22859),
	.c(myLocX_f_7_),
	.d(n22820));
   na02f04 U23997 (.o(n18865),
	.a(n18127),
	.b(west_input_NIB_storage_data_f_0__46_));
   ao22f04 U23998 (.o(n18868),
	.a(n18959),
	.b(west_input_NIB_storage_data_f_3__47_),
	.c(n18127),
	.d(west_input_NIB_storage_data_f_0__47_));
   ao22f08 U24000 (.o(n18867),
	.a(FE_OFN24764_n18960),
	.b(west_input_NIB_storage_data_f_2__47_),
	.c(n18828),
	.d(west_input_NIB_storage_data_f_1__47_));
   na02f10 U24001 (.o(n23323),
	.a(n18868),
	.b(n18867));
   na02f06 U24002 (.o(n18967),
	.a(n18873),
	.b(n20432));
   in01f03 U24003 (.o(n19725),
	.a(myLocX_f_6_));
   ao22f10 U24004 (.o(n20430),
	.a(n19701),
	.b(n23323),
	.c(n19725),
	.d(n18881));
   na02f20 U24007 (.o(n21465),
	.a(n18887),
	.b(n18886));
   no02f20 U24008 (.o(n18891),
	.a(n19666),
	.b(FE_RN_25));
   ao22f20 U24009 (.o(n18904),
	.a(FE_RN_64),
	.b(west_input_NIB_storage_data_f_3__57_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__57_));
   ao12f10 U24010 (.o(n18890),
	.a(myChipID_f_7_),
	.b(n20642),
	.c(n18904));
   ao12f20 U24012 (.o(n18889),
	.a(myChipID_f_10_),
	.b(n20747),
	.c(n20746));
   no04f20 U24013 (.o(n18903),
	.a(n18892),
	.b(n18891),
	.c(n18890),
	.d(n18889));
   no02f20 U24014 (.o(n18898),
	.a(n18995),
	.b(n18893));
   in01f10 U24015 (.o(n18899),
	.a(n23993));
   ao22f20 U24016 (.o(n18900),
	.a(FE_OFN53_n19355),
	.b(n18899),
	.c(n19633),
	.d(n23317));
   na04f40 U24017 (.o(n18947),
	.a(n18903),
	.b(n18902),
	.c(n18901),
	.d(n18900));
   in01f10 U24018 (.o(n20643),
	.a(n18904));
   no02f20 U24019 (.o(n18907),
	.a(FE_OFN73_n19631),
	.b(n20643));
   ao22f20 U24020 (.o(n18906),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__52_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__52_));
   ao22f20 U24021 (.o(n18905),
	.a(FE_OFN24763_n18960),
	.b(west_input_NIB_storage_data_f_2__52_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__52_));
   ao22f10 U24022 (.o(n18920),
	.a(n18907),
	.b(n20642),
	.c(n19647),
	.d(n21162));
   ao22f10 U24023 (.o(n18908),
	.a(FE_OFN24763_n18960),
	.b(west_input_NIB_storage_data_f_2__51_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__51_));
   na02f20 U24024 (.o(n21696),
	.a(n18909),
	.b(n18908));
   in01f10 U24025 (.o(n18914),
	.a(n21696));
   ao22f10 U24026 (.o(n18912),
	.a(FE_RN_64),
	.b(west_input_NIB_storage_data_f_3__63_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__63_));
   ao22f20 U24028 (.o(n18918),
	.a(myChipID_f_1_),
	.b(n18914),
	.c(myChipID_f_13_),
	.d(n18913));
   na04f40 U24031 (.o(n18946),
	.a(n18920),
	.b(n18919),
	.c(n18918),
	.d(n18917));
   no03f40 U24032 (.o(n24002),
	.a(n18926),
	.b(n18925),
	.c(n18924));
   ao22f10 U24033 (.o(n18944),
	.a(myChipID_f_11_),
	.b(n24002),
	.c(n19347),
	.d(FE_RN_65));
   no02f20 U24034 (.o(n18934),
	.a(n18995),
	.b(n18928));
   na02f40 U24035 (.o(n18930),
	.a(FE_RN_32),
	.b(west_input_NIB_storage_data_f_0__50_));
   no03f40 U24036 (.o(n18937),
	.a(n18934),
	.b(n18933),
	.c(n18932));
   ao22f20 U24037 (.o(n18943),
	.a(myChipID_f_0_),
	.b(n18937),
	.c(n19584),
	.d(n18935));
   in01f10 U24038 (.o(n18936),
	.a(n20746));
   no02f20 U24039 (.o(n18938),
	.a(n19387),
	.b(n18936));
   in01f20 U24040 (.o(n23340),
	.a(n18937));
   ao22f20 U24041 (.o(n18942),
	.a(n18938),
	.b(n20747),
	.c(n19657),
	.d(n23340));
   na04f40 U24042 (.o(n18945),
	.a(n18944),
	.b(n18943),
	.c(n18942),
	.d(n18941));
   ao22f10 U24043 (.o(n20589),
	.a(west_input_control_count_zero_f),
	.b(west_input_control_thanks_all_f),
	.c(west_input_control_header_last_f),
	.d(n20566));
   na02f10 U24044 (.o(n18948),
	.a(n20437),
	.b(FE_OFN24832_n25232));
   no02f20 U24045 (.o(n19014),
	.a(n20227),
	.b(n18948));
   no03f10 U24046 (.o(n19864),
	.a(n18967),
	.b(n18966),
	.c(n20429));
   oa12f10 U24047 (.o(n18981),
	.a(n18979),
	.b(n18980),
	.c(FE_RN_47));
   ao22f06 U24048 (.o(n18987),
	.a(FE_RN_8),
	.b(west_input_NIB_storage_data_f_3__38_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__38_));
   no04f10 U24049 (.o(n19010),
	.a(n20231),
	.b(n20230),
	.c(n20263),
	.d(n20229));
   na04f20 U24050 (.o(n19011),
	.a(n20437),
	.b(n19864),
	.c(n20233),
	.d(n19010));
   na02f20 U24051 (.o(n19013),
	.a(n19012),
	.b(n19011));
   no02f40 U24052 (.o(n23400),
	.a(n19014),
	.b(n19013));
   na02f10 U24053 (.o(n20259),
	.a(east_output_current_route_connection_1_),
	.b(n20318));
   no02f20 U24054 (.o(n19020),
	.a(east_output_current_route_connection_0_),
	.b(n20259));
   no02f10 U24055 (.o(n19022),
	.a(n19021),
	.b(n20259));
   no02f10 U24056 (.o(n19053),
	.a(n19030),
	.b(n19029));
   no03f06 U24057 (.o(n19032),
	.a(n19031),
	.b(n19064),
	.c(n20377));
   no02f10 U24058 (.o(n19034),
	.a(FE_RN_4),
	.b(n19033));
   no04f10 U24059 (.o(n19049),
	.a(n20286),
	.b(n19830),
	.c(n19829),
	.d(n20270));
   na03f10 U24060 (.o(n19050),
	.a(n20417),
	.b(n19049),
	.c(n20466));
   in01f01 U24061 (.o(n19061),
	.a(north_output_space_is_one_f));
   no02f10 U24062 (.o(n19070),
	.a(n25018),
	.b(n19067));
   no02f20 U24063 (.o(n19071),
	.a(north_input_NIB_head_ptr_f_1_),
	.b(n25109));
   in01f02 U24065 (.o(n19072),
	.a(north_input_NIB_storage_data_f_1__41_));
   no02f40 U24067 (.o(n19073),
	.a(north_input_NIB_head_ptr_f_0_),
	.b(FE_RN_45));
   in01f02 U24070 (.o(n19077),
	.a(north_input_NIB_storage_data_f_3__41_));
   na02f40 U24071 (.o(n19225),
	.a(north_input_NIB_head_ptr_f_0_),
	.b(north_input_NIB_head_ptr_f_1_));
   no02f40 U24074 (.o(n19075),
	.a(north_input_NIB_head_ptr_f_0_),
	.b(north_input_NIB_head_ptr_f_1_));
   na02f03 U24077 (.o(n19076),
	.a(FE_OFN24769_n19075),
	.b(north_input_NIB_storage_data_f_0__41_));
   oa12f08 U24080 (.o(n19134),
	.a(n19080),
	.b(n19081),
	.c(n19225));
   no02f08 U24081 (.o(n20158),
	.a(n19083),
	.b(n19082));
   ao22f04 U24083 (.o(n19085),
	.a(FE_OFN51_n19193),
	.b(north_input_NIB_storage_data_f_3__39_),
	.c(FE_OFN24769_n19075),
	.d(north_input_NIB_storage_data_f_0__39_));
   ao22f04 U24085 (.o(n19084),
	.a(FE_RN_11),
	.b(north_input_NIB_storage_data_f_2__39_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__39_));
   na02f08 U24088 (.o(n21141),
	.a(n19088),
	.b(n19087));
   no02f08 U24089 (.o(n19129),
	.a(n19133),
	.b(n19089));
   ao22f03 U24090 (.o(n19091),
	.a(FE_OFN24769_n19075),
	.b(north_input_NIB_storage_data_f_0__35_),
	.c(FE_RN_11),
	.d(north_input_NIB_storage_data_f_2__35_));
   ao22f06 U24091 (.o(n19090),
	.a(FE_OFN51_n19193),
	.b(north_input_NIB_storage_data_f_3__35_),
	.c(n24364),
	.d(north_input_NIB_storage_data_f_1__35_));
   na02f10 U24092 (.o(n19123),
	.a(n19091),
	.b(n19090));
   ao22f04 U24093 (.o(n19098),
	.a(FE_OFN51_n19193),
	.b(north_input_NIB_storage_data_f_3__37_),
	.c(FE_OFN24769_n19075),
	.d(north_input_NIB_storage_data_f_0__37_));
   na02f08 U24094 (.o(n20784),
	.a(n19098),
	.b(n19097));
   no02f06 U24095 (.o(n19127),
	.a(n19321),
	.b(n20784));
   in01f02 U24096 (.o(n19103),
	.a(north_input_NIB_storage_data_f_1__31_));
   in01f04 U24098 (.o(n19106),
	.a(north_input_NIB_storage_data_f_3__31_));
   na02f06 U24099 (.o(n19105),
	.a(FE_OFN24770_n19075),
	.b(north_input_NIB_storage_data_f_0__31_));
   oa12f04 U24100 (.o(n19107),
	.a(n19105),
	.b(n19106),
	.c(n19225));
   in01f02 U24101 (.o(n19110),
	.a(north_input_NIB_storage_data_f_1__30_));
   in01f02 U24102 (.o(n19113),
	.a(north_input_NIB_storage_data_f_3__30_));
   na02f08 U24103 (.o(n19121),
	.a(n19321),
	.b(n20784));
   na02f08 U24104 (.o(n19124),
	.a(FE_OFN67_n19548),
	.b(n23967));
   no02f10 U24105 (.o(n19126),
	.a(myLocY_f_0_),
	.b(n22829));
   na02f10 U24106 (.o(n19144),
	.a(n21893),
	.b(n20158));
   na02f06 U24107 (.o(n19130),
	.a(n19129),
	.b(n19128));
   ao22f10 U24108 (.o(n19148),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__53_),
	.c(FE_OFN24769_n19075),
	.d(north_input_NIB_storage_data_f_0__53_));
   ao22f08 U24110 (.o(n19151),
	.a(FE_RN_10),
	.b(north_input_NIB_storage_data_f_3__51_),
	.c(FE_OFN24773_n19075),
	.d(north_input_NIB_storage_data_f_0__51_));
   ao22f10 U24111 (.o(n19154),
	.a(FE_OFN24774_n19073),
	.b(north_input_NIB_storage_data_f_2__52_),
	.c(FE_OFN25610_n19071),
	.d(north_input_NIB_storage_data_f_1__52_));
   ao22f06 U24113 (.o(n19156),
	.a(n21865),
	.b(north_input_NIB_storage_data_f_2__58_),
	.c(FE_OFN25610_n19071),
	.d(north_input_NIB_storage_data_f_1__58_));
   ao22f10 U24114 (.o(n19155),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__58_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__58_));
   no02f20 U24115 (.o(n19164),
	.a(FE_OFN24776_n19073),
	.b(n19157));
   no02f10 U24116 (.o(n19163),
	.a(n19223),
	.b(n19158));
   na02f20 U24117 (.o(n19160),
	.a(FE_OFN24768_n19075),
	.b(north_input_NIB_storage_data_f_0__50_));
   ao22f20 U24118 (.o(n19167),
	.a(FE_OFN96_n21865),
	.b(north_input_NIB_storage_data_f_2__56_),
	.c(FE_OFN25610_n19071),
	.d(north_input_NIB_storage_data_f_1__56_));
   in01f10 U24119 (.o(n19168),
	.a(n23613));
   no02f08 U24120 (.o(n19169),
	.a(n19635),
	.b(n23613));
   no02f10 U24121 (.o(n19184),
	.a(n19170),
	.b(n19169));
   ao22f10 U24122 (.o(n19171),
	.a(FE_RN_10),
	.b(north_input_NIB_storage_data_f_3__54_),
	.c(FE_OFN24773_n19075),
	.d(north_input_NIB_storage_data_f_0__54_));
   no02f20 U24123 (.o(n19173),
	.a(FE_OFN53_n19355),
	.b(n23994));
   ao12f10 U24124 (.o(n19183),
	.a(n19173),
	.b(FE_OFN53_n19355),
	.c(n23994));
   ao22f10 U24125 (.o(n19174),
	.a(FE_RN_10),
	.b(north_input_NIB_storage_data_f_3__61_),
	.c(FE_OFN24773_n19075),
	.d(north_input_NIB_storage_data_f_0__61_));
   no02f20 U24126 (.o(n19176),
	.a(n19584),
	.b(n24003));
   ao12f10 U24127 (.o(n19182),
	.a(n19176),
	.b(n19584),
	.c(n24003));
   ao22f08 U24128 (.o(n19178),
	.a(FE_OFN24774_n19073),
	.b(north_input_NIB_storage_data_f_2__62_),
	.c(FE_OFN25610_n19071),
	.d(north_input_NIB_storage_data_f_1__62_));
   na02f10 U24129 (.o(n21408),
	.a(n19178),
	.b(n19177));
   na02f10 U24130 (.o(n19188),
	.a(n19180),
	.b(n19179));
   na04f20 U24131 (.o(n19202),
	.a(n19184),
	.b(n19183),
	.c(n19182),
	.d(n19181));
   ao22f10 U24132 (.o(n19186),
	.a(n21865),
	.b(north_input_NIB_storage_data_f_2__55_),
	.c(FE_OFN25610_n19071),
	.d(north_input_NIB_storage_data_f_1__55_));
   ao22f10 U24133 (.o(n19185),
	.a(FE_RN_10),
	.b(north_input_NIB_storage_data_f_3__55_),
	.c(FE_OFN24772_n19075),
	.d(north_input_NIB_storage_data_f_0__55_));
   ao22f10 U24134 (.o(n19190),
	.a(n21865),
	.b(north_input_NIB_storage_data_f_2__63_),
	.c(FE_OFN25610_n19071),
	.d(north_input_NIB_storage_data_f_1__63_));
   ao22f10 U24135 (.o(n19199),
	.a(n22869),
	.b(myChipID_f_7_),
	.c(n19617),
	.d(n23510));
   in01f08 U24136 (.o(n19191),
	.a(n23510));
   ao22f10 U24137 (.o(n19198),
	.a(n21485),
	.b(myChipID_f_5_),
	.c(n19191),
	.d(myChipID_f_13_));
   ao22f20 U24138 (.o(n19195),
	.a(FE_OFN96_n21865),
	.b(north_input_NIB_storage_data_f_2__60_),
	.c(FE_OFN25610_n19071),
	.d(north_input_NIB_storage_data_f_1__60_));
   ao22f20 U24139 (.o(n19194),
	.a(FE_OFN48_n19193),
	.b(north_input_NIB_storage_data_f_3__60_),
	.c(FE_OFN24773_n19075),
	.d(north_input_NIB_storage_data_f_0__60_));
   na02f20 U24140 (.o(n23542),
	.a(n19195),
	.b(n19194));
   na04f40 U24141 (.o(n19201),
	.a(n19200),
	.b(n19199),
	.c(n19198),
	.d(n19197));
   no03f40 U24142 (.o(n20152),
	.a(n19203),
	.b(n19202),
	.c(n19201));
   na02f08 U24143 (.o(n19230),
	.a(n19205),
	.b(n19204));
   ao22f06 U24144 (.o(n19207),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__43_),
	.c(FE_OFN24770_n19075),
	.d(north_input_NIB_storage_data_f_0__43_));
   no02f10 U24146 (.o(n19233),
	.a(n20394),
	.b(n20392));
   no02f10 U24147 (.o(n19228),
	.a(myLocX_f_6_),
	.b(n22860));
   ao22f06 U24148 (.o(n19238),
	.a(FE_OFN51_n19193),
	.b(north_input_NIB_storage_data_f_3__49_),
	.c(FE_RN_11),
	.d(north_input_NIB_storage_data_f_2__49_));
   no02f10 U24150 (.o(n19232),
	.a(myLocX_f_0_),
	.b(FE_OFN25638_n19230));
   na04f20 U24151 (.o(n19242),
	.a(n20389),
	.b(n19233),
	.c(n20400),
	.d(n20301));
   no02f10 U24152 (.o(n19236),
	.a(n19234),
	.b(myLocX_f_2_));
   na02f10 U24153 (.o(n20298),
	.a(n20395),
	.b(n20303));
   no03f20 U24154 (.o(n19243),
	.a(n19242),
	.b(n20387),
	.c(n20298));
   na02f20 U24155 (.o(n20297),
	.a(n20152),
	.b(n19243));
   no02f10 U24156 (.o(n20110),
	.a(n19244),
	.b(n20297));
   no02f40 U24158 (.o(n20504),
	.a(FE_RN_9),
	.b(n20109));
   no02f01 U24159 (.o(n19249),
	.a(south_output_space_is_one_f),
	.b(south_output_space_yummy_f));
   in01f01 U24160 (.o(n19250),
	.a(south_output_space_yummy_f));
   in01f02 U24162 (.o(n19259),
	.a(east_input_NIB_storage_data_f_2__43_));
   no02f40 U24163 (.o(n19932),
	.a(east_input_NIB_head_ptr_f_0_),
	.b(east_input_NIB_head_ptr_f_1_));
   in01f02 U24165 (.o(n19258),
	.a(east_input_NIB_storage_data_f_0__43_));
   na02f40 U24167 (.o(n20506),
	.a(east_input_NIB_head_ptr_f_1_),
	.b(east_input_NIB_head_ptr_f_0_));
   ao22f10 U24173 (.o(n19266),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__44_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__44_));
   na02f10 U24174 (.o(n19269),
	.a(FE_OFN24777_n19932),
	.b(east_input_NIB_storage_data_f_0__42_));
   na02f08 U24178 (.o(n19282),
	.a(n19795),
	.b(n19281));
   oa22f04 U24179 (.o(n19288),
	.a(FE_OFN25663_n19914),
	.b(n19285),
	.c(n20506),
	.d(n19284));
   oa22f08 U24180 (.o(n19287),
	.a(n21858),
	.b(n19286),
	.c(FE_OFN60_n19435),
	.d(n24919));
   no02f10 U24181 (.o(n22819),
	.a(n19288),
	.b(n19287));
   no02f08 U24182 (.o(n19411),
	.a(myLocX_f_7_),
	.b(n22819));
   oa22f04 U24183 (.o(n19293),
	.a(FE_OFN25663_n19914),
	.b(n19290),
	.c(n20506),
	.d(n19289));
   oa22f08 U24184 (.o(n19292),
	.a(n21858),
	.b(n19291),
	.c(n19435),
	.d(n24909));
   in01f01 U24185 (.o(n19297),
	.a(east_input_NIB_storage_data_f_2__30_));
   in01f01 U24186 (.o(n19296),
	.a(east_input_NIB_storage_data_f_3__30_));
   in01f01 U24187 (.o(n19298),
	.a(east_input_NIB_storage_data_f_0__30_));
   in01f02 U24188 (.o(n24787),
	.a(east_input_NIB_storage_data_f_1__30_));
   in01f01 U24189 (.o(n19301),
	.a(east_input_NIB_storage_data_f_3__32_));
   oa22f01 U24190 (.o(n19305),
	.a(FE_OFN25664_n19914),
	.b(n19302),
	.c(n20506),
	.d(n19301));
   in01f01 U24191 (.o(n19303),
	.a(east_input_NIB_storage_data_f_0__32_));
   in01f02 U24192 (.o(n24887),
	.a(east_input_NIB_storage_data_f_1__32_));
   oa22f01 U24193 (.o(n19304),
	.a(n21858),
	.b(n19303),
	.c(n19435),
	.d(n24887));
   ao22f01 U24194 (.o(n19307),
	.a(FE_RN_69),
	.b(east_input_NIB_storage_data_f_1__31_),
	.c(n19400),
	.d(east_input_NIB_storage_data_f_3__31_));
   na02f03 U24196 (.o(n19310),
	.a(FE_OFN24777_n19932),
	.b(east_input_NIB_storage_data_f_0__34_));
   ao22f06 U24197 (.o(n19317),
	.a(FE_OFN24777_n19932),
	.b(east_input_NIB_storage_data_f_0__36_),
	.c(n19400),
	.d(east_input_NIB_storage_data_f_3__36_));
   ao22f04 U24198 (.o(n19320),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__37_),
	.c(n19400),
	.d(east_input_NIB_storage_data_f_3__37_));
   na02f20 U24199 (.o(n25519),
	.a(n19332),
	.b(n19331));
   no02f10 U24200 (.o(n19336),
	.a(n19622),
	.b(n25519));
   in01f10 U24201 (.o(n22904),
	.a(n25519));
   no02f20 U24202 (.o(n19335),
	.a(myChipID_f_9_),
	.b(n22904));
   ao22f20 U24203 (.o(n21289),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__50_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__50_));
   ao22f10 U24204 (.o(n21288),
	.a(FE_OFN24780_n19932),
	.b(east_input_NIB_storage_data_f_0__50_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__50_));
   ao12f20 U24205 (.o(n19334),
	.a(myChipID_f_0_),
	.b(n21289),
	.c(n21288));
   ao22f20 U24206 (.o(n21295),
	.a(FE_OFN25661_n19914),
	.b(east_input_NIB_storage_data_f_2__63_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__63_));
   ao22f10 U24207 (.o(n21294),
	.a(FE_OFN24780_n19932),
	.b(east_input_NIB_storage_data_f_0__63_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__63_));
   ao12f20 U24208 (.o(n19333),
	.a(myChipID_f_13_),
	.b(n21295),
	.c(n21294));
   no02f10 U24209 (.o(n19341),
	.a(FE_OFN25663_n19914),
	.b(n19337));
   no02f10 U24210 (.o(n19340),
	.a(FE_RN_57),
	.b(n24765));
   ao22f10 U24211 (.o(n19360),
	.a(n22889),
	.b(myChipID_f_12_),
	.c(n19635),
	.d(n23611));
   ao22f10 U24212 (.o(n19344),
	.a(FE_OFN24780_n19932),
	.b(east_input_NIB_storage_data_f_0__51_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__51_));
   na02f10 U24213 (.o(n25512),
	.a(n19345),
	.b(n19344));
   na02f20 U24214 (.o(n19349),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__54_));
   oa22f20 U24215 (.o(n19356),
	.a(n19594),
	.b(FE_RN_14),
	.c(FE_OFN53_n19355),
	.d(n19354));
   ao22f10 U24216 (.o(n19363),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__61_),
	.c(FE_RN_69),
	.d(east_input_NIB_storage_data_f_1__61_));
   na02f20 U24217 (.o(n19372),
	.a(n19363),
	.b(n19362));
   no02f20 U24219 (.o(n19365),
	.a(n19657),
	.b(n19364));
   ao22f20 U24220 (.o(n19391),
	.a(myChipID_f_11_),
	.b(n24001),
	.c(n21289),
	.d(n19365));
   no02f06 U24221 (.o(n19370),
	.a(FE_OFN25663_n19914),
	.b(n19366));
   na02f10 U24222 (.o(n19367),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__57_));
   oa12f10 U24223 (.o(n19369),
	.a(n19367),
	.b(n20506),
	.c(n19368));
   no03f20 U24224 (.o(n22866),
	.a(n19371),
	.b(n19370),
	.c(n19369));
   ao22f10 U24225 (.o(n19390),
	.a(n22866),
	.b(myChipID_f_7_),
	.c(n19584),
	.d(n19372));
   na02f20 U24226 (.o(n19374),
	.a(FE_OFN24780_n19932),
	.b(east_input_NIB_storage_data_f_0__53_));
   ao22f20 U24227 (.o(n19389),
	.a(myChipID_f_3_),
	.b(n19379),
	.c(FE_OFN73_n19631),
	.d(n19378));
   in01f10 U24228 (.o(n23330),
	.a(n19379));
   na02f10 U24229 (.o(n19381),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__60_));
   ao22f20 U24230 (.o(n19388),
	.a(n19666),
	.b(n23330),
	.c(n19387),
	.d(n19386));
   na04f40 U24231 (.o(n19409),
	.a(n19391),
	.b(n19390),
	.c(n19389),
	.d(n19388));
   ao22f10 U24232 (.o(n19392),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__52_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__52_));
   in01f10 U24233 (.o(n21163),
	.a(n19394));
   ao22f20 U24234 (.o(n19396),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__55_),
	.c(FE_OCPN25813_FE_OFN24735_n19306),
	.d(east_input_NIB_storage_data_f_1__55_));
   ao22f10 U24235 (.o(n19395),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__55_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__55_));
   ao22f20 U24236 (.o(n19406),
	.a(myChipID_f_2_),
	.b(n21163),
	.c(n19633),
	.d(n23316));
   no02f20 U24237 (.o(n19398),
	.a(n19617),
	.b(n19397));
   ao22f20 U24238 (.o(n19405),
	.a(myChipID_f_5_),
	.b(n19399),
	.c(n21295),
	.d(n19398));
   ao22f10 U24240 (.o(n19401),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__58_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__58_));
   na02f20 U24241 (.o(n23586),
	.a(n19402),
	.b(n19401));
   no02f10 U24242 (.o(n19403),
	.a(n19575),
	.b(n23586));
   ao12f10 U24243 (.o(n19404),
	.a(n19403),
	.b(n19575),
	.c(n23586));
   na03f20 U24244 (.o(n19444),
	.a(n20147),
	.b(n20514),
	.c(n20252));
   no02f10 U24245 (.o(n22881),
	.a(n19420),
	.b(n19419));
   no02f10 U24247 (.o(n22925),
	.a(n19431),
	.b(n19430));
   na02f08 U24248 (.o(n19812),
	.a(myLocY_f_7_),
	.b(n22925));
   no02f10 U24249 (.o(n19810),
	.a(myLocY_f_7_),
	.b(n22925));
   no02f06 U24250 (.o(n19440),
	.a(myLocY_f_5_),
	.b(n22851));
   na02f02 U24251 (.o(n19448),
	.a(east_input_control_thanks_all_f),
	.b(east_input_control_count_zero_f));
   no02f20 U24252 (.o(n19465),
	.a(n26016),
	.b(n26019));
   in01f01 U24253 (.o(n25112),
	.a(proc_input_NIB_elements_in_array_f_0_));
   na02s01 U24254 (.o(n25044),
	.a(n25974),
	.b(proc_input_NIB_elements_in_array_f_0_));
   no04f02 U24255 (.o(n19467),
	.a(reset),
	.b(proc_input_NIB_elements_in_array_f_1_),
	.c(n18408),
	.d(n18407));
   na02f02 U24256 (.o(n2848),
	.a(n19470),
	.b(n19469));
   no02f10 U24257 (.o(n25992),
	.a(n23400),
	.b(n20323));
   in01f01 U24258 (.o(n19482),
	.a(n19481));
   in01s01 U24259 (.o(n25268),
	.a(south_input_NIB_elements_in_array_f_0_));
   in01s01 U24260 (.o(n25897),
	.a(validIn_S));
   no02s01 U24261 (.o(n25347),
	.a(south_input_NIB_elements_in_array_f_0_),
	.b(validIn_S));
   in01f02 U24262 (.o(n19491),
	.a(n19485));
   na03f01 U24263 (.o(n19486),
	.a(south_input_NIB_elements_in_array_f_2_),
	.b(south_input_NIB_elements_in_array_f_1_),
	.c(n17888));
   in01f02 U24264 (.o(n19490),
	.a(n19487));
   in01s01 U24265 (.o(n25345),
	.a(south_input_NIB_elements_in_array_f_1_));
   no02s01 U24266 (.o(n19488),
	.a(south_input_NIB_elements_in_array_f_2_),
	.b(n25345));
   ao22s01 U24267 (.o(n19489),
	.a(n19488),
	.b(south_input_NIB_elements_in_array_f_0_),
	.c(south_input_NIB_elements_in_array_f_2_),
	.d(n25345));
   oa22f02 U24268 (.o(n3003),
	.a(n19492),
	.b(n19491),
	.c(n19490),
	.d(n18606));
   na02f40 U24271 (.o(n19507),
	.a(proc_input_NIB_head_ptr_f_2_),
	.b(n19496));
   na02f10 U24273 (.o(n19497),
	.a(proc_input_NIB_head_ptr_f_2_),
	.b(proc_input_NIB_head_ptr_f_1_));
   no03f20 U24274 (.o(n19498),
	.a(proc_input_NIB_head_ptr_f_3_),
	.b(n20508),
	.c(n19497));
   no02f40 U24275 (.o(n19499),
	.a(proc_input_NIB_head_ptr_f_1_),
	.b(proc_input_NIB_head_ptr_f_0_));
   na02f40 U24277 (.o(n19505),
	.a(proc_input_NIB_head_ptr_f_2_),
	.b(proc_input_NIB_head_ptr_f_3_));
   no02f20 U24278 (.o(n19500),
	.a(n19506),
	.b(n19505));
   no02f40 U24280 (.o(n19501),
	.a(proc_input_NIB_head_ptr_f_3_),
	.b(proc_input_NIB_head_ptr_f_2_));
   na02f40 U24283 (.o(n25072),
	.a(proc_input_NIB_head_ptr_f_0_),
	.b(proc_input_NIB_head_ptr_f_1_));
   na02f80 U24284 (.o(n25140),
	.a(proc_input_NIB_head_ptr_f_1_),
	.b(n20508));
   no02f40 U24285 (.o(n19503),
	.a(n19507),
	.b(n25140));
   na04f10 U24294 (.o(n19559),
	.a(n19558),
	.b(n19557),
	.c(n19556),
	.d(n19555));
   ao22f08 U24296 (.o(n19570),
	.a(n17754),
	.b(proc_input_NIB_storage_data_f_3__58_),
	.c(FE_OFN165_n24129),
	.d(proc_input_NIB_storage_data_f_1__58_));
   ao22f08 U24298 (.o(n19573),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__58_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__58_));
   ao22f08 U24299 (.o(n19572),
	.a(FE_OCPN25947_n19595),
	.b(proc_input_NIB_storage_data_f_15__58_),
	.c(FE_OCPN25924_n19547),
	.d(proc_input_NIB_storage_data_f_11__58_));
   ao22f08 U24300 (.o(n19582),
	.a(FE_OCPN25962_n18039),
	.b(proc_input_NIB_storage_data_f_10__61_),
	.c(FE_OFN168_n24343),
	.d(proc_input_NIB_storage_data_f_8__61_));
   ao22f06 U24301 (.o(n19586),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__51_),
	.c(FE_OCPN25814_FE_OFN186_n24453),
	.d(proc_input_NIB_storage_data_f_2__51_));
   na02f10 U24302 (.o(n19587),
	.a(proc_input_NIB_storage_data_f_9__51_),
	.b(FE_OFN25681_n17814));
   ao22f20 U24303 (.o(n19593),
	.a(FE_OCPN25836_n24342),
	.b(proc_input_NIB_storage_data_f_0__51_),
	.c(FE_OFN25673_n18033),
	.d(proc_input_NIB_storage_data_f_11__51_));
   ao22f10 U24304 (.o(n19596),
	.a(FE_OCPN25814_FE_OFN186_n24453),
	.b(proc_input_NIB_storage_data_f_2__63_),
	.c(FE_OFN25673_n18033),
	.d(proc_input_NIB_storage_data_f_11__63_));
   na02f10 U24305 (.o(n19605),
	.a(n19604),
	.b(n19603));
   ao22f08 U24306 (.o(n19610),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__60_),
	.c(FE_OFN20_n17779),
	.d(proc_input_NIB_storage_data_f_7__60_));
   ao22f08 U24307 (.o(n19607),
	.a(FE_OFN25681_n17814),
	.b(proc_input_NIB_storage_data_f_9__60_),
	.c(FE_OCPN25924_n19547),
	.d(proc_input_NIB_storage_data_f_11__60_));
   na04f20 U24308 (.o(n19616),
	.a(n19610),
	.b(n19609),
	.c(n19608),
	.d(n19607));
   na04f20 U24310 (.o(n19615),
	.a(n19614),
	.b(n19613),
	.c(n19612),
	.d(n19611));
   na02f10 U24311 (.o(n19626),
	.a(n19619),
	.b(n19618));
   in01f08 U24312 (.o(n19623),
	.a(n25520));
   oa22f20 U24313 (.o(n19624),
	.a(myChipID_f_9_),
	.b(n19623),
	.c(myChipID_f_10_),
	.d(n18102));
   oa22f20 U24314 (.o(n19652),
	.a(myChipID_f_7_),
	.b(n22873),
	.c(n19630),
	.d(n18101));
   oa22f20 U24315 (.o(n19651),
	.a(myChipID_f_6_),
	.b(n23619),
	.c(n19632),
	.d(FE_OFN73_n19631));
   ao22f08 U24317 (.o(n19658),
	.a(FE_OCPN25968_n19500),
	.b(proc_input_NIB_storage_data_f_12__53_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__53_));
   ao22f08 U24320 (.o(n19661),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__53_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__53_));
   no04f20 U24321 (.o(n19671),
	.a(n19670),
	.b(n19669),
	.c(n19668),
	.d(n19667));
   na02f06 U24322 (.o(n19723),
	.a(n19683),
	.b(n19682));
   no02f08 U24323 (.o(n20362),
	.a(n20374),
	.b(n20375));
   na02f10 U24324 (.o(n20361),
	.a(n19703),
	.b(n20366));
   ao22f04 U24325 (.o(n19710),
	.a(FE_OCPN25949_n18039),
	.b(proc_input_NIB_storage_data_f_10__42_),
	.c(FE_OFN156_n24129),
	.d(proc_input_NIB_storage_data_f_1__42_));
   ao22f06 U24326 (.o(n19714),
	.a(n24060),
	.b(proc_input_NIB_storage_data_f_9__42_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__42_));
   no02f10 U24327 (.o(n20368),
	.a(myLocX_f_3_),
	.b(n19734));
   na02f02 U24328 (.o(n19754),
	.a(n19753),
	.b(n19752));
   na02f02 U24329 (.o(n19774),
	.a(n19773),
	.b(n19772));
   no02f06 U24330 (.o(n19782),
	.a(n19781),
	.b(n19780));
   in01f02 U24331 (.o(n19859),
	.a(n19784));
   in01m02 U24332 (.o(n19791),
	.a(n20250));
   na02f04 U24333 (.o(n19821),
	.a(n20245),
	.b(n19791));
   na03f10 U24334 (.o(n19801),
	.a(n19825),
	.b(n19793),
	.c(n19792));
   na02f04 U24336 (.o(n19798),
	.a(n19797),
	.b(n19820));
   in01f04 U24337 (.o(n19799),
	.a(n19798));
   na02f10 U24338 (.o(n19800),
	.a(FE_RN_6),
	.b(n19799));
   in01f02 U24339 (.o(n23486),
	.a(n25002));
   oa12m02 U24340 (.o(n19843),
	.a(n19840),
	.b(n19842),
	.c(n19841));
   no02f04 U24341 (.o(n19889),
	.a(n20344),
	.b(n19858));
   no02f04 U24342 (.o(n24976),
	.a(n19861),
	.b(n19860));
   in01f01 U24343 (.o(n19863),
	.a(proc_input_control_header_last_f));
   na02f02 U24344 (.o(n19862),
	.a(proc_input_control_thanks_all_f),
	.b(proc_input_control_count_zero_f));
   na02f01 U24345 (.o(n19870),
	.a(n21426),
	.b(n23479));
   no02f02 U24346 (.o(n19872),
	.a(n24996),
	.b(n19870));
   in01f01 U24347 (.o(n19875),
	.a(n19874));
   na02f02 U24348 (.o(n20189),
	.a(n19876),
	.b(n19875));
   na02f04 U24351 (.o(n21431),
	.a(n19913),
	.b(n19912));
   na02f02 U24352 (.o(n19915),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__26_));
   oa22f01 U24356 (.o(n19919),
	.a(n21858),
	.b(n19918),
	.c(n20506),
	.d(n19917));
   na02f01 U24358 (.o(n19923),
	.a(FE_OFN24800_n20506),
	.b(east_input_NIB_storage_data_f_3__25_));
   na02f01 U24359 (.o(n19922),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__25_));
   na02f02 U24360 (.o(n19928),
	.a(n19923),
	.b(n19922));
   na02f01 U24361 (.o(n19926),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__25_));
   na02f02 U24362 (.o(n19925),
	.a(FE_RN_69),
	.b(east_input_NIB_storage_data_f_1__25_));
   na02f02 U24363 (.o(n19927),
	.a(n19926),
	.b(n19925));
   na02f01 U24364 (.o(n19931),
	.a(FE_OFN24800_n20506),
	.b(east_input_NIB_storage_data_f_3__27_));
   na02f01 U24365 (.o(n19930),
	.a(FE_OFN25662_n19914),
	.b(east_input_NIB_storage_data_f_2__27_));
   na02f02 U24366 (.o(n19937),
	.a(n19931),
	.b(n19930));
   na02f01 U24367 (.o(n19935),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__27_));
   na02f01 U24368 (.o(n19934),
	.a(FE_RN_69),
	.b(east_input_NIB_storage_data_f_1__27_));
   in01s01 U24369 (.o(n19951),
	.a(east_input_control_count_one_f));
   no02f01 U24370 (.o(n19950),
	.a(east_input_control_thanks_all_f),
	.b(east_input_control_tail_last_f));
   ao12f02 U24371 (.o(n19952),
	.a(n19950),
	.b(east_input_control_thanks_all_f),
	.c(n19951));
   na02f01 U24372 (.o(n19956),
	.a(n20343),
	.b(n19955));
   in01s01 U24373 (.o(n20563),
	.a(south_input_control_thanks_all_f));
   na02m02 U24374 (.o(n19986),
	.a(n19982),
	.b(n19981));
   na02f08 U24375 (.o(n25231),
	.a(n19993),
	.b(n19992));
   na02f06 U24376 (.o(n24029),
	.a(n19995),
	.b(n19994));
   na02f06 U24377 (.o(n23951),
	.a(n19997),
	.b(n19996));
   no02f04 U24378 (.o(n20000),
	.a(n23951),
	.b(n23621));
   in01s01 U24379 (.o(n20005),
	.a(west_input_control_count_one_f));
   no02s01 U24380 (.o(n20004),
	.a(west_input_control_thanks_all_f),
	.b(west_input_control_tail_last_f));
   na02f02 U24381 (.o(n20023),
	.a(n20022),
	.b(n20021));
   no02f06 U24382 (.o(n20116),
	.a(n25026),
	.b(n20111));
   oa22f02 U24383 (.o(south_output_control_N467),
	.a(n20125),
	.b(n20124),
	.c(n20123),
	.d(n24988));
   no02f10 U24384 (.o(n25994),
	.a(n23400),
	.b(n20324));
   no03f20 U24385 (.o(n26017),
	.a(n20529),
	.b(n20528),
	.c(n20531));
   in01s01 U24386 (.o(n25379),
	.a(west_input_NIB_elements_in_array_f_1_));
   no02s01 U24387 (.o(n20126),
	.a(west_input_NIB_elements_in_array_f_2_),
	.b(n25379));
   ao22s01 U24388 (.o(n20128),
	.a(n20126),
	.b(west_input_NIB_elements_in_array_f_0_),
	.c(west_input_NIB_elements_in_array_f_2_),
	.d(n25379));
   na03s01 U24389 (.o(n20129),
	.a(west_input_NIB_elements_in_array_f_2_),
	.b(west_input_NIB_elements_in_array_f_1_),
	.c(n17888));
   in01s01 U24390 (.o(n25234),
	.a(west_input_NIB_elements_in_array_f_0_));
   in01s01 U24391 (.o(n25929),
	.a(validIn_W));
   no02m01 U24392 (.o(n20148),
	.a(n25003),
	.b(n25002));
   no02f04 U24393 (.o(n20151),
	.a(n20149),
	.b(n20148));
   no03f02 U24394 (.o(n20179),
	.a(n20408),
	.b(n25010),
	.c(n20292));
   na02f02 U24395 (.o(n20171),
	.a(n20170),
	.b(n20169));
   no03f03 U24396 (.o(n20174),
	.a(n20173),
	.b(n20172),
	.c(n20171));
   in01f06 U24397 (.o(n20178),
	.a(n20177));
   ao12f02 U24398 (.o(n20188),
	.a(n20181),
	.b(n20183),
	.c(n20182));
   no02f02 U24399 (.o(n20194),
	.a(n20188),
	.b(n20187));
   no02f01 U24400 (.o(n20192),
	.a(n20190),
	.b(n20189));
   na03f01 U24401 (.o(n20197),
	.a(FE_OFN24833_n25232),
	.b(n20196),
	.c(n23479));
   no02m02 U24402 (.o(n20237),
	.a(n20265),
	.b(n20228));
   no03m02 U24403 (.o(n20232),
	.a(n20231),
	.b(n20230),
	.c(n20229));
   na02m02 U24404 (.o(n20260),
	.a(n20233),
	.b(n20232));
   in01m01 U24405 (.o(n20234),
	.a(n20260));
   na02m02 U24406 (.o(n20235),
	.a(n20450),
	.b(n20234));
   na03m02 U24407 (.o(n20239),
	.a(n25003),
	.b(n25001),
	.c(n23486));
   ao12f04 U24408 (.o(n20249),
	.a(n20244),
	.b(n20246),
	.c(n20245));
   oa12f02 U24409 (.o(n20253),
	.a(n20248),
	.b(n20250),
	.c(n20249));
   ao22f04 U24410 (.o(n20256),
	.a(n20254),
	.b(n20253),
	.c(n20252),
	.d(n20251));
   na02f02 U24412 (.o(n20290),
	.a(n20289),
	.b(n20288));
   oa12f04 U24413 (.o(n25393),
	.a(n20290),
	.b(n25007),
	.c(n20291));
   no02f06 U24415 (.o(n20311),
	.a(n20294),
	.b(n20295));
   oa22f06 U24416 (.o(n20316),
	.a(n20315),
	.b(n20314),
	.c(n20313),
	.d(n25397));
   no02f02 U24417 (.o(n20322),
	.a(n25017),
	.b(n20517));
   no03f10 U24418 (.o(n20326),
	.a(n20325),
	.b(n20548),
	.c(n20547));
   na02s01 U24419 (.o(n20327),
	.a(east_output_current_route_connection_0_),
	.b(FE_OFN25598_reset));
   in01f02 U24420 (.o(n25830),
	.a(validIn_N));
   in01s01 U24421 (.o(n25289),
	.a(north_input_NIB_elements_in_array_f_0_));
   na02m02 U24422 (.o(n20340),
	.a(n22517),
	.b(n24959));
   na02f02 U24423 (.o(n24974),
	.a(n22518),
	.b(n24952));
   in01s01 U24424 (.o(n20353),
	.a(n25176));
   na02s02 U24425 (.o(n25168),
	.a(west_output_current_route_connection_1_),
	.b(n20531));
   oa22f08 U24426 (.o(n20354),
	.a(n20531),
	.b(n25079),
	.c(n22216),
	.d(n25168));
   oa12f04 U24427 (.o(n20359),
	.a(n20357),
	.b(n20427),
	.c(n20358));
   na02f08 U24428 (.o(n20530),
	.a(n20360),
	.b(n20359));
   no03f06 U24429 (.o(n20367),
	.a(n20365),
	.b(n18099),
	.c(n20364));
   ao22f06 U24430 (.o(n20386),
	.a(n20373),
	.b(n20372),
	.c(n20371),
	.d(n20370));
   ao12f02 U24431 (.o(n20380),
	.a(n20377),
	.b(n20379),
	.c(n20378));
   no03m02 U24432 (.o(n20399),
	.a(n20389),
	.b(n20388),
	.c(n20387));
   oa12m02 U24433 (.o(n20398),
	.a(n20395),
	.b(n20397),
	.c(n20396));
   no02f03 U24434 (.o(n20405),
	.a(n20402),
	.b(n20401));
   no02f08 U24435 (.o(n20412),
	.a(n23035),
	.b(n25009));
   no02f04 U24436 (.o(n20455),
	.a(n17755),
	.b(FE_RN_23));
   no02s02 U24437 (.o(n20416),
	.a(n20415),
	.b(n20414));
   na02f01 U24438 (.o(n25154),
	.a(n20424),
	.b(n20423));
   no02f04 U24439 (.o(n20454),
	.a(FE_OFN94_n21695),
	.b(FE_OCPN25831_n20535));
   no02f10 U24440 (.o(n20534),
	.a(n20428),
	.b(n21907));
   oa12m02 U24441 (.o(n20436),
	.a(n20433),
	.b(n20435),
	.c(n20434));
   ao12f02 U24442 (.o(n20441),
	.a(n20438),
	.b(n20440),
	.c(n20439));
   na04f04 U24443 (.o(n20457),
	.a(n25180),
	.b(n25170),
	.c(n25496),
	.d(n25172));
   in01s01 U24444 (.o(n20494),
	.a(south_output_space_count_f_2_));
   in01s01 U24445 (.o(n20480),
	.a(south_output_space_valid_f));
   in01s01 U24446 (.o(n20492),
	.a(south_output_space_count_f_0_));
   no02f01 U24447 (.o(n20496),
	.a(n20491),
	.b(n20492));
   na02s01 U24448 (.o(n20481),
	.a(n20494),
	.b(n20489));
   in01s01 U24449 (.o(n20497),
	.a(n20493));
   no02m01 U24450 (.o(n20495),
	.a(south_output_space_count_f_0_),
	.b(south_output_space_count_f_1_));
   na02s01 U24451 (.o(n20486),
	.a(n20497),
	.b(n20495));
   in01s01 U24452 (.o(n20490),
	.a(south_output_space_N44));
   in01s01 U24453 (.o(n20485),
	.a(n20496));
   na02s01 U24454 (.o(n20488),
	.a(n20485),
	.b(n20484));
   no02f08 U24455 (.o(n25998),
	.a(n20529),
	.b(n20513));
   na02s01 U24456 (.o(n20511),
	.a(east_input_NIB_elements_in_array_f_1_),
	.b(n25315));
   in01f04 U24457 (.o(n25339),
	.a(n25997));
   na02f02 U24458 (.o(n20521),
	.a(n20520),
	.b(n20519));
   no02f02 U24459 (.o(n2438),
	.a(n20527),
	.b(n20526));
   no02f02 U24460 (.o(n25183),
	.a(FE_RN_23),
	.b(FE_OFN393_n19446));
   no02f04 U24461 (.o(n25174),
	.a(FE_OFN526_n24731),
	.b(n25175));
   in01s01 U24462 (.o(n20549),
	.a(east_output_control_planned_f));
   in01s01 U24463 (.o(n20752),
	.a(south_input_control_count_f_0_));
   na02s02 U24464 (.o(n23550),
	.a(n20563),
	.b(n22912));
   ao12s01 U24465 (.o(n20567),
	.a(n20630),
	.b(west_input_control_count_f_0_),
	.c(n20566));
   no02s01 U24466 (.o(n20568),
	.a(FE_OFN24831_n25232),
	.b(n20567));
   no02f01 U24467 (.o(n26012),
	.a(reset),
	.b(n20569));
   na02f01 U24468 (.o(n21886),
	.a(north_input_control_thanks_all_f),
	.b(n20737));
   in01s01 U24469 (.o(n20719),
	.a(north_input_control_count_f_0_));
   na02m01 U24470 (.o(n21887),
	.a(n20648),
	.b(n20737));
   na02f01 U24471 (.o(n20571),
	.a(n25433),
	.b(n20570));
   in01s01 U24472 (.o(n20573),
	.a(east_input_control_count_f_0_));
   ao22f01 U24473 (.o(n20575),
	.a(east_input_control_thanks_all_f),
	.b(n20573),
	.c(east_input_control_count_f_0_),
	.d(n21151));
   no02f01 U24474 (.o(n21565),
	.a(FE_OFN5_reset),
	.b(FE_OFN100_n21907));
   no02f01 U24475 (.o(n21657),
	.a(proc_input_control_count_f_0_),
	.b(n21688));
   ao12f01 U24476 (.o(n20576),
	.a(n21657),
	.b(proc_input_control_count_f_0_),
	.c(n21688));
   na02f02 U24477 (.o(n21689),
	.a(FE_OFN571_n25463),
	.b(FE_OFN947_n25096));
   na02f02 U24478 (.o(n21694),
	.a(FE_OFN428_n22902),
	.b(FE_OFN571_n25463));
   in01s01 U24479 (.o(n20577),
	.a(myLocY_4_));
   no02f01 U24480 (.o(N8),
	.a(FE_OFN25647_reset),
	.b(n20577));
   in01s01 U24481 (.o(n20578),
	.a(myLocY_0_));
   no02f01 U24482 (.o(N4),
	.a(FE_OFN25647_reset),
	.b(n20578));
   in01s01 U24483 (.o(n20579),
	.a(yummyIn_N));
   no02f01 U24484 (.o(north_output_space_N45),
	.a(FE_OFN25601_reset),
	.b(n20579));
   in01s01 U24485 (.o(n20580),
	.a(myChipID_11_));
   no02f01 U24486 (.o(N31),
	.a(FE_OFN25647_reset),
	.b(n20580));
   in01s01 U24487 (.o(n20581),
	.a(myLocX_4_));
   no02f01 U24488 (.o(N16),
	.a(FE_OFN25647_reset),
	.b(n20581));
   in01s01 U24489 (.o(n20582),
	.a(myLocX_6_));
   no02f01 U24490 (.o(N18),
	.a(FE_OFN25647_reset),
	.b(n20582));
   in01s01 U24491 (.o(n20583),
	.a(myLocX_0_));
   no02f01 U24492 (.o(N12),
	.a(FE_OFN8_reset),
	.b(n20583));
   in01s01 U24493 (.o(n20584),
	.a(myChipID_12_));
   no02f01 U24494 (.o(N32),
	.a(FE_OFN25647_reset),
	.b(n20584));
   in01s01 U24495 (.o(n20585),
	.a(myLocY_5_));
   no02f01 U24496 (.o(N9),
	.a(FE_OFN5_reset),
	.b(n20585));
   in01s01 U24497 (.o(n20586),
	.a(myChipID_9_));
   no02f01 U24498 (.o(N29),
	.a(FE_OFN25647_reset),
	.b(n20586));
   in01s01 U24499 (.o(n20587),
	.a(myChipID_2_));
   no02f01 U24500 (.o(N22),
	.a(FE_OFN25647_reset),
	.b(n20587));
   in01s01 U24501 (.o(n20588),
	.a(yummyIn_W));
   no02f01 U24502 (.o(west_output_space_N45),
	.a(FE_OFN25601_reset),
	.b(n20588));
   na02s01 U24503 (.o(west_input_control_N49),
	.a(FE_OFN25598_reset),
	.b(n20589));
   no02f01 U24504 (.o(n20591),
	.a(FE_OFN5_reset),
	.b(n20590));
   in01s01 U24505 (.o(south_input_control_N49),
	.a(n20591));
   in01s01 U24506 (.o(n20592),
	.a(myChipID_1_));
   no02f01 U24507 (.o(N21),
	.a(FE_OFN25647_reset),
	.b(n20592));
   in01s01 U24508 (.o(n20593),
	.a(myChipID_0_));
   no02f01 U24509 (.o(N20),
	.a(FE_OFN25647_reset),
	.b(n20593));
   in01s01 U24510 (.o(n20594),
	.a(myChipID_8_));
   no02f01 U24511 (.o(N28),
	.a(FE_OFN25647_reset),
	.b(n20594));
   in01s01 U24512 (.o(n20595),
	.a(myLocY_7_));
   no02f01 U24513 (.o(N11),
	.a(FE_OFN5_reset),
	.b(n20595));
   in01s01 U24514 (.o(n20596),
	.a(myLocX_7_));
   no02f01 U24515 (.o(N19),
	.a(FE_OFN25647_reset),
	.b(n20596));
   in01s01 U24516 (.o(n20597),
	.a(yummyIn_S));
   no02f01 U24517 (.o(south_output_space_N45),
	.a(reset),
	.b(n20597));
   in01s01 U24518 (.o(n20598),
	.a(myLocX_2_));
   no02f01 U24519 (.o(N14),
	.a(FE_OFN8_reset),
	.b(n20598));
   in01s01 U24520 (.o(n20599),
	.a(myChipID_3_));
   no02f01 U24521 (.o(N23),
	.a(FE_OFN25647_reset),
	.b(n20599));
   in01s01 U24522 (.o(n20600),
	.a(myLocX_3_));
   no02f01 U24523 (.o(N15),
	.a(reset),
	.b(n20600));
   in01s01 U24524 (.o(n20601),
	.a(myLocX_5_));
   no02f01 U24525 (.o(N17),
	.a(FE_OFN5_reset),
	.b(n20601));
   in01s01 U24526 (.o(n20602),
	.a(yummyIn_E));
   no02f01 U24527 (.o(east_output_space_N45),
	.a(FE_OFN25601_reset),
	.b(n20602));
   in01s01 U24528 (.o(n20603),
	.a(myLocX_1_));
   no02f01 U24529 (.o(N13),
	.a(FE_OFN25647_reset),
	.b(n20603));
   in01s01 U24530 (.o(n20604),
	.a(myChipID_6_));
   no02f01 U24531 (.o(N26),
	.a(FE_OFN25647_reset),
	.b(n20604));
   no02f01 U24532 (.o(N33),
	.a(FE_OFN25647_reset),
	.b(n20605));
   in01s01 U24533 (.o(n20606),
	.a(myChipID_7_));
   no02f01 U24534 (.o(N27),
	.a(FE_OFN25647_reset),
	.b(n20606));
   in01s01 U24535 (.o(n20607),
	.a(myChipID_4_));
   no02f01 U24536 (.o(N24),
	.a(FE_OFN25647_reset),
	.b(n20607));
   no02f01 U24537 (.o(N10),
	.a(FE_OFN5_reset),
	.b(n20608));
   in01s01 U24538 (.o(n20609),
	.a(myChipID_5_));
   no02f01 U24539 (.o(N25),
	.a(FE_OFN25647_reset),
	.b(n20609));
   in01s01 U24540 (.o(n20610),
	.a(myLocY_2_));
   no02f01 U24541 (.o(N6),
	.a(FE_OFN25647_reset),
	.b(n20610));
   in01s01 U24542 (.o(n20611),
	.a(myLocY_1_));
   no02f01 U24543 (.o(N5),
	.a(FE_OFN25647_reset),
	.b(n20611));
   in01s01 U24544 (.o(n20612),
	.a(myLocY_3_));
   no02f01 U24545 (.o(N7),
	.a(FE_OFN25647_reset),
	.b(n20612));
   in01s01 U24546 (.o(n20613),
	.a(myChipID_10_));
   no02f01 U24547 (.o(N30),
	.a(FE_OFN25647_reset),
	.b(n20613));
   in01s01 U24548 (.o(n20614),
	.a(yummyIn_P));
   no02f01 U24549 (.o(proc_output_space_N45),
	.a(reset),
	.b(n20614));
   in01s01 U24550 (.o(n20629),
	.a(west_input_control_count_f_1_));
   in01s01 U24551 (.o(n20615),
	.a(n20630));
   no03f01 U24552 (.o(west_input_control_N42),
	.a(FE_OFN25647_reset),
	.b(n21538),
	.c(n20617));
   no02f01 U24553 (.o(n20619),
	.a(FE_OFN5_reset),
	.b(n20618));
   in01s01 U24554 (.o(north_input_control_N49),
	.a(n20619));
   no02f01 U24555 (.o(n20621),
	.a(FE_OFN8_reset),
	.b(n20620));
   in01s01 U24556 (.o(proc_input_control_N49),
	.a(n20621));
   no02f01 U24557 (.o(n20623),
	.a(FE_OFN5_reset),
	.b(n20622));
   in01s01 U24558 (.o(east_input_control_N49),
	.a(n20623));
   na02s01 U24559 (.o(n20625),
	.a(west_input_control_count_f_3_),
	.b(n20633));
   in01s01 U24560 (.o(n20626),
	.a(n20625));
   ao12f01 U24561 (.o(west_input_control_N44),
	.a(FE_OFN25647_reset),
	.b(n20628),
	.c(n20627));
   na02s01 U24562 (.o(n20631),
	.a(n20630),
	.b(n20629));
   na02s01 U24563 (.o(n20632),
	.a(west_input_control_count_f_2_),
	.b(n20631));
   no02f01 U24564 (.o(west_input_control_N43),
	.a(FE_OFN25647_reset),
	.b(n20635));
   na02s01 U24565 (.o(n21384),
	.a(south_input_control_thanks_all_f),
	.b(n21385));
   in01s01 U24566 (.o(n20637),
	.a(n21384));
   in01s01 U24567 (.o(n20636),
	.a(south_input_control_count_f_2_));
   ao22s01 U24568 (.o(n20638),
	.a(south_input_control_count_f_2_),
	.b(n20637),
	.c(n21384),
	.d(n20636));
   na02s01 U24569 (.o(n20639),
	.a(n20638),
	.b(n22912));
   no02s01 U24570 (.o(n20647),
	.a(n20646),
	.b(n20645));
   in01s01 U24571 (.o(n20698),
	.a(north_input_control_count_f_2_));
   na02s01 U24572 (.o(n20650),
	.a(n20699),
	.b(n20698));
   in01s01 U24573 (.o(n20651),
	.a(n20650));
   in01s01 U24574 (.o(n20649),
	.a(north_input_control_count_f_3_));
   ao22s01 U24575 (.o(n20652),
	.a(north_input_control_count_f_3_),
	.b(n20651),
	.c(n20650),
	.d(n20649));
   na02s01 U24576 (.o(n20653),
	.a(n20652),
	.b(n20737));
   ao12f01 U24577 (.o(north_input_control_N44),
	.a(FE_OFN5_reset),
	.b(n20654),
	.c(n20653));
   na02f01 U24578 (.o(n20655),
	.a(north_input_NIB_tail_ptr_f_1_),
	.b(n25826));
   in01s01 U24579 (.o(n21277),
	.a(dataIn_N_56_));
   na02f01 U24580 (.o(n20657),
	.a(north_input_NIB_storage_data_f_2__56_),
	.b(FE_OFN25876_n25842));
   in01s01 U24581 (.o(n21280),
	.a(dataIn_N_52_));
   na02f01 U24582 (.o(n20658),
	.a(north_input_NIB_storage_data_f_2__52_),
	.b(FE_OFN25876_n25842));
   in01s01 U24583 (.o(n21274),
	.a(dataIn_N_57_));
   na02f01 U24584 (.o(n20659),
	.a(north_input_NIB_storage_data_f_2__57_),
	.b(FE_OFN25876_n25842));
   in01s01 U24585 (.o(n22630),
	.a(dataIn_N_43_));
   na02f01 U24586 (.o(n20660),
	.a(north_input_NIB_storage_data_f_2__43_),
	.b(FE_OFN1087_n20656));
   in01s01 U24587 (.o(n21282),
	.a(dataIn_N_50_));
   na02f01 U24588 (.o(n20661),
	.a(north_input_NIB_storage_data_f_2__50_),
	.b(FE_OFN1087_n20656));
   in01s01 U24589 (.o(n22636),
	.a(dataIn_N_46_));
   na02f01 U24590 (.o(n20662),
	.a(north_input_NIB_storage_data_f_2__46_),
	.b(FE_OFN1087_n20656));
   in01s01 U24591 (.o(n21254),
	.a(dataIn_N_55_));
   na02f01 U24592 (.o(n20663),
	.a(north_input_NIB_storage_data_f_2__55_),
	.b(FE_OFN25876_n25842));
   in01s01 U24593 (.o(n22646),
	.a(dataIn_N_39_));
   na02f01 U24594 (.o(n20664),
	.a(north_input_NIB_storage_data_f_2__39_),
	.b(FE_OFN1087_n20656));
   in01s01 U24595 (.o(n21270),
	.a(dataIn_N_54_));
   na02f01 U24596 (.o(n20665),
	.a(north_input_NIB_storage_data_f_2__54_),
	.b(FE_OFN25876_n25842));
   in01s01 U24597 (.o(n21248),
	.a(dataIn_N_29_));
   na02f01 U24598 (.o(n20667),
	.a(north_input_NIB_storage_data_f_2__49_),
	.b(FE_OFN1087_n20656));
   in01s01 U24599 (.o(n21264),
	.a(dataIn_N_41_));
   na02f01 U24600 (.o(n20668),
	.a(north_input_NIB_storage_data_f_2__41_),
	.b(FE_OFN1087_n20656));
   in01s01 U24601 (.o(n22654),
	.a(dataIn_N_37_));
   na02f01 U24602 (.o(n20669),
	.a(north_input_NIB_storage_data_f_2__37_),
	.b(FE_OFN1087_n20656));
   in01s01 U24603 (.o(n21256),
	.a(dataIn_N_58_));
   na02f01 U24604 (.o(n20670),
	.a(north_input_NIB_storage_data_f_2__58_),
	.b(FE_OFN25876_n25842));
   in01s01 U24605 (.o(n21232),
	.a(dataIn_N_25_));
   na02f01 U24606 (.o(n20671),
	.a(north_input_NIB_storage_data_f_2__25_),
	.b(FE_OFN1087_n20656));
   in01s01 U24607 (.o(n22656),
	.a(dataIn_N_36_));
   na02f01 U24608 (.o(n20672),
	.a(north_input_NIB_storage_data_f_2__36_),
	.b(FE_OFN1087_n20656));
   in01s01 U24609 (.o(n22644),
	.a(dataIn_N_35_));
   na02f01 U24610 (.o(n20673),
	.a(north_input_NIB_storage_data_f_2__35_),
	.b(FE_OFN1087_n20656));
   in01s01 U24611 (.o(n21272),
	.a(dataIn_N_44_));
   na02f01 U24612 (.o(n20675),
	.a(north_input_NIB_storage_data_f_2__34_),
	.b(FE_OFN1087_n20656));
   in01s01 U24613 (.o(n22650),
	.a(dataIn_N_42_));
   na02f01 U24614 (.o(n20676),
	.a(north_input_NIB_storage_data_f_2__42_),
	.b(FE_OFN1087_n20656));
   in01s01 U24615 (.o(n21239),
	.a(dataIn_N_51_));
   na02f01 U24616 (.o(n20677),
	.a(north_input_NIB_storage_data_f_2__51_),
	.b(FE_OFN25876_n25842));
   in01s01 U24617 (.o(n22640),
	.a(dataIn_N_32_));
   na02f01 U24618 (.o(n20678),
	.a(north_input_NIB_storage_data_f_2__32_),
	.b(FE_OFN1087_n20656));
   in01s01 U24619 (.o(n21237),
	.a(dataIn_N_31_));
   na02f01 U24620 (.o(n20679),
	.a(north_input_NIB_storage_data_f_2__31_),
	.b(FE_OFN1087_n20656));
   in01s01 U24621 (.o(n22638),
	.a(dataIn_N_38_));
   na02f01 U24622 (.o(n20680),
	.a(north_input_NIB_storage_data_f_2__38_),
	.b(FE_OFN1087_n20656));
   in01s01 U24623 (.o(n22444),
	.a(dataIn_N_61_));
   na02f01 U24624 (.o(n20681),
	.a(north_input_NIB_storage_data_f_2__61_),
	.b(FE_OFN25876_n25842));
   in01s01 U24625 (.o(n21243),
	.a(dataIn_N_28_));
   na02f01 U24626 (.o(n20682),
	.a(north_input_NIB_storage_data_f_2__28_),
	.b(FE_OFN1087_n20656));
   in01s01 U24627 (.o(n21250),
	.a(dataIn_N_27_));
   na02f01 U24628 (.o(n20683),
	.a(north_input_NIB_storage_data_f_2__27_),
	.b(FE_OFN1087_n20656));
   na02f01 U24629 (.o(n20684),
	.a(north_input_NIB_storage_data_f_2__26_),
	.b(FE_OFN1087_n20656));
   in01s01 U24630 (.o(n21241),
	.a(dataIn_N_63_));
   na02f01 U24631 (.o(n20685),
	.a(north_input_NIB_storage_data_f_2__63_),
	.b(FE_OFN25876_n25842));
   in01s01 U24632 (.o(n22642),
	.a(dataIn_N_59_));
   in01s01 U24633 (.o(n22632),
	.a(dataIn_N_45_));
   na02f01 U24634 (.o(n20687),
	.a(north_input_NIB_storage_data_f_2__45_),
	.b(FE_OFN1087_n20656));
   in01s01 U24635 (.o(n22652),
	.a(dataIn_N_48_));
   na02f01 U24636 (.o(n20688),
	.a(north_input_NIB_storage_data_f_2__48_),
	.b(FE_OFN1087_n20656));
   in01s01 U24637 (.o(n21234),
	.a(dataIn_N_47_));
   na02f01 U24638 (.o(n20689),
	.a(north_input_NIB_storage_data_f_2__47_),
	.b(FE_OFN1087_n20656));
   in01s01 U24639 (.o(n21226),
	.a(dataIn_N_22_));
   na02f01 U24640 (.o(n20690),
	.a(north_input_NIB_storage_data_f_2__22_),
	.b(FE_OFN1087_n20656));
   in01s01 U24641 (.o(n21246),
	.a(dataIn_N_62_));
   na02f01 U24642 (.o(n20691),
	.a(north_input_NIB_storage_data_f_2__62_),
	.b(FE_OFN25876_n25842));
   in01s01 U24643 (.o(n21262),
	.a(dataIn_N_40_));
   na02f01 U24644 (.o(n20692),
	.a(north_input_NIB_storage_data_f_2__40_),
	.b(FE_OFN1087_n20656));
   in01s01 U24645 (.o(n21259),
	.a(dataIn_N_30_));
   na02f01 U24646 (.o(n20693),
	.a(north_input_NIB_storage_data_f_2__30_),
	.b(FE_OFN1087_n20656));
   in01s01 U24647 (.o(n21224),
	.a(dataIn_N_24_));
   na02f01 U24648 (.o(n20694),
	.a(north_input_NIB_storage_data_f_2__24_),
	.b(FE_OFN1087_n20656));
   in01s01 U24649 (.o(n21222),
	.a(dataIn_N_23_));
   na02f01 U24650 (.o(n20695),
	.a(north_input_NIB_storage_data_f_2__23_),
	.b(FE_OFN1087_n20656));
   in01s01 U24651 (.o(n21287),
	.a(dataIn_N_60_));
   na02f01 U24652 (.o(n20696),
	.a(north_input_NIB_storage_data_f_2__60_),
	.b(FE_OFN25876_n25842));
   in01s01 U24653 (.o(n21285),
	.a(dataIn_N_53_));
   na02f01 U24654 (.o(n20697),
	.a(north_input_NIB_storage_data_f_2__53_),
	.b(FE_OFN1087_n20656));
   in01s01 U24655 (.o(n20702),
	.a(n24031));
   na02s02 U24656 (.o(n20724),
	.a(n21893),
	.b(n25433));
   in01s01 U24657 (.o(n20700),
	.a(n20699));
   ao22s01 U24658 (.o(n20701),
	.a(north_input_control_count_f_2_),
	.b(n20700),
	.c(FE_OFN25845_n20699),
	.d(n20698));
   oa22s01 U24659 (.o(north_input_control_N43),
	.a(n20702),
	.b(n20724),
	.c(n20701),
	.d(n20711));
   in01s01 U24660 (.o(n20706),
	.a(n23949));
   in01s01 U24661 (.o(n20723),
	.a(n21887));
   in01s01 U24662 (.o(n20722),
	.a(n21886));
   no02f01 U24663 (.o(n21888),
	.a(north_input_control_count_f_2_),
	.b(north_input_control_count_f_3_));
   na02f02 U24664 (.o(n20734),
	.a(n21888),
	.b(n20703));
   oa22f01 U24665 (.o(north_input_control_N47),
	.a(n20706),
	.b(n20724),
	.c(FE_OFN5_reset),
	.d(n21896));
   in01s01 U24666 (.o(n20713),
	.a(n23957));
   na02s01 U24667 (.o(n20740),
	.a(north_input_control_thanks_all_f),
	.b(n20707));
   no02m01 U24668 (.o(n20709),
	.a(north_input_control_count_f_6_),
	.b(n20740));
   in01s01 U24669 (.o(n20708),
	.a(north_input_control_count_f_7_));
   ao22m01 U24670 (.o(n20712),
	.a(north_input_control_count_f_7_),
	.b(n20710),
	.c(n20709),
	.d(n20708));
   oa22m01 U24671 (.o(north_input_control_N48),
	.a(n20713),
	.b(n20724),
	.c(n20712),
	.d(n20711));
   in01s01 U24672 (.o(n20718),
	.a(n23524));
   in01s01 U24673 (.o(n20716),
	.a(north_input_control_count_f_4_));
   na02s01 U24674 (.o(n20714),
	.a(n20734),
	.b(n20716));
   oa12s01 U24675 (.o(n20715),
	.a(n20714),
	.b(n20716),
	.c(n20734));
   in01s01 U24676 (.o(n20717),
	.a(n21890));
   oa22f01 U24677 (.o(north_input_control_N45),
	.a(n20718),
	.b(n20724),
	.c(FE_OFN5_reset),
	.d(n20717));
   in01s01 U24678 (.o(n20725),
	.a(n23620));
   in01s01 U24679 (.o(n20720),
	.a(north_input_control_count_f_1_));
   ao22s01 U24680 (.o(n20721),
	.a(north_input_control_count_f_0_),
	.b(n20720),
	.c(north_input_control_count_f_1_),
	.d(n20719));
   oa22f01 U24681 (.o(north_input_control_N42),
	.a(n20725),
	.b(n20724),
	.c(FE_OFN5_reset),
	.d(n21897));
   na02s01 U24682 (.o(n20729),
	.a(n24970),
	.b(n20728));
   no02f01 U24683 (.o(n20733),
	.a(n20732),
	.b(n20731));
   no02s01 U24684 (.o(n20735),
	.a(north_input_control_count_f_4_),
	.b(n20734));
   ao12s01 U24685 (.o(north_input_control_N46),
	.a(n20738),
	.b(n20740),
	.c(n20739));
   na02f01 U24686 (.o(n20743),
	.a(n20742),
	.b(n20741));
   in01f01 U24687 (.o(n20744),
	.a(n20743));
   in01s01 U24688 (.o(n20754),
	.a(south_input_control_count_f_1_));
   oa22s01 U24689 (.o(n25238),
	.a(south_input_control_count_f_0_),
	.b(n20754),
	.c(south_input_control_count_f_1_),
	.d(n20752));
   no02s01 U24690 (.o(n20757),
	.a(n25250),
	.b(n25238));
   no02s01 U24692 (.o(n20755),
	.a(n23550),
	.b(n20754));
   no02f01 U24693 (.o(south_input_control_N42),
	.a(FE_OFN5_reset),
	.b(n20758));
   no02f01 U24694 (.o(n20762),
	.a(n20761),
	.b(n20760));
   no02f01 U24695 (.o(n20765),
	.a(n20764),
	.b(n20763));
   in01f02 U24696 (.o(n23527),
	.a(n20766));
   na02f01 U24697 (.o(n20773),
	.a(n20767),
	.b(n23527));
   no02s01 U24698 (.o(n20769),
	.a(east_input_control_count_f_3_),
	.b(east_input_control_count_f_2_));
   na02s01 U24699 (.o(n20770),
	.a(n21584),
	.b(n20769));
   in01s01 U24700 (.o(n21577),
	.a(n20770));
   in01s01 U24701 (.o(n21576),
	.a(east_input_control_count_f_4_));
   ao12f01 U24702 (.o(east_input_control_N45),
	.a(FE_OFN5_reset),
	.b(n20773),
	.c(n20772));
   na02f01 U24703 (.o(n20776),
	.a(n20775),
	.b(n20774));
   in01s01 U24704 (.o(n20777),
	.a(n20776));
   no02f01 U24705 (.o(n20780),
	.a(n20779),
	.b(n20778));
   no02f01 U24706 (.o(n20783),
	.a(n20782),
	.b(n20781));
   no02f02 U24707 (.o(n20787),
	.a(n20786),
	.b(n20785));
   no02f02 U24708 (.o(n20790),
	.a(n20789),
	.b(n20788));
   in01s01 U24709 (.o(n25896),
	.a(south_input_NIB_tail_ptr_f_0_));
   no02f01 U24710 (.o(n20795),
	.a(south_input_NIB_tail_ptr_f_1_),
	.b(n25896));
   in01s01 U24711 (.o(n21024),
	.a(dataIn_S_30_));
   na02f01 U24712 (.o(n20798),
	.a(south_input_NIB_storage_data_f_1__30_),
	.b(FE_OFN25785_n17770));
   oa12s01 U24713 (.o(n10008),
	.a(n20798),
	.b(FE_OFN25785_n17770),
	.c(n21024));
   in01s01 U24714 (.o(n21005),
	.a(dataIn_S_27_));
   na02s01 U24715 (.o(n20799),
	.a(south_input_NIB_storage_data_f_1__27_),
	.b(FE_OFN25785_n17770));
   oa12s01 U24716 (.o(n10023),
	.a(n20799),
	.b(FE_OFN25785_n17770),
	.c(n21005));
   in01s01 U24717 (.o(n21030),
	.a(dataIn_S_28_));
   na02s01 U24718 (.o(n20800),
	.a(south_input_NIB_storage_data_f_1__28_),
	.b(FE_OFN25785_n17770));
   in01s01 U24719 (.o(n21007),
	.a(dataIn_S_62_));
   na02m01 U24720 (.o(n20801),
	.a(south_input_NIB_storage_data_f_1__62_),
	.b(FE_OFN25853_FE_OFN899_n17770));
   oa12s01 U24721 (.o(n9848),
	.a(n20801),
	.b(FE_OFN25853_FE_OFN899_n17770),
	.c(n21007));
   in01s01 U24722 (.o(n22679),
	.a(dataIn_S_48_));
   na02s01 U24723 (.o(n20802),
	.a(south_input_NIB_storage_data_f_1__48_),
	.b(FE_OFN25785_n17770));
   oa12s01 U24724 (.o(n9918),
	.a(n20802),
	.b(FE_OFN25785_n17770),
	.c(n22679));
   in01s01 U24725 (.o(n21009),
	.a(dataIn_S_25_));
   na02f02 U24726 (.o(n20803),
	.a(south_input_NIB_storage_data_f_1__25_),
	.b(FE_OFN25785_n17770));
   oa12s01 U24727 (.o(n10033),
	.a(n20803),
	.b(FE_OFN25785_n17770),
	.c(n21009));
   in01s01 U24728 (.o(n21035),
	.a(dataIn_S_50_));
   na02m01 U24729 (.o(n20804),
	.a(south_input_NIB_storage_data_f_1__50_),
	.b(FE_OFN25850_FE_OFN899_n17770));
   oa12f01 U24730 (.o(n9908),
	.a(n20804),
	.b(FE_OFN25850_FE_OFN899_n17770),
	.c(n21035));
   in01s01 U24731 (.o(n21040),
	.a(dataIn_S_54_));
   na02m01 U24732 (.o(n20805),
	.a(south_input_NIB_storage_data_f_1__54_),
	.b(FE_OFN25857_FE_OFN899_n17770));
   oa12s01 U24733 (.o(n9888),
	.a(n20805),
	.b(FE_OFN25857_FE_OFN899_n17770),
	.c(n21040));
   in01s01 U24734 (.o(n21014),
	.a(dataIn_S_55_));
   na02m01 U24735 (.o(n20806),
	.a(south_input_NIB_storage_data_f_1__55_),
	.b(FE_OFN25857_FE_OFN899_n17770));
   oa12s01 U24736 (.o(n9883),
	.a(n20806),
	.b(FE_OFN25857_FE_OFN899_n17770),
	.c(n21014));
   in01s01 U24737 (.o(n21049),
	.a(dataIn_S_29_));
   na02s01 U24738 (.o(n20807),
	.a(south_input_NIB_storage_data_f_1__29_),
	.b(FE_OFN25785_n17770));
   oa12s01 U24739 (.o(n10013),
	.a(n20807),
	.b(FE_OFN25785_n17770),
	.c(n21049));
   in01s01 U24740 (.o(n21026),
	.a(dataIn_S_57_));
   na02m01 U24741 (.o(n20808),
	.a(south_input_NIB_storage_data_f_1__57_),
	.b(FE_OFN25849_FE_OFN899_n17770));
   oa12s01 U24742 (.o(n9873),
	.a(n20808),
	.b(FE_OFN25849_FE_OFN899_n17770),
	.c(n21026));
   in01f01 U24743 (.o(n21044),
	.a(dataIn_S_24_));
   na02s01 U24744 (.o(n20809),
	.a(south_input_NIB_storage_data_f_1__24_),
	.b(FE_OFN25785_n17770));
   oa12s01 U24745 (.o(n10038),
	.a(n20809),
	.b(FE_OFN25785_n17770),
	.c(n21044));
   in01s01 U24746 (.o(n21018),
	.a(dataIn_S_59_));
   na02m01 U24747 (.o(n20810),
	.a(south_input_NIB_storage_data_f_1__59_),
	.b(FE_OFN25850_FE_OFN899_n17770));
   oa12f01 U24748 (.o(n9863),
	.a(n20810),
	.b(FE_OFN25850_FE_OFN899_n17770),
	.c(n21018));
   in01s01 U24749 (.o(n21020),
	.a(dataIn_S_40_));
   na02s01 U24750 (.o(n20811),
	.a(south_input_NIB_storage_data_f_1__40_),
	.b(FE_OFN899_n17770));
   oa12s01 U24751 (.o(n9958),
	.a(n20811),
	.b(FE_OFN899_n17770),
	.c(n21020));
   in01s01 U24752 (.o(n21012),
	.a(dataIn_S_61_));
   na02m01 U24753 (.o(n20812),
	.a(south_input_NIB_storage_data_f_1__61_),
	.b(FE_OFN25857_FE_OFN899_n17770));
   oa12s01 U24754 (.o(n9853),
	.a(n20812),
	.b(FE_OFN25857_FE_OFN899_n17770),
	.c(n21012));
   no02f01 U24755 (.o(n20813),
	.a(south_input_NIB_tail_ptr_f_0_),
	.b(south_input_NIB_tail_ptr_f_1_));
   in01s01 U24756 (.o(n21037),
	.a(dataIn_S_56_));
   na02s01 U24757 (.o(n20816),
	.a(south_input_NIB_storage_data_f_0__56_),
	.b(FE_OFN403_n20815));
   oa12s01 U24758 (.o(n9558),
	.a(n20816),
	.b(FE_OFN403_n20815),
	.c(n21037));
   in01s01 U24759 (.o(n22690),
	.a(dataIn_S_38_));
   na02f01 U24760 (.o(n20817),
	.a(south_input_NIB_storage_data_f_1__38_),
	.b(FE_OFN25785_n17770));
   oa12s01 U24761 (.o(n9968),
	.a(n20817),
	.b(FE_OFN25785_n17770),
	.c(n22690));
   in01s01 U24762 (.o(n21028),
	.a(dataIn_S_22_));
   na02s01 U24763 (.o(n20818),
	.a(south_input_NIB_storage_data_f_0__22_),
	.b(FE_OFN952_n25916));
   oa12s01 U24764 (.o(n9728),
	.a(n20818),
	.b(FE_OFN952_n25916),
	.c(n21028));
   in01s01 U24765 (.o(n22482),
	.a(dataIn_S_52_));
   na02m01 U24766 (.o(n20819),
	.a(south_input_NIB_storage_data_f_1__52_),
	.b(FE_OFN25854_FE_OFN899_n17770));
   oa12s01 U24767 (.o(n9898),
	.a(n20819),
	.b(FE_OFN25854_FE_OFN899_n17770),
	.c(n22482));
   in01s01 U24768 (.o(n21042),
	.a(dataIn_S_53_));
   na02m01 U24769 (.o(n20820),
	.a(south_input_NIB_storage_data_f_1__53_),
	.b(FE_OFN899_n17770));
   oa12s01 U24770 (.o(n9893),
	.a(n20820),
	.b(FE_OFN899_n17770),
	.c(n21042));
   in01s01 U24771 (.o(n21046),
	.a(dataIn_S_23_));
   na02f01 U24772 (.o(n20821),
	.a(south_input_NIB_storage_data_f_1__23_),
	.b(FE_OFN25785_n17770));
   oa12s01 U24773 (.o(n10043),
	.a(n20821),
	.b(FE_OFN25785_n17770),
	.c(n21046));
   na02s01 U24774 (.o(n20822),
	.a(south_input_NIB_storage_data_f_0__23_),
	.b(FE_OFN952_n25916));
   oa12s01 U24775 (.o(n9723),
	.a(n20822),
	.b(FE_OFN952_n25916),
	.c(n21046));
   na02s01 U24776 (.o(n20823),
	.a(south_input_NIB_storage_data_f_0__24_),
	.b(FE_OFN952_n25916));
   in01f01 U24777 (.o(n21032),
	.a(dataIn_S_26_));
   na02f01 U24778 (.o(n20824),
	.a(south_input_NIB_storage_data_f_1__26_),
	.b(FE_OFN25785_n17770));
   oa12s01 U24779 (.o(n10028),
	.a(n20824),
	.b(FE_OFN25785_n17770),
	.c(n21032));
   na02s01 U24780 (.o(n20825),
	.a(south_input_NIB_storage_data_f_0__25_),
	.b(FE_OFN952_n25916));
   oa12s01 U24781 (.o(n9713),
	.a(n20825),
	.b(FE_OFN952_n25916),
	.c(n21009));
   na02s01 U24782 (.o(n20826),
	.a(south_input_NIB_storage_data_f_0__26_),
	.b(FE_OFN952_n25916));
   oa12s01 U24783 (.o(n9708),
	.a(n20826),
	.b(FE_OFN952_n25916),
	.c(n21032));
   na02s01 U24784 (.o(n20827),
	.a(south_input_NIB_storage_data_f_0__27_),
	.b(FE_OFN952_n25916));
   oa12s01 U24785 (.o(n9703),
	.a(n20827),
	.b(FE_OFN952_n25916),
	.c(n21005));
   na02s01 U24786 (.o(n20828),
	.a(south_input_NIB_storage_data_f_0__28_),
	.b(FE_OFN952_n25916));
   oa12s01 U24787 (.o(n9698),
	.a(n20828),
	.b(FE_OFN952_n25916),
	.c(n21030));
   oa12s01 U24788 (.o(n9693),
	.a(n20829),
	.b(FE_OFN952_n25916),
	.c(n21049));
   na02s01 U24789 (.o(n20830),
	.a(south_input_NIB_storage_data_f_1__49_),
	.b(FE_OFN25785_n17770));
   oa12s01 U24790 (.o(n9913),
	.a(n20830),
	.b(FE_OFN25785_n17770),
	.c(n20998));
   na02s01 U24791 (.o(n20831),
	.a(south_input_NIB_storage_data_f_0__30_),
	.b(FE_OFN952_n25916));
   oa12s01 U24792 (.o(n9688),
	.a(n20831),
	.b(FE_OFN952_n25916),
	.c(n21024));
   in01s01 U24793 (.o(n22688),
	.a(dataIn_S_41_));
   na02s01 U24794 (.o(n20832),
	.a(south_input_NIB_storage_data_f_1__41_),
	.b(FE_OFN25785_n17770));
   oa12s01 U24795 (.o(n9953),
	.a(n20832),
	.b(FE_OFN25785_n17770),
	.c(n22688));
   na02s01 U24796 (.o(n20833),
	.a(south_input_NIB_storage_data_f_0__38_),
	.b(FE_OFN952_n25916));
   oa12s01 U24797 (.o(n9648),
	.a(n20833),
	.b(FE_OFN952_n25916),
	.c(n22690));
   na02s01 U24798 (.o(n20834),
	.a(south_input_NIB_storage_data_f_0__40_),
	.b(FE_OFN403_n20815));
   oa12s01 U24799 (.o(n9638),
	.a(n20834),
	.b(FE_OFN403_n20815),
	.c(n21020));
   na02s01 U24800 (.o(n20835),
	.a(south_input_NIB_storage_data_f_0__41_),
	.b(FE_OFN952_n25916));
   oa12s01 U24801 (.o(n9633),
	.a(n20835),
	.b(FE_OFN952_n25916),
	.c(n22688));
   na02s01 U24802 (.o(n20836),
	.a(south_input_NIB_storage_data_f_0__48_),
	.b(FE_OFN952_n25916));
   oa12s01 U24803 (.o(n9598),
	.a(n20836),
	.b(FE_OFN952_n25916),
	.c(n22679));
   na02s01 U24804 (.o(n20837),
	.a(south_input_NIB_storage_data_f_0__49_),
	.b(FE_OFN952_n25916));
   oa12s01 U24805 (.o(n9593),
	.a(n20837),
	.b(FE_OFN952_n25916),
	.c(n20998));
   na02s01 U24806 (.o(n20838),
	.a(south_input_NIB_storage_data_f_0__50_),
	.b(FE_OFN403_n20815));
   oa12s01 U24807 (.o(n9588),
	.a(n20838),
	.b(FE_OFN403_n20815),
	.c(n21035));
   na02s01 U24808 (.o(n20839),
	.a(south_input_NIB_storage_data_f_0__52_),
	.b(FE_OFN403_n20815));
   oa12s01 U24809 (.o(n9578),
	.a(n20839),
	.b(FE_OFN403_n20815),
	.c(n22482));
   na02m01 U24810 (.o(n20840),
	.a(south_input_NIB_storage_data_f_1__56_),
	.b(FE_OFN25855_FE_OFN899_n17770));
   oa12s01 U24811 (.o(n9878),
	.a(n20840),
	.b(FE_OFN25855_FE_OFN899_n17770),
	.c(n21037));
   na02s01 U24812 (.o(n20841),
	.a(south_input_NIB_storage_data_f_0__53_),
	.b(FE_OFN403_n20815));
   oa12s01 U24813 (.o(n9573),
	.a(n20841),
	.b(FE_OFN403_n20815),
	.c(n21042));
   in01s01 U24814 (.o(n21022),
	.a(dataIn_S_58_));
   na02m01 U24815 (.o(n20842),
	.a(south_input_NIB_storage_data_f_1__58_),
	.b(FE_OFN25857_FE_OFN899_n17770));
   na02s01 U24816 (.o(n20843),
	.a(south_input_NIB_storage_data_f_0__54_),
	.b(FE_OFN403_n20815));
   in01s01 U24817 (.o(n21016),
	.a(dataIn_S_60_));
   na02m01 U24818 (.o(n20844),
	.a(south_input_NIB_storage_data_f_1__60_),
	.b(FE_OFN25850_FE_OFN899_n17770));
   oa12f01 U24819 (.o(n9858),
	.a(n20844),
	.b(FE_OFN25850_FE_OFN899_n17770),
	.c(n21016));
   na02s01 U24820 (.o(n20845),
	.a(south_input_NIB_storage_data_f_0__55_),
	.b(FE_OFN403_n20815));
   oa12s01 U24821 (.o(n9563),
	.a(n20845),
	.b(FE_OFN403_n20815),
	.c(n21014));
   na02s01 U24822 (.o(n20846),
	.a(south_input_NIB_storage_data_f_0__60_),
	.b(FE_OFN403_n20815));
   oa12s01 U24823 (.o(n9538),
	.a(n20846),
	.b(FE_OFN403_n20815),
	.c(n21016));
   na02s01 U24824 (.o(n20847),
	.a(south_input_NIB_storage_data_f_0__57_),
	.b(FE_OFN403_n20815));
   oa12s01 U24825 (.o(n9553),
	.a(n20847),
	.b(FE_OFN403_n20815),
	.c(n21026));
   na02s01 U24826 (.o(n20848),
	.a(south_input_NIB_storage_data_f_0__58_),
	.b(FE_OFN403_n20815));
   oa12s01 U24827 (.o(n9548),
	.a(n20848),
	.b(FE_OFN403_n20815),
	.c(n21022));
   na02s01 U24828 (.o(n20849),
	.a(south_input_NIB_storage_data_f_0__59_),
	.b(FE_OFN403_n20815));
   oa12s01 U24829 (.o(n9543),
	.a(n20849),
	.b(FE_OFN403_n20815),
	.c(n21018));
   na02f01 U24830 (.o(n20850),
	.a(south_input_NIB_storage_data_f_1__22_),
	.b(FE_OFN25785_n17770));
   oa12s01 U24831 (.o(n10048),
	.a(n20850),
	.b(FE_OFN25785_n17770),
	.c(n21028));
   na02s01 U24832 (.o(n20851),
	.a(south_input_NIB_storage_data_f_0__62_),
	.b(FE_OFN403_n20815));
   oa12s01 U24833 (.o(n9528),
	.a(n20851),
	.b(FE_OFN403_n20815),
	.c(n21007));
   na02s01 U24834 (.o(n20852),
	.a(south_input_NIB_storage_data_f_0__61_),
	.b(FE_OFN403_n20815));
   oa12s01 U24835 (.o(n9533),
	.a(n20852),
	.b(FE_OFN403_n20815),
	.c(n21012));
   in01s01 U24836 (.o(n21072),
	.a(dataIn_W_63_));
   na02s01 U24837 (.o(n20856),
	.a(west_input_NIB_storage_data_f_0__63_),
	.b(FE_OFN25750_FE_OFN24796_n20854));
   oa12s01 U24838 (.o(n8233),
	.a(n20856),
	.b(FE_OFN25750_FE_OFN24796_n20854),
	.c(n21072));
   in01f01 U24839 (.o(n25928),
	.a(west_input_NIB_tail_ptr_f_0_));
   no02f01 U24840 (.o(n20857),
	.a(west_input_NIB_tail_ptr_f_1_),
	.b(n25928));
   in01s01 U24841 (.o(n21086),
	.a(dataIn_W_50_));
   na02s01 U24842 (.o(n20860),
	.a(west_input_NIB_storage_data_f_1__50_),
	.b(FE_OFN381_n17772));
   oa12f01 U24843 (.o(n8618),
	.a(n20860),
	.b(FE_OFN381_n17772),
	.c(n21086));
   in01s01 U24844 (.o(n21095),
	.a(dataIn_W_61_));
   na02f01 U24845 (.o(n20861),
	.a(west_input_NIB_storage_data_f_0__61_),
	.b(FE_OFN25748_FE_OFN24796_n20854));
   oa12f01 U24846 (.o(n8243),
	.a(n20861),
	.b(FE_OFN25748_FE_OFN24796_n20854),
	.c(n21095));
   in01s01 U24847 (.o(n21097),
	.a(dataIn_W_60_));
   na02s01 U24848 (.o(n20862),
	.a(west_input_NIB_storage_data_f_0__60_),
	.b(FE_OFN25750_FE_OFN24796_n20854));
   oa12s01 U24849 (.o(n8248),
	.a(n20862),
	.b(FE_OFN25750_FE_OFN24796_n20854),
	.c(n21097));
   in01s01 U24850 (.o(n22717),
	.a(dataIn_W_52_));
   na02s01 U24851 (.o(n20863),
	.a(west_input_NIB_storage_data_f_0__52_),
	.b(FE_OFN25750_FE_OFN24796_n20854));
   oa12s01 U24852 (.o(n8288),
	.a(n20863),
	.b(FE_OFN25750_FE_OFN24796_n20854),
	.c(n22717));
   in01s01 U24853 (.o(n21084),
	.a(dataIn_W_51_));
   na02s01 U24854 (.o(n20864),
	.a(west_input_NIB_storage_data_f_0__51_),
	.b(FE_OFN25750_FE_OFN24796_n20854));
   na02f01 U24855 (.o(n20865),
	.a(west_input_NIB_storage_data_f_0__50_),
	.b(FE_OFN25747_FE_OFN24796_n20854));
   oa12f01 U24856 (.o(n8298),
	.a(n20865),
	.b(FE_OFN25747_FE_OFN24796_n20854),
	.c(n21086));
   in01s01 U24857 (.o(n21091),
	.a(dataIn_W_49_));
   na02f01 U24858 (.o(n20866),
	.a(west_input_NIB_storage_data_f_0__49_),
	.b(FE_OFN25747_FE_OFN24796_n20854));
   oa12f01 U24859 (.o(n8303),
	.a(n20866),
	.b(FE_OFN25747_FE_OFN24796_n20854),
	.c(n21091));
   in01s01 U24860 (.o(n21099),
	.a(dataIn_W_48_));
   na02f01 U24861 (.o(n20867),
	.a(west_input_NIB_storage_data_f_0__48_),
	.b(FE_OFN25747_FE_OFN24796_n20854));
   oa12f01 U24862 (.o(n8308),
	.a(n20867),
	.b(FE_OFN25747_FE_OFN24796_n20854),
	.c(n21099));
   na02s01 U24863 (.o(n20868),
	.a(west_input_NIB_storage_data_f_0__47_),
	.b(FE_OFN25747_FE_OFN24796_n20854));
   oa12f01 U24864 (.o(n8313),
	.a(n20868),
	.b(FE_OFN25747_FE_OFN24796_n20854),
	.c(n21125));
   in01s01 U24865 (.o(n21101),
	.a(dataIn_W_45_));
   na02f01 U24866 (.o(n20869),
	.a(west_input_NIB_storage_data_f_0__45_),
	.b(FE_OFN25748_FE_OFN24796_n20854));
   oa12f01 U24867 (.o(n8323),
	.a(n20869),
	.b(FE_OFN25748_FE_OFN24796_n20854),
	.c(n21101));
   in01s01 U24868 (.o(n22486),
	.a(dataIn_W_44_));
   na02f01 U24869 (.o(n20870),
	.a(west_input_NIB_storage_data_f_0__44_),
	.b(FE_OFN25748_FE_OFN24796_n20854));
   oa12f01 U24870 (.o(n8328),
	.a(n20870),
	.b(FE_OFN25748_FE_OFN24796_n20854),
	.c(n22486));
   in01s01 U24871 (.o(n21129),
	.a(dataIn_W_43_));
   na02f01 U24872 (.o(n20871),
	.a(west_input_NIB_storage_data_f_0__43_),
	.b(FE_OFN25748_FE_OFN24796_n20854));
   oa12f01 U24873 (.o(n8333),
	.a(n20871),
	.b(FE_OFN25748_FE_OFN24796_n20854),
	.c(n21129));
   in01s01 U24874 (.o(n21105),
	.a(dataIn_W_42_));
   na02f01 U24875 (.o(n20872),
	.a(west_input_NIB_storage_data_f_0__42_),
	.b(FE_OFN25747_FE_OFN24796_n20854));
   oa12f01 U24876 (.o(n8338),
	.a(n20872),
	.b(FE_OFN25747_FE_OFN24796_n20854),
	.c(n21105));
   in01s01 U24877 (.o(n21107),
	.a(dataIn_W_41_));
   na02f01 U24878 (.o(n20873),
	.a(west_input_NIB_storage_data_f_0__41_),
	.b(FE_OFN25748_FE_OFN24796_n20854));
   oa12f01 U24879 (.o(n8343),
	.a(n20873),
	.b(FE_OFN25748_FE_OFN24796_n20854),
	.c(n21107));
   in01s01 U24880 (.o(n21109),
	.a(dataIn_W_40_));
   na02f01 U24881 (.o(n20874),
	.a(west_input_NIB_storage_data_f_0__40_),
	.b(FE_OFN25747_FE_OFN24796_n20854));
   oa12f01 U24882 (.o(n8348),
	.a(n20874),
	.b(FE_OFN25747_FE_OFN24796_n20854),
	.c(n21109));
   in01s01 U24883 (.o(n21111),
	.a(dataIn_W_39_));
   na02s01 U24884 (.o(n20875),
	.a(west_input_NIB_storage_data_f_0__39_),
	.b(FE_OFN25751_FE_OFN24796_n20854));
   oa12f01 U24885 (.o(n8353),
	.a(n20875),
	.b(FE_OFN25751_FE_OFN24796_n20854),
	.c(n21111));
   in01s01 U24886 (.o(n21113),
	.a(dataIn_W_38_));
   na02s01 U24887 (.o(n20876),
	.a(west_input_NIB_storage_data_f_0__38_),
	.b(FE_OFN25753_FE_OFN24796_n20854));
   oa12f01 U24888 (.o(n8358),
	.a(n20876),
	.b(FE_OFN25753_FE_OFN24796_n20854),
	.c(n21113));
   in01s01 U24889 (.o(n21115),
	.a(dataIn_W_37_));
   na02f01 U24890 (.o(n20877),
	.a(west_input_NIB_storage_data_f_0__37_),
	.b(FE_OFN25747_FE_OFN24796_n20854));
   oa12f01 U24891 (.o(n8363),
	.a(n20877),
	.b(FE_OFN25747_FE_OFN24796_n20854),
	.c(n21115));
   in01s01 U24892 (.o(n21117),
	.a(dataIn_W_36_));
   na02s01 U24893 (.o(n20878),
	.a(west_input_NIB_storage_data_f_0__36_),
	.b(FE_OFN25751_FE_OFN24796_n20854));
   in01s01 U24894 (.o(n21119),
	.a(dataIn_W_35_));
   na02f01 U24895 (.o(n20879),
	.a(west_input_NIB_storage_data_f_0__35_),
	.b(FE_OFN25748_FE_OFN24796_n20854));
   oa12f01 U24896 (.o(n8373),
	.a(n20879),
	.b(FE_OFN25748_FE_OFN24796_n20854),
	.c(n21119));
   in01s01 U24897 (.o(n21121),
	.a(dataIn_W_34_));
   na02s01 U24898 (.o(n20880),
	.a(west_input_NIB_storage_data_f_0__34_),
	.b(FE_OFN25753_FE_OFN24796_n20854));
   oa12s01 U24899 (.o(n8378),
	.a(n20880),
	.b(FE_OFN25753_FE_OFN24796_n20854),
	.c(n21121));
   in01s01 U24900 (.o(n22749),
	.a(dataIn_W_32_));
   na02f01 U24901 (.o(n20881),
	.a(west_input_NIB_storage_data_f_0__32_),
	.b(FE_OFN25748_FE_OFN24796_n20854));
   oa12f01 U24902 (.o(n8388),
	.a(n20881),
	.b(FE_OFN25748_FE_OFN24796_n20854),
	.c(n22749));
   in01f01 U24903 (.o(n22714),
	.a(dataIn_W_31_));
   na02f01 U24904 (.o(n20882),
	.a(west_input_NIB_storage_data_f_0__31_),
	.b(FE_OFN25747_FE_OFN24796_n20854));
   oa12f01 U24905 (.o(n8393),
	.a(n20882),
	.b(FE_OFN25747_FE_OFN24796_n20854),
	.c(n22714));
   in01s01 U24906 (.o(n22739),
	.a(dataIn_W_29_));
   na02s01 U24907 (.o(n20883),
	.a(west_input_NIB_storage_data_f_0__29_),
	.b(FE_OFN25749_FE_OFN24796_n20854));
   oa12s01 U24908 (.o(n8403),
	.a(n20883),
	.b(FE_OFN25749_FE_OFN24796_n20854),
	.c(n22739));
   na02s01 U24909 (.o(n20884),
	.a(west_input_NIB_storage_data_f_1__63_),
	.b(FE_OFN382_n17772));
   oa12s01 U24910 (.o(n8553),
	.a(n20884),
	.b(FE_OFN382_n17772),
	.c(n21072));
   na02s01 U24911 (.o(n20885),
	.a(west_input_NIB_storage_data_f_1__62_),
	.b(FE_OFN382_n17772));
   oa12s01 U24912 (.o(n8558),
	.a(n20885),
	.b(FE_OFN382_n17772),
	.c(n21093));
   na02f01 U24913 (.o(n20886),
	.a(west_input_NIB_storage_data_f_1__61_),
	.b(FE_OFN381_n17772));
   oa12f01 U24914 (.o(n8563),
	.a(n20886),
	.b(FE_OFN381_n17772),
	.c(n21095));
   na02s01 U24915 (.o(n20887),
	.a(west_input_NIB_storage_data_f_1__60_),
	.b(FE_OFN382_n17772));
   oa12s01 U24916 (.o(n8568),
	.a(n20887),
	.b(FE_OFN382_n17772),
	.c(n21097));
   in01s01 U24917 (.o(n21127),
	.a(dataIn_W_56_));
   na02s01 U24918 (.o(n20888),
	.a(west_input_NIB_storage_data_f_1__56_),
	.b(FE_OFN382_n17772));
   oa12s01 U24919 (.o(n8588),
	.a(n20888),
	.b(FE_OFN382_n17772),
	.c(n21127));
   in01s01 U24920 (.o(n22557),
	.a(dataIn_W_54_));
   na02f01 U24921 (.o(n20889),
	.a(west_input_NIB_storage_data_f_1__54_),
	.b(FE_OFN381_n17772));
   oa12f01 U24922 (.o(n8598),
	.a(n20889),
	.b(FE_OFN381_n17772),
	.c(n22557));
   na02s01 U24923 (.o(n20890),
	.a(west_input_NIB_storage_data_f_0__62_),
	.b(FE_OFN25750_FE_OFN24796_n20854));
   oa12s01 U24924 (.o(n8238),
	.a(n20890),
	.b(FE_OFN25750_FE_OFN24796_n20854),
	.c(n21093));
   na02s01 U24925 (.o(n20891),
	.a(west_input_NIB_storage_data_f_1__51_),
	.b(FE_OFN382_n17772));
   oa12s01 U24926 (.o(n8613),
	.a(n20891),
	.b(FE_OFN382_n17772),
	.c(n21084));
   na02f01 U24927 (.o(n20892),
	.a(west_input_NIB_storage_data_f_1__49_),
	.b(FE_OFN381_n17772));
   oa12f01 U24928 (.o(n8623),
	.a(n20892),
	.b(FE_OFN381_n17772),
	.c(n21091));
   na02f01 U24929 (.o(n20893),
	.a(west_input_NIB_storage_data_f_1__48_),
	.b(FE_OFN381_n17772));
   oa12f01 U24930 (.o(n8628),
	.a(n20893),
	.b(FE_OFN381_n17772),
	.c(n21099));
   na02s01 U24931 (.o(n20894),
	.a(west_input_NIB_storage_data_f_1__47_),
	.b(FE_OFN381_n17772));
   oa12f01 U24932 (.o(n8633),
	.a(n20894),
	.b(FE_OFN381_n17772),
	.c(n21125));
   na02s01 U24933 (.o(n20895),
	.a(west_input_NIB_storage_data_f_1__39_),
	.b(FE_OFN381_n17772));
   oa12s01 U24934 (.o(n8673),
	.a(n20895),
	.b(FE_OFN381_n17772),
	.c(n21111));
   na02s01 U24935 (.o(n20896),
	.a(west_input_NIB_storage_data_f_1__52_),
	.b(FE_OFN382_n17772));
   oa12s01 U24936 (.o(n8608),
	.a(n20896),
	.b(FE_OFN382_n17772),
	.c(n22717));
   na02f01 U24937 (.o(n20897),
	.a(west_input_NIB_storage_data_f_1__31_),
	.b(FE_OFN381_n17772));
   oa12f01 U24938 (.o(n8713),
	.a(n20897),
	.b(FE_OFN381_n17772),
	.c(n22714));
   in01s01 U24939 (.o(n22726),
	.a(dataIn_W_25_));
   na02s01 U24940 (.o(n20898),
	.a(west_input_NIB_storage_data_f_1__25_),
	.b(FE_OFN381_n17772));
   na02f01 U24941 (.o(n20899),
	.a(west_input_NIB_storage_data_f_1__45_),
	.b(FE_OFN381_n17772));
   oa12f01 U24942 (.o(n8643),
	.a(n20899),
	.b(FE_OFN381_n17772),
	.c(n21101));
   na02s01 U24943 (.o(n20900),
	.a(west_input_NIB_storage_data_f_1__38_),
	.b(FE_OFN381_n17772));
   oa12s01 U24944 (.o(n8678),
	.a(n20900),
	.b(FE_OFN381_n17772),
	.c(n21113));
   na02s01 U24945 (.o(n20901),
	.a(west_input_NIB_storage_data_f_1__37_),
	.b(FE_OFN381_n17772));
   oa12f01 U24946 (.o(n8683),
	.a(n20901),
	.b(FE_OFN381_n17772),
	.c(n21115));
   na02s01 U24947 (.o(n20902),
	.a(west_input_NIB_storage_data_f_1__36_),
	.b(FE_OFN381_n17772));
   oa12s01 U24948 (.o(n8688),
	.a(n20902),
	.b(FE_OFN381_n17772),
	.c(n21117));
   na02s01 U24949 (.o(n20903),
	.a(west_input_NIB_storage_data_f_1__41_),
	.b(FE_OFN381_n17772));
   oa12f01 U24950 (.o(n8663),
	.a(n20903),
	.b(FE_OFN381_n17772),
	.c(n21107));
   na02f01 U24951 (.o(n20904),
	.a(west_input_NIB_storage_data_f_1__35_),
	.b(FE_OFN381_n17772));
   oa12f01 U24952 (.o(n8693),
	.a(n20904),
	.b(FE_OFN381_n17772),
	.c(n21119));
   na02s01 U24953 (.o(n20905),
	.a(west_input_NIB_storage_data_f_1__34_),
	.b(FE_OFN381_n17772));
   oa12s01 U24954 (.o(n8698),
	.a(n20905),
	.b(FE_OFN381_n17772),
	.c(n21121));
   na02f01 U24955 (.o(n20906),
	.a(west_input_NIB_storage_data_f_1__40_),
	.b(FE_OFN381_n17772));
   na02f01 U24956 (.o(n20907),
	.a(west_input_NIB_storage_data_f_1__44_),
	.b(FE_OFN381_n17772));
   oa12f01 U24957 (.o(n8648),
	.a(n20907),
	.b(FE_OFN381_n17772),
	.c(n22486));
   na02f01 U24958 (.o(n20908),
	.a(west_input_NIB_storage_data_f_1__42_),
	.b(FE_OFN381_n17772));
   oa12f01 U24959 (.o(n8658),
	.a(n20908),
	.b(FE_OFN381_n17772),
	.c(n21105));
   na02s01 U24960 (.o(n20909),
	.a(west_input_NIB_storage_data_f_0__56_),
	.b(FE_OFN25750_FE_OFN24796_n20854));
   oa12s01 U24961 (.o(n8268),
	.a(n20909),
	.b(FE_OFN25750_FE_OFN24796_n20854),
	.c(n21127));
   na02f01 U24962 (.o(n20910),
	.a(west_input_NIB_storage_data_f_1__43_),
	.b(FE_OFN381_n17772));
   oa12f01 U24963 (.o(n8653),
	.a(n20910),
	.b(FE_OFN381_n17772),
	.c(n21129));
   no02f02 U24964 (.o(n20918),
	.a(n20917),
	.b(n20916));
   no02f01 U24965 (.o(n20922),
	.a(n20921),
	.b(n20920));
   no02f02 U24966 (.o(n20925),
	.a(n20924),
	.b(n20923));
   no02f02 U24968 (.o(n20931),
	.a(n20930),
	.b(n20929));
   in01s01 U24969 (.o(n20932),
	.a(north_input_NIB_tail_ptr_f_1_));
   na02s01 U24970 (.o(n20935),
	.a(north_input_NIB_storage_data_f_0__40_),
	.b(n20934));
   oa12s01 U24971 (.o(n12218),
	.a(n20935),
	.b(n20934),
	.c(n21262));
   na02s01 U24972 (.o(n20936),
	.a(north_input_NIB_storage_data_f_0__29_),
	.b(n20934));
   oa12s01 U24973 (.o(n12273),
	.a(n20936),
	.b(n20934),
	.c(n21248));
   na02s01 U24974 (.o(n20937),
	.a(north_input_NIB_storage_data_f_0__56_),
	.b(n17771));
   oa12s01 U24975 (.o(n12138),
	.a(n20937),
	.b(n17771),
	.c(n21277));
   na02s01 U24976 (.o(n20938),
	.a(north_input_NIB_storage_data_f_0__44_),
	.b(n20934));
   oa12s01 U24977 (.o(n12198),
	.a(n20938),
	.b(n20934),
	.c(n21272));
   na02s01 U24978 (.o(n20939),
	.a(north_input_NIB_storage_data_f_0__31_),
	.b(n20934));
   oa12s01 U24979 (.o(n12263),
	.a(n20939),
	.b(n20934),
	.c(n21237));
   na02s01 U24980 (.o(n20940),
	.a(north_input_NIB_storage_data_f_0__53_),
	.b(n20934));
   oa12s01 U24981 (.o(n12153),
	.a(n20940),
	.b(n20934),
	.c(n21285));
   na02s01 U24982 (.o(n20941),
	.a(north_input_NIB_storage_data_f_0__30_),
	.b(n20934));
   na02s01 U24983 (.o(n20942),
	.a(north_input_NIB_storage_data_f_0__25_),
	.b(n20934));
   oa12s01 U24984 (.o(n12293),
	.a(n20942),
	.b(n20934),
	.c(n21232));
   oa12s01 U24985 (.o(n12183),
	.a(n20943),
	.b(n20934),
	.c(n21234));
   na02s01 U24986 (.o(n20944),
	.a(north_input_NIB_storage_data_f_0__28_),
	.b(n20934));
   oa12s01 U24987 (.o(n12278),
	.a(n20944),
	.b(n20934),
	.c(n21243));
   na02s01 U24988 (.o(n20945),
	.a(north_input_NIB_storage_data_f_0__52_),
	.b(n17771));
   oa12s01 U24989 (.o(n12158),
	.a(n20945),
	.b(n17771),
	.c(n21280));
   na02s01 U24990 (.o(n20946),
	.a(north_input_NIB_storage_data_f_0__51_),
	.b(n17771));
   oa12s01 U24991 (.o(n12163),
	.a(n20946),
	.b(n17771),
	.c(n21239));
   na02s01 U24992 (.o(n20947),
	.a(north_input_NIB_storage_data_f_0__22_),
	.b(n20934));
   oa12s01 U24993 (.o(n12308),
	.a(n20947),
	.b(n20934),
	.c(n21226));
   na02s01 U24994 (.o(n20948),
	.a(north_input_NIB_storage_data_f_0__55_),
	.b(n17771));
   oa12s01 U24995 (.o(n12143),
	.a(n20948),
	.b(n17771),
	.c(n21254));
   na02s01 U24996 (.o(n20949),
	.a(north_input_NIB_storage_data_f_0__27_),
	.b(n20934));
   oa12s01 U24997 (.o(n12283),
	.a(n20949),
	.b(n20934),
	.c(n21250));
   na02s01 U24998 (.o(n20950),
	.a(north_input_NIB_storage_data_f_0__57_),
	.b(n17771));
   oa12s01 U24999 (.o(n12133),
	.a(n20950),
	.b(n17771),
	.c(n21274));
   na02s01 U25000 (.o(n20951),
	.a(north_input_NIB_storage_data_f_0__58_),
	.b(n17771));
   oa12s01 U25001 (.o(n12128),
	.a(n20951),
	.b(n17771),
	.c(n21256));
   na02s01 U25002 (.o(n20952),
	.a(north_input_NIB_storage_data_f_0__60_),
	.b(n17771));
   oa12s01 U25003 (.o(n12108),
	.a(n20953),
	.b(n17771),
	.c(n21246));
   na02s01 U25004 (.o(n20954),
	.a(north_input_NIB_storage_data_f_0__63_),
	.b(n17771));
   oa12s01 U25005 (.o(n12103),
	.a(n20954),
	.b(n17771),
	.c(n21241));
   na02s01 U25006 (.o(n20955),
	.a(north_input_NIB_storage_data_f_0__26_),
	.b(n20934));
   oa12s01 U25007 (.o(n12288),
	.a(n20955),
	.b(n20934),
	.c(n21266));
   na02s01 U25008 (.o(n20956),
	.a(north_input_NIB_storage_data_f_0__23_),
	.b(n20934));
   oa12s01 U25009 (.o(n12303),
	.a(n20956),
	.b(n20934),
	.c(n21222));
   na02s01 U25010 (.o(n20957),
	.a(north_input_NIB_storage_data_f_0__54_),
	.b(n17771));
   oa12s01 U25011 (.o(n12148),
	.a(n20957),
	.b(n17771),
	.c(n21270));
   na02s01 U25012 (.o(n20958),
	.a(north_input_NIB_storage_data_f_0__41_),
	.b(n20934));
   oa12s01 U25013 (.o(n12213),
	.a(n20958),
	.b(n20934),
	.c(n21264));
   na02s01 U25014 (.o(n20959),
	.a(north_input_NIB_storage_data_f_0__24_),
	.b(n20934));
   oa12s01 U25015 (.o(n12298),
	.a(n20959),
	.b(n20934),
	.c(n21224));
   na02s01 U25016 (.o(n20960),
	.a(north_input_NIB_storage_data_f_0__50_),
	.b(n20934));
   oa12s01 U25017 (.o(n12168),
	.a(n20960),
	.b(n20934),
	.c(n21282));
   in01s01 U25020 (.o(n20969),
	.a(south_input_NIB_tail_ptr_f_1_));
   no02f02 U25021 (.o(n20994),
	.a(n20970),
	.b(n20969));
   in01s01 U25022 (.o(n22686),
	.a(dataIn_S_63_));
   na02f01 U25023 (.o(n20973),
	.a(south_input_NIB_storage_data_f_2__63_),
	.b(n25905));
   na02f01 U25024 (.o(n20974),
	.a(south_input_NIB_storage_data_f_2__28_),
	.b(FE_OFN84_n20972));
   oa12f01 U25025 (.o(n10338),
	.a(n20974),
	.b(n21030),
	.c(FE_OFN84_n20972));
   na02f02 U25026 (.o(n20975),
	.a(south_input_NIB_storage_data_f_2__60_),
	.b(n25905));
   oa12f01 U25027 (.o(n10178),
	.a(n20975),
	.b(n25905),
	.c(n21016));
   na02f01 U25028 (.o(n20976),
	.a(south_input_NIB_storage_data_f_2__61_),
	.b(n25905));
   oa12f01 U25029 (.o(n10173),
	.a(n20976),
	.b(n25905),
	.c(n21012));
   na02f01 U25030 (.o(n20977),
	.a(south_input_NIB_storage_data_f_2__58_),
	.b(n25905));
   oa12f01 U25031 (.o(n10188),
	.a(n20977),
	.b(n25905),
	.c(n21022));
   na02f01 U25032 (.o(n20978),
	.a(south_input_NIB_storage_data_f_2__59_),
	.b(n25905));
   oa12f01 U25033 (.o(n10183),
	.a(n20978),
	.b(n25905),
	.c(n21018));
   na02f01 U25034 (.o(n20979),
	.a(south_input_NIB_storage_data_f_2__56_),
	.b(n25905));
   oa12f01 U25035 (.o(n10198),
	.a(n20979),
	.b(n25905),
	.c(n21037));
   na02f01 U25036 (.o(n20980),
	.a(south_input_NIB_storage_data_f_2__55_),
	.b(n25905));
   oa12f01 U25037 (.o(n10203),
	.a(n20980),
	.b(n25905),
	.c(n21014));
   na02f01 U25038 (.o(n20981),
	.a(south_input_NIB_storage_data_f_2__54_),
	.b(n25905));
   oa12f01 U25039 (.o(n10208),
	.a(n20981),
	.b(n25905),
	.c(n21040));
   na02f01 U25040 (.o(n20982),
	.a(south_input_NIB_storage_data_f_2__53_),
	.b(n25905));
   oa12f01 U25041 (.o(n10213),
	.a(n20982),
	.b(n25905),
	.c(n21042));
   in01s01 U25042 (.o(n22484),
	.a(dataIn_S_51_));
   na02f01 U25043 (.o(n20983),
	.a(south_input_NIB_storage_data_f_2__51_),
	.b(n25905));
   oa12f01 U25044 (.o(n10223),
	.a(n20983),
	.b(n25905),
	.c(n22484));
   na02f01 U25045 (.o(n20984),
	.a(south_input_NIB_storage_data_f_2__62_),
	.b(n25905));
   na02f01 U25046 (.o(n20985),
	.a(south_input_NIB_storage_data_f_2__50_),
	.b(n25905));
   oa12f01 U25047 (.o(n10228),
	.a(n20985),
	.b(n25905),
	.c(n21035));
   na02f01 U25048 (.o(n20986),
	.a(south_input_NIB_storage_data_f_2__49_),
	.b(FE_OFN84_n20972));
   oa12f01 U25049 (.o(n10233),
	.a(n20986),
	.b(FE_OFN84_n20972),
	.c(n20998));
   na02f01 U25050 (.o(n20987),
	.a(south_input_NIB_storage_data_f_2__40_),
	.b(n25905));
   oa12f01 U25051 (.o(n10278),
	.a(n20987),
	.b(n25905),
	.c(n21020));
   in01s01 U25052 (.o(n22582),
	.a(dataIn_S_39_));
   na02f01 U25053 (.o(n20988),
	.a(south_input_NIB_storage_data_f_2__39_),
	.b(FE_OFN84_n20972));
   oa12f01 U25054 (.o(n10283),
	.a(n20988),
	.b(FE_OFN84_n20972),
	.c(n22582));
   na02f01 U25055 (.o(n20989),
	.a(south_input_NIB_storage_data_f_2__34_),
	.b(FE_OFN84_n20972));
   na02f01 U25056 (.o(n20990),
	.a(south_input_NIB_storage_data_f_2__30_),
	.b(FE_OFN84_n20972));
   oa12f01 U25057 (.o(n10328),
	.a(n20990),
	.b(FE_OFN84_n20972),
	.c(n21024));
   na02f01 U25058 (.o(n20991),
	.a(south_input_NIB_storage_data_f_2__29_),
	.b(FE_OFN84_n20972));
   oa12f01 U25059 (.o(n10333),
	.a(n20991),
	.b(FE_OFN84_n20972),
	.c(n21049));
   na02f01 U25060 (.o(n20992),
	.a(south_input_NIB_storage_data_f_2__57_),
	.b(n25905));
   oa12f01 U25061 (.o(n10193),
	.a(n20992),
	.b(n25905),
	.c(n21026));
   oa12f01 U25062 (.o(n10343),
	.a(n20993),
	.b(FE_OFN84_n20972),
	.c(n21005));
   na02f02 U25063 (.o(n20995),
	.a(n20994),
	.b(south_input_NIB_tail_ptr_f_0_));
   na02s01 U25064 (.o(n20997),
	.a(south_input_NIB_storage_data_f_3__49_),
	.b(n17769));
   oa12s01 U25065 (.o(n10553),
	.a(n20997),
	.b(n20998),
	.c(n17769));
   na02f01 U25066 (.o(n20999),
	.a(south_input_NIB_storage_data_f_2__26_),
	.b(FE_OFN84_n20972));
   oa12f01 U25067 (.o(n10348),
	.a(n20999),
	.b(FE_OFN84_n20972),
	.c(n21032));
   na02f01 U25068 (.o(n21000),
	.a(south_input_NIB_storage_data_f_2__25_),
	.b(FE_OFN84_n20972));
   na02f01 U25069 (.o(n21001),
	.a(south_input_NIB_storage_data_f_2__24_),
	.b(FE_OFN84_n20972));
   na02f01 U25070 (.o(n21002),
	.a(south_input_NIB_storage_data_f_2__23_),
	.b(FE_OFN84_n20972));
   na02f01 U25071 (.o(n21003),
	.a(south_input_NIB_storage_data_f_2__22_),
	.b(FE_OFN84_n20972));
   na02s01 U25072 (.o(n21004),
	.a(south_input_NIB_storage_data_f_3__27_),
	.b(n17769));
   oa12s01 U25073 (.o(n10663),
	.a(n21004),
	.b(n21005),
	.c(n17769));
   na02s01 U25074 (.o(n21006),
	.a(south_input_NIB_storage_data_f_3__62_),
	.b(FE_OFN896_n17769));
   oa12s01 U25075 (.o(n10488),
	.a(n21006),
	.b(n21007),
	.c(FE_OFN896_n17769));
   na02s01 U25076 (.o(n21008),
	.a(south_input_NIB_storage_data_f_3__25_),
	.b(n17769));
   oa12s01 U25077 (.o(n10673),
	.a(n21008),
	.b(n21009),
	.c(n17769));
   na02s01 U25078 (.o(n21010),
	.a(south_input_NIB_storage_data_f_3__41_),
	.b(n17769));
   oa12s01 U25079 (.o(n10593),
	.a(n21010),
	.b(n17769),
	.c(n22688));
   na02s01 U25080 (.o(n21011),
	.a(south_input_NIB_storage_data_f_3__61_),
	.b(FE_OFN896_n17769));
   oa12s01 U25081 (.o(n10493),
	.a(n21011),
	.b(n21012),
	.c(FE_OFN896_n17769));
   na02s01 U25082 (.o(n21013),
	.a(south_input_NIB_storage_data_f_3__55_),
	.b(FE_OFN896_n17769));
   oa12s01 U25083 (.o(n10523),
	.a(n21013),
	.b(n21014),
	.c(FE_OFN896_n17769));
   na02s01 U25084 (.o(n21015),
	.a(south_input_NIB_storage_data_f_3__60_),
	.b(FE_OFN896_n17769));
   oa12s01 U25085 (.o(n10498),
	.a(n21015),
	.b(n21016),
	.c(FE_OFN896_n17769));
   na02s01 U25086 (.o(n21017),
	.a(south_input_NIB_storage_data_f_3__59_),
	.b(FE_OFN896_n17769));
   oa12s01 U25087 (.o(n10503),
	.a(n21017),
	.b(n21018),
	.c(FE_OFN896_n17769));
   na02s01 U25088 (.o(n21019),
	.a(south_input_NIB_storage_data_f_3__40_),
	.b(FE_OFN896_n17769));
   oa12s01 U25089 (.o(n10598),
	.a(n21019),
	.b(n21020),
	.c(FE_OFN896_n17769));
   na02s01 U25090 (.o(n21021),
	.a(south_input_NIB_storage_data_f_3__58_),
	.b(FE_OFN896_n17769));
   oa12s01 U25091 (.o(n10508),
	.a(n21021),
	.b(n21022),
	.c(FE_OFN896_n17769));
   na02s01 U25092 (.o(n21023),
	.a(south_input_NIB_storage_data_f_3__30_),
	.b(n17769));
   oa12s01 U25093 (.o(n10648),
	.a(n21023),
	.b(n21024),
	.c(n17769));
   na02s01 U25094 (.o(n21025),
	.a(south_input_NIB_storage_data_f_3__57_),
	.b(FE_OFN896_n17769));
   oa12s01 U25095 (.o(n10513),
	.a(n21025),
	.b(n21026),
	.c(FE_OFN896_n17769));
   na02s01 U25096 (.o(n21027),
	.a(south_input_NIB_storage_data_f_3__22_),
	.b(n17769));
   oa12s01 U25097 (.o(n10688),
	.a(n21027),
	.b(n21028),
	.c(n17769));
   na02s01 U25098 (.o(n21029),
	.a(south_input_NIB_storage_data_f_3__28_),
	.b(n17769));
   oa12s01 U25099 (.o(n10658),
	.a(n21029),
	.b(n17769),
	.c(n21030));
   oa12s01 U25100 (.o(n10668),
	.a(n21031),
	.b(n21032),
	.c(n17769));
   na02s01 U25101 (.o(n21033),
	.a(south_input_NIB_storage_data_f_3__52_),
	.b(FE_OFN896_n17769));
   oa12s01 U25102 (.o(n10538),
	.a(n21033),
	.b(n22482),
	.c(FE_OFN896_n17769));
   na02s01 U25103 (.o(n21034),
	.a(south_input_NIB_storage_data_f_3__50_),
	.b(FE_OFN896_n17769));
   oa12s01 U25104 (.o(n10548),
	.a(n21034),
	.b(n21035),
	.c(FE_OFN896_n17769));
   na02s01 U25105 (.o(n21036),
	.a(south_input_NIB_storage_data_f_3__56_),
	.b(FE_OFN896_n17769));
   oa12s01 U25106 (.o(n10518),
	.a(n21036),
	.b(n21037),
	.c(FE_OFN896_n17769));
   na02s01 U25107 (.o(n21038),
	.a(south_input_NIB_storage_data_f_3__48_),
	.b(n17769));
   oa12s01 U25108 (.o(n10558),
	.a(n21038),
	.b(n22679),
	.c(n17769));
   na02s01 U25109 (.o(n21039),
	.a(south_input_NIB_storage_data_f_3__54_),
	.b(FE_OFN896_n17769));
   oa12s01 U25110 (.o(n10528),
	.a(n21039),
	.b(n21040),
	.c(FE_OFN896_n17769));
   na02s01 U25111 (.o(n21041),
	.a(south_input_NIB_storage_data_f_3__53_),
	.b(FE_OFN896_n17769));
   oa12s01 U25112 (.o(n10533),
	.a(n21041),
	.b(n21042),
	.c(FE_OFN896_n17769));
   na02s01 U25113 (.o(n21043),
	.a(south_input_NIB_storage_data_f_3__24_),
	.b(n17769));
   oa12s01 U25114 (.o(n10678),
	.a(n21043),
	.b(n21044),
	.c(n17769));
   na02s01 U25115 (.o(n21045),
	.a(south_input_NIB_storage_data_f_3__23_),
	.b(n17769));
   oa12s01 U25116 (.o(n10683),
	.a(n21045),
	.b(n21046),
	.c(n17769));
   na02s01 U25117 (.o(n21047),
	.a(south_input_NIB_storage_data_f_3__39_),
	.b(n17769));
   oa12s01 U25118 (.o(n10603),
	.a(n21047),
	.b(n22582),
	.c(n17769));
   na02s01 U25119 (.o(n21048),
	.a(south_input_NIB_storage_data_f_3__29_),
	.b(n17769));
   oa12s01 U25120 (.o(n10653),
	.a(n21048),
	.b(n21049),
	.c(n17769));
   in01s01 U25121 (.o(n21050),
	.a(west_input_NIB_tail_ptr_f_1_));
   no02f02 U25122 (.o(n21068),
	.a(n21051),
	.b(n21050));
   na02f01 U25123 (.o(n21054),
	.a(west_input_NIB_storage_data_f_2__60_),
	.b(FE_OFN25791_n21053));
   na02f01 U25124 (.o(n21055),
	.a(west_input_NIB_storage_data_f_2__50_),
	.b(FE_OFN25792_n21053));
   oa12f01 U25125 (.o(n8938),
	.a(n21055),
	.b(FE_OFN25792_n21053),
	.c(n21086));
   na02f01 U25126 (.o(n21056),
	.a(west_input_NIB_storage_data_f_2__39_),
	.b(n21053));
   oa12f01 U25127 (.o(n8993),
	.a(n21056),
	.b(n21053),
	.c(n21111));
   in01s01 U25128 (.o(n22488),
	.a(dataIn_W_53_));
   na02f01 U25129 (.o(n21057),
	.a(west_input_NIB_storage_data_f_2__53_),
	.b(FE_OFN25792_n21053));
   oa12f01 U25130 (.o(n8923),
	.a(n21057),
	.b(FE_OFN25792_n21053),
	.c(n22488));
   na02f01 U25131 (.o(n21058),
	.a(west_input_NIB_storage_data_f_2__61_),
	.b(FE_OFN25792_n21053));
   oa12f01 U25132 (.o(n8883),
	.a(n21058),
	.b(FE_OFN25792_n21053),
	.c(n21095));
   na02f01 U25133 (.o(n21059),
	.a(west_input_NIB_storage_data_f_2__36_),
	.b(n21053));
   na02f01 U25134 (.o(n21060),
	.a(west_input_NIB_storage_data_f_2__38_),
	.b(FE_OFN25794_n21053));
   na02f01 U25135 (.o(n21061),
	.a(west_input_NIB_storage_data_f_2__63_),
	.b(FE_OFN25791_n21053));
   na02f01 U25136 (.o(n21062),
	.a(west_input_NIB_storage_data_f_2__35_),
	.b(FE_OFN25792_n21053));
   na02f01 U25137 (.o(n21063),
	.a(west_input_NIB_storage_data_f_2__62_),
	.b(FE_OFN25791_n21053));
   oa12f01 U25138 (.o(n8878),
	.a(n21063),
	.b(FE_OFN25791_n21053),
	.c(n21093));
   na02f01 U25139 (.o(n21064),
	.a(west_input_NIB_storage_data_f_2__45_),
	.b(FE_OFN25792_n21053));
   na02f01 U25140 (.o(n21065),
	.a(west_input_NIB_storage_data_f_2__34_),
	.b(FE_OFN25794_n21053));
   na02f01 U25141 (.o(n21066),
	.a(west_input_NIB_storage_data_f_2__29_),
	.b(n21053));
   in01s01 U25142 (.o(n22751),
	.a(dataIn_W_26_));
   na02f01 U25143 (.o(n21067),
	.a(west_input_NIB_storage_data_f_2__26_),
	.b(n21053));
   na02f01 U25144 (.o(n21071),
	.a(west_input_NIB_storage_data_f_3__63_),
	.b(FE_OFN24767_n21069));
   na02f01 U25145 (.o(n21073),
	.a(west_input_NIB_storage_data_f_2__42_),
	.b(FE_OFN25792_n21053));
   oa12f01 U25146 (.o(n8978),
	.a(n21073),
	.b(n21105),
	.c(FE_OFN25792_n21053));
   na02f01 U25147 (.o(n21074),
	.a(west_input_NIB_storage_data_f_2__41_),
	.b(FE_OFN25792_n21053));
   oa12f01 U25148 (.o(n8983),
	.a(n21074),
	.b(FE_OFN25792_n21053),
	.c(n21107));
   na02f01 U25149 (.o(n21075),
	.a(west_input_NIB_storage_data_f_2__40_),
	.b(FE_OFN25792_n21053));
   oa12f01 U25150 (.o(n8988),
	.a(n21075),
	.b(FE_OFN25792_n21053),
	.c(n21109));
   na02f01 U25151 (.o(n21076),
	.a(west_input_NIB_storage_data_f_3__54_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25152 (.o(n9238),
	.a(n21076),
	.b(n22557),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U25153 (.o(n21077),
	.a(west_input_NIB_storage_data_f_2__56_),
	.b(FE_OFN25791_n21053));
   oa12f01 U25154 (.o(n8908),
	.a(n21077),
	.b(FE_OFN25791_n21053),
	.c(n21127));
   na02f01 U25155 (.o(n21078),
	.a(west_input_NIB_storage_data_f_2__37_),
	.b(FE_OFN25792_n21053));
   na02f01 U25156 (.o(n21079),
	.a(west_input_NIB_storage_data_f_2__54_),
	.b(FE_OFN25792_n21053));
   oa12f01 U25157 (.o(n8918),
	.a(n21079),
	.b(FE_OFN25792_n21053),
	.c(n22557));
   na02f01 U25158 (.o(n21080),
	.a(west_input_NIB_storage_data_f_2__49_),
	.b(FE_OFN25792_n21053));
   oa12f01 U25159 (.o(n8943),
	.a(n21080),
	.b(FE_OFN25792_n21053),
	.c(n21091));
   na02f01 U25160 (.o(n21081),
	.a(west_input_NIB_storage_data_f_3__52_),
	.b(FE_OFN24767_n21069));
   oa12f01 U25161 (.o(n9248),
	.a(n21081),
	.b(n22717),
	.c(FE_OFN24767_n21069));
   na02f01 U25162 (.o(n21082),
	.a(west_input_NIB_storage_data_f_2__51_),
	.b(FE_OFN25791_n21053));
   oa12f01 U25163 (.o(n8933),
	.a(n21082),
	.b(FE_OFN25791_n21053),
	.c(n21084));
   na02f01 U25164 (.o(n21083),
	.a(west_input_NIB_storage_data_f_3__51_),
	.b(FE_OFN24767_n21069));
   oa12f01 U25165 (.o(n9253),
	.a(n21083),
	.b(n21084),
	.c(FE_OFN24767_n21069));
   na02f01 U25166 (.o(n21085),
	.a(west_input_NIB_storage_data_f_3__50_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25167 (.o(n9258),
	.a(n21085),
	.b(n21086),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U25168 (.o(n21087),
	.a(west_input_NIB_storage_data_f_2__48_),
	.b(FE_OFN25792_n21053));
   oa12f01 U25169 (.o(n8948),
	.a(n21087),
	.b(FE_OFN25792_n21053),
	.c(n21099));
   na02f01 U25170 (.o(n21088),
	.a(west_input_NIB_storage_data_f_2__47_),
	.b(FE_OFN25792_n21053));
   oa12f01 U25171 (.o(n8953),
	.a(n21088),
	.b(FE_OFN25792_n21053),
	.c(n21125));
   in01s01 U25172 (.o(n22743),
	.a(dataIn_W_46_));
   na02f01 U25173 (.o(n21089),
	.a(west_input_NIB_storage_data_f_2__46_),
	.b(FE_OFN25792_n21053));
   oa12f01 U25174 (.o(n8958),
	.a(n21089),
	.b(FE_OFN25792_n21053),
	.c(n22743));
   na02f01 U25175 (.o(n21090),
	.a(west_input_NIB_storage_data_f_3__49_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U25176 (.o(n21092),
	.a(west_input_NIB_storage_data_f_3__62_),
	.b(FE_OFN24767_n21069));
   oa12f01 U25177 (.o(n9198),
	.a(n21092),
	.b(n21093),
	.c(FE_OFN24767_n21069));
   na02f01 U25178 (.o(n21094),
	.a(west_input_NIB_storage_data_f_3__61_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25179 (.o(n9203),
	.a(n21094),
	.b(n21095),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U25180 (.o(n21096),
	.a(west_input_NIB_storage_data_f_3__60_),
	.b(FE_OFN24767_n21069));
   oa12f01 U25181 (.o(n9208),
	.a(n21096),
	.b(n21097),
	.c(FE_OFN24767_n21069));
   na02f01 U25182 (.o(n21098),
	.a(west_input_NIB_storage_data_f_3__48_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U25183 (.o(n21100),
	.a(west_input_NIB_storage_data_f_3__45_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25184 (.o(n9283),
	.a(n21100),
	.b(FE_OFN25866_FE_OFN24766_n21069),
	.c(n21101));
   na02f01 U25185 (.o(n21102),
	.a(west_input_NIB_storage_data_f_3__44_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25186 (.o(n9288),
	.a(n21102),
	.b(n22486),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U25187 (.o(n21103),
	.a(west_input_NIB_storage_data_f_3__43_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25188 (.o(n9293),
	.a(n21103),
	.b(FE_OFN25866_FE_OFN24766_n21069),
	.c(n21129));
   na02f01 U25189 (.o(n21104),
	.a(west_input_NIB_storage_data_f_3__42_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25190 (.o(n9298),
	.a(n21104),
	.b(FE_OFN25866_FE_OFN24766_n21069),
	.c(n21105));
   na02f01 U25191 (.o(n21106),
	.a(west_input_NIB_storage_data_f_3__41_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25192 (.o(n9303),
	.a(n21106),
	.b(n21107),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U25193 (.o(n21108),
	.a(west_input_NIB_storage_data_f_3__40_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25194 (.o(n9308),
	.a(n21108),
	.b(n21109),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U25195 (.o(n21110),
	.a(west_input_NIB_storage_data_f_3__39_),
	.b(FE_OFN24766_n21069));
   oa12f01 U25196 (.o(n9313),
	.a(n21110),
	.b(n21111),
	.c(FE_OFN24766_n21069));
   na02f01 U25197 (.o(n21112),
	.a(west_input_NIB_storage_data_f_3__38_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25198 (.o(n9318),
	.a(n21112),
	.b(n21113),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U25199 (.o(n21114),
	.a(west_input_NIB_storage_data_f_3__37_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25200 (.o(n9323),
	.a(n21114),
	.b(n21115),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U25201 (.o(n21116),
	.a(west_input_NIB_storage_data_f_3__36_),
	.b(FE_OFN25862_FE_OFN24766_n21069));
   oa12f01 U25202 (.o(n9328),
	.a(n21116),
	.b(n21117),
	.c(FE_OFN25862_FE_OFN24766_n21069));
   na02f01 U25203 (.o(n21118),
	.a(west_input_NIB_storage_data_f_3__35_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25204 (.o(n9333),
	.a(n21118),
	.b(n21119),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U25205 (.o(n21120),
	.a(west_input_NIB_storage_data_f_3__34_),
	.b(FE_OFN24766_n21069));
   oa12f01 U25206 (.o(n9338),
	.a(n21120),
	.b(FE_OFN24766_n21069),
	.c(n21121));
   na02f01 U25207 (.o(n21123),
	.a(west_input_NIB_storage_data_f_3__25_),
	.b(FE_OFN24766_n21069));
   na02f01 U25208 (.o(n21124),
	.a(west_input_NIB_storage_data_f_3__47_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U25209 (.o(n9273),
	.a(n21124),
	.b(n21125),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U25210 (.o(n21126),
	.a(west_input_NIB_storage_data_f_3__56_),
	.b(FE_OFN24767_n21069));
   oa12f01 U25211 (.o(n9228),
	.a(n21126),
	.b(n21127),
	.c(FE_OFN24767_n21069));
   na02f01 U25212 (.o(n21128),
	.a(west_input_NIB_storage_data_f_2__43_),
	.b(FE_OFN25792_n21053));
   oa12f01 U25213 (.o(n8973),
	.a(n21128),
	.b(n21129),
	.c(FE_OFN25792_n21053));
   na02f02 U25215 (.o(n21136),
	.a(n21135),
	.b(n21134));
   no02f02 U25217 (.o(n21140),
	.a(n21139),
	.b(n21138));
   no02f01 U25218 (.o(n21147),
	.a(n21146),
	.b(n21145));
   na03f03 U25219 (.o(dataOut_E_46_),
	.a(n21150),
	.b(n21149),
	.c(n21148));
   in01s01 U25220 (.o(n21570),
	.a(east_input_control_count_f_6_));
   na02f01 U25221 (.o(n21899),
	.a(east_input_control_thanks_all_f),
	.b(FE_OFN100_n21907));
   na02s01 U25222 (.o(n21153),
	.a(n21902),
	.b(n21156));
   na02s01 U25223 (.o(n21152),
	.a(n21570),
	.b(n21153));
   in01s01 U25224 (.o(east_input_control_N47),
	.a(n21155));
   ao12s01 U25225 (.o(n21158),
	.a(n21156),
	.b(east_input_control_count_f_0_),
	.c(east_input_control_count_f_1_));
   in01s01 U25226 (.o(n21157),
	.a(east_input_control_count_f_1_));
   in01s01 U25227 (.o(east_input_control_N42),
	.a(n21159));
   in01f01 U25228 (.o(n23632),
	.a(n21161));
   na02f01 U25229 (.o(n21166),
	.a(n21165),
	.b(n21164));
   ao22f01 U25231 (.o(n21169),
	.a(FE_OFN42_n19022),
	.b(n23632),
	.c(n19019),
	.d(n23630));
   ao22f01 U25232 (.o(n21168),
	.a(FE_OFN35_n19017),
	.b(n23629),
	.c(n19020),
	.d(FE_OFN479_n23631));
   na02f02 U25233 (.o(n21170),
	.a(n21169),
	.b(n21168));
   in01s01 U25234 (.o(n21171),
	.a(n21170));
   na02s01 U25235 (.o(n21172),
	.a(north_input_NIB_tail_ptr_f_1_),
	.b(north_input_NIB_tail_ptr_f_0_));
   na02f01 U25236 (.o(n21176),
	.a(north_input_NIB_storage_data_f_3__57_),
	.b(FE_OFN86_n21175));
   oa12f01 U25237 (.o(n13098),
	.a(n21177),
	.b(FE_OFN86_n21175),
	.c(n21277));
   na02f01 U25238 (.o(n21178),
	.a(north_input_NIB_storage_data_f_3__55_),
	.b(FE_OFN86_n21175));
   oa12f01 U25239 (.o(n13103),
	.a(n21178),
	.b(FE_OFN86_n21175),
	.c(n21254));
   na02f01 U25240 (.o(n21179),
	.a(north_input_NIB_storage_data_f_3__22_),
	.b(n25836));
   na02f01 U25241 (.o(n21180),
	.a(north_input_NIB_storage_data_f_3__52_),
	.b(FE_OFN86_n21175));
   oa12f01 U25242 (.o(n13118),
	.a(n21180),
	.b(FE_OFN86_n21175),
	.c(n21280));
   na02f01 U25243 (.o(n21181),
	.a(north_input_NIB_storage_data_f_3__51_),
	.b(FE_OFN86_n21175));
   oa12f01 U25244 (.o(n13123),
	.a(n21181),
	.b(FE_OFN86_n21175),
	.c(n21239));
   na02f01 U25245 (.o(n21182),
	.a(north_input_NIB_storage_data_f_3__25_),
	.b(n25836));
   oa12f01 U25246 (.o(n13253),
	.a(n21182),
	.b(n25836),
	.c(n21232));
   na02f01 U25247 (.o(n21183),
	.a(north_input_NIB_storage_data_f_3__54_),
	.b(FE_OFN86_n21175));
   oa12f01 U25248 (.o(n13108),
	.a(n21183),
	.b(FE_OFN86_n21175),
	.c(n21270));
   na02f01 U25249 (.o(n21184),
	.a(north_input_NIB_storage_data_f_3__53_),
	.b(n25836));
   oa12f01 U25250 (.o(n13113),
	.a(n21184),
	.b(n25836),
	.c(n21285));
   na02f01 U25251 (.o(n21185),
	.a(north_input_NIB_storage_data_f_3__58_),
	.b(FE_OFN86_n21175));
   na02f01 U25252 (.o(n21186),
	.a(north_input_NIB_storage_data_f_3__59_),
	.b(FE_OFN86_n21175));
   oa12f01 U25253 (.o(n13083),
	.a(n21186),
	.b(FE_OFN86_n21175),
	.c(n22642));
   na02f01 U25254 (.o(n21187),
	.a(north_input_NIB_storage_data_f_3__39_),
	.b(n25836));
   oa12f01 U25255 (.o(n13183),
	.a(n21187),
	.b(n25836),
	.c(n22646));
   na02f01 U25256 (.o(n21188),
	.a(north_input_NIB_storage_data_f_3__60_),
	.b(FE_OFN86_n21175));
   oa12f01 U25257 (.o(n13078),
	.a(n21188),
	.b(FE_OFN86_n21175),
	.c(n21287));
   na02f01 U25258 (.o(n21189),
	.a(north_input_NIB_storage_data_f_3__61_),
	.b(FE_OFN86_n21175));
   oa12f01 U25259 (.o(n13073),
	.a(n21189),
	.b(FE_OFN86_n21175),
	.c(n22444));
   na02f01 U25260 (.o(n21190),
	.a(north_input_NIB_storage_data_f_3__62_),
	.b(FE_OFN86_n21175));
   oa12f01 U25261 (.o(n13068),
	.a(n21190),
	.b(FE_OFN86_n21175),
	.c(n21246));
   na02f01 U25262 (.o(n21191),
	.a(north_input_NIB_storage_data_f_3__63_),
	.b(FE_OFN86_n21175));
   oa12f01 U25263 (.o(n13063),
	.a(n21191),
	.b(FE_OFN86_n21175),
	.c(n21241));
   na02f01 U25264 (.o(n21192),
	.a(north_input_NIB_storage_data_f_3__48_),
	.b(n25836));
   oa12f01 U25265 (.o(n13138),
	.a(n21192),
	.b(n25836),
	.c(n22652));
   na02f01 U25266 (.o(n21193),
	.a(north_input_NIB_storage_data_f_3__49_),
	.b(n25836));
   oa12f01 U25267 (.o(n13133),
	.a(n21193),
	.b(n25836),
	.c(n22634));
   na02f01 U25268 (.o(n21194),
	.a(north_input_NIB_storage_data_f_3__47_),
	.b(n25836));
   oa12f01 U25269 (.o(n13143),
	.a(n21194),
	.b(n25836),
	.c(n21234));
   na02f01 U25270 (.o(n21195),
	.a(north_input_NIB_storage_data_f_3__46_),
	.b(n25836));
   oa12f01 U25271 (.o(n13148),
	.a(n21195),
	.b(n25836),
	.c(n22636));
   na02f01 U25272 (.o(n21196),
	.a(north_input_NIB_storage_data_f_3__45_),
	.b(n25836));
   oa12f01 U25273 (.o(n13153),
	.a(n21196),
	.b(n25836),
	.c(n22632));
   na02f01 U25274 (.o(n21197),
	.a(north_input_NIB_storage_data_f_3__44_),
	.b(n25836));
   oa12f01 U25275 (.o(n13158),
	.a(n21197),
	.b(n25836),
	.c(n21272));
   na02f01 U25276 (.o(n21198),
	.a(north_input_NIB_storage_data_f_3__43_),
	.b(n25836));
   na02f01 U25277 (.o(n21199),
	.a(north_input_NIB_storage_data_f_3__42_),
	.b(n25836));
   na02f01 U25278 (.o(n21200),
	.a(north_input_NIB_storage_data_f_3__41_),
	.b(n25836));
   oa12f01 U25279 (.o(n13173),
	.a(n21200),
	.b(n25836),
	.c(n21264));
   na02f01 U25280 (.o(n21201),
	.a(north_input_NIB_storage_data_f_3__40_),
	.b(n25836));
   oa12f01 U25281 (.o(n13178),
	.a(n21201),
	.b(n25836),
	.c(n21262));
   na02f01 U25282 (.o(n21202),
	.a(north_input_NIB_storage_data_f_3__38_),
	.b(n25836));
   oa12f01 U25283 (.o(n13188),
	.a(n21202),
	.b(n25836),
	.c(n22638));
   na02f01 U25284 (.o(n21203),
	.a(north_input_NIB_storage_data_f_3__27_),
	.b(n25836));
   na02f01 U25285 (.o(n21204),
	.a(north_input_NIB_storage_data_f_3__26_),
	.b(n25836));
   oa12f01 U25286 (.o(n13248),
	.a(n21204),
	.b(n25836),
	.c(n21266));
   na02f01 U25287 (.o(n21205),
	.a(north_input_NIB_storage_data_f_3__34_),
	.b(n25836));
   oa12f01 U25288 (.o(n13208),
	.a(n21205),
	.b(n25836),
	.c(n22648));
   na02f01 U25289 (.o(n21206),
	.a(north_input_NIB_storage_data_f_3__37_),
	.b(n25836));
   oa12f01 U25290 (.o(n13193),
	.a(n21206),
	.b(n25836),
	.c(n22654));
   na02f01 U25291 (.o(n21207),
	.a(north_input_NIB_storage_data_f_3__24_),
	.b(n25836));
   na02f01 U25292 (.o(n21208),
	.a(north_input_NIB_storage_data_f_3__31_),
	.b(n25836));
   oa12f01 U25293 (.o(n13223),
	.a(n21208),
	.b(n25836),
	.c(n21237));
   na02f01 U25294 (.o(n21209),
	.a(north_input_NIB_storage_data_f_3__35_),
	.b(n25836));
   oa12f01 U25295 (.o(n13203),
	.a(n21209),
	.b(n25836),
	.c(n22644));
   na02f01 U25296 (.o(n21210),
	.a(north_input_NIB_storage_data_f_3__23_),
	.b(n25836));
   na02f01 U25297 (.o(n21211),
	.a(north_input_NIB_storage_data_f_3__28_),
	.b(n25836));
   na02f01 U25298 (.o(n21212),
	.a(north_input_NIB_storage_data_f_3__36_),
	.b(n25836));
   oa12f01 U25299 (.o(n13198),
	.a(n21212),
	.b(n25836),
	.c(n22656));
   na02f01 U25300 (.o(n21213),
	.a(north_input_NIB_storage_data_f_3__29_),
	.b(n25836));
   oa12f01 U25301 (.o(n13233),
	.a(n21213),
	.b(n25836),
	.c(n21248));
   na02f01 U25302 (.o(n21214),
	.a(north_input_NIB_storage_data_f_3__50_),
	.b(n25836));
   oa12f01 U25303 (.o(n13128),
	.a(n21214),
	.b(n25836),
	.c(n21282));
   na02f01 U25304 (.o(n21215),
	.a(north_input_NIB_storage_data_f_3__30_),
	.b(n25836));
   oa12f01 U25305 (.o(n13228),
	.a(n21215),
	.b(n25836),
	.c(n21259));
   na02f01 U25306 (.o(n21216),
	.a(north_input_NIB_storage_data_f_3__32_),
	.b(n25836));
   oa12f01 U25307 (.o(n13218),
	.a(n21216),
	.b(n25836),
	.c(n22640));
   in01s01 U25308 (.o(n25829),
	.a(north_input_NIB_tail_ptr_f_0_));
   no02f01 U25309 (.o(n21217),
	.a(north_input_NIB_tail_ptr_f_1_),
	.b(n25829));
   na02f01 U25310 (.o(n21221),
	.a(north_input_NIB_storage_data_f_1__23_),
	.b(FE_OFN88_n21220));
   na02f01 U25311 (.o(n21225),
	.a(north_input_NIB_storage_data_f_1__22_),
	.b(FE_OFN88_n21220));
   na02f01 U25312 (.o(n21227),
	.a(north_input_NIB_storage_data_f_1__36_),
	.b(FE_OFN88_n21220));
   na02f01 U25313 (.o(n21229),
	.a(north_input_NIB_storage_data_f_1__61_),
	.b(n25848));
   na02f01 U25314 (.o(n21230),
	.a(north_input_NIB_storage_data_f_1__32_),
	.b(FE_OFN88_n21220));
   na02f01 U25315 (.o(n21231),
	.a(north_input_NIB_storage_data_f_1__25_),
	.b(FE_OFN88_n21220));
   na02f01 U25316 (.o(n21233),
	.a(north_input_NIB_storage_data_f_1__47_),
	.b(FE_OFN88_n21220));
   na02f01 U25317 (.o(n21235),
	.a(north_input_NIB_storage_data_f_1__42_),
	.b(FE_OFN88_n21220));
   na02f01 U25318 (.o(n21236),
	.a(north_input_NIB_storage_data_f_1__31_),
	.b(FE_OFN88_n21220));
   na02f01 U25319 (.o(n21238),
	.a(north_input_NIB_storage_data_f_1__51_),
	.b(n25848));
   na02f01 U25320 (.o(n21240),
	.a(north_input_NIB_storage_data_f_1__63_),
	.b(n25848));
   na02f01 U25321 (.o(n21242),
	.a(north_input_NIB_storage_data_f_1__28_),
	.b(FE_OFN88_n21220));
   na02f01 U25322 (.o(n21244),
	.a(north_input_NIB_storage_data_f_1__46_),
	.b(FE_OFN88_n21220));
   na02f01 U25323 (.o(n21245),
	.a(north_input_NIB_storage_data_f_1__62_),
	.b(n25848));
   na02f01 U25324 (.o(n21247),
	.a(north_input_NIB_storage_data_f_1__29_),
	.b(FE_OFN88_n21220));
   na02f01 U25325 (.o(n21249),
	.a(north_input_NIB_storage_data_f_1__27_),
	.b(FE_OFN88_n21220));
   na02f01 U25326 (.o(n21251),
	.a(north_input_NIB_storage_data_f_1__59_),
	.b(n25848));
   na02f01 U25327 (.o(n21252),
	.a(north_input_NIB_storage_data_f_1__35_),
	.b(FE_OFN88_n21220));
   na02f01 U25328 (.o(n21253),
	.a(north_input_NIB_storage_data_f_1__55_),
	.b(n25848));
   na02f01 U25329 (.o(n21255),
	.a(north_input_NIB_storage_data_f_1__58_),
	.b(n25848));
   na02f01 U25330 (.o(n21257),
	.a(north_input_NIB_storage_data_f_1__37_),
	.b(FE_OFN88_n21220));
   na02f01 U25331 (.o(n21258),
	.a(north_input_NIB_storage_data_f_1__30_),
	.b(FE_OFN88_n21220));
   na02f01 U25332 (.o(n21260),
	.a(north_input_NIB_storage_data_f_1__34_),
	.b(FE_OFN88_n21220));
   na02f01 U25333 (.o(n21261),
	.a(north_input_NIB_storage_data_f_1__40_),
	.b(FE_OFN88_n21220));
   na02f01 U25334 (.o(n21263),
	.a(north_input_NIB_storage_data_f_1__41_),
	.b(FE_OFN88_n21220));
   na02f01 U25335 (.o(n21265),
	.a(north_input_NIB_storage_data_f_1__26_),
	.b(FE_OFN88_n21220));
   na02f01 U25336 (.o(n21267),
	.a(north_input_NIB_storage_data_f_1__48_),
	.b(FE_OFN88_n21220));
   na02f01 U25337 (.o(n21268),
	.a(north_input_NIB_storage_data_f_1__38_),
	.b(FE_OFN88_n21220));
   na02f01 U25338 (.o(n21271),
	.a(north_input_NIB_storage_data_f_1__44_),
	.b(FE_OFN88_n21220));
   na02f01 U25339 (.o(n21273),
	.a(north_input_NIB_storage_data_f_1__57_),
	.b(n25848));
   na02f01 U25340 (.o(n21275),
	.a(north_input_NIB_storage_data_f_1__45_),
	.b(FE_OFN88_n21220));
   na02f01 U25341 (.o(n21276),
	.a(north_input_NIB_storage_data_f_1__56_),
	.b(n25848));
   na02f01 U25342 (.o(n21278),
	.a(north_input_NIB_storage_data_f_1__49_),
	.b(FE_OFN88_n21220));
   na02f01 U25343 (.o(n21279),
	.a(north_input_NIB_storage_data_f_1__52_),
	.b(n25848));
   na02f01 U25344 (.o(n21281),
	.a(north_input_NIB_storage_data_f_1__50_),
	.b(FE_OFN88_n21220));
   na02f01 U25345 (.o(n21283),
	.a(north_input_NIB_storage_data_f_1__43_),
	.b(FE_OFN88_n21220));
   na02f01 U25346 (.o(n21284),
	.a(north_input_NIB_storage_data_f_1__53_),
	.b(FE_OFN88_n21220));
   na02f01 U25347 (.o(n21286),
	.a(north_input_NIB_storage_data_f_1__60_),
	.b(n25848));
   na03f02 U25348 (.o(dataOut_E_50_),
	.a(n21292),
	.b(n21291),
	.c(n21290));
   na03m02 U25350 (.o(dataOut_E_63_),
	.a(n21298),
	.b(n21297),
	.c(n21296));
   ao22f01 U25351 (.o(n21302),
	.a(n18077),
	.b(proc_input_NIB_storage_data_f_5__5_),
	.c(FE_OFN20_n17779),
	.d(proc_input_NIB_storage_data_f_7__5_));
   ao22f02 U25352 (.o(n21301),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__5_),
	.c(FE_OCPN25834_n),
	.d(proc_input_NIB_storage_data_f_0__5_));
   ao22f01 U25353 (.o(n21300),
	.a(n19709),
	.b(proc_input_NIB_storage_data_f_3__5_),
	.c(FE_OFN25604_n19530),
	.d(proc_input_NIB_storage_data_f_13__5_));
   ao22f01 U25354 (.o(n21299),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__5_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__5_));
   ao22f01 U25355 (.o(n21306),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__5_),
	.c(n17743),
	.d(proc_input_NIB_storage_data_f_4__5_));
   ao22f01 U25356 (.o(n21305),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__5_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__5_));
   ao22f01 U25357 (.o(n21304),
	.a(FE_OFN25635_n19595),
	.b(proc_input_NIB_storage_data_f_15__5_),
	.c(FE_RN_51),
	.d(proc_input_NIB_storage_data_f_1__5_));
   ao22f01 U25358 (.o(n21303),
	.a(n24060),
	.b(proc_input_NIB_storage_data_f_9__5_),
	.c(FE_OFN25645_n21748),
	.d(proc_input_NIB_storage_data_f_8__5_));
   ao22f01 U25359 (.o(n21310),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__5_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__5_));
   ao22f01 U25360 (.o(n21309),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__5_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__5_));
   na02f03 U25361 (.o(n23974),
	.a(n21310),
	.b(n21309));
   ao22f01 U25362 (.o(n21312),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__5_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__5_));
   ao22f01 U25363 (.o(n21311),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__5_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__5_));
   na02f02 U25364 (.o(n23975),
	.a(n21312),
	.b(n21311));
   ao22f01 U25365 (.o(n21314),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__5_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__5_));
   ao22f01 U25366 (.o(n21313),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__5_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__5_));
   na02f03 U25367 (.o(n23977),
	.a(n21314),
	.b(n21313));
   ao22f01 U25368 (.o(n21316),
	.a(FE_RN_17),
	.b(south_input_NIB_storage_data_f_2__5_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__5_));
   na02f02 U25369 (.o(n23976),
	.a(n21317),
	.b(n21316));
   na02f02 U25370 (.o(n21320),
	.a(n21319),
	.b(n21318));
   in01s01 U25371 (.o(n21321),
	.a(n21320));
   ao22f01 U25372 (.o(n21323),
	.a(n19019),
	.b(n23975),
	.c(n19017),
	.d(n23974));
   na03f02 U25374 (.o(dataOut_N_63_),
	.a(n21328),
	.b(n21327),
	.c(n21326));
   na03f02 U25375 (.o(dataOut_N_50_),
	.a(n21331),
	.b(n21330),
	.c(n21329));
   na02f01 U25377 (.o(n21336),
	.a(n21335),
	.b(n21334));
   na02f01 U25379 (.o(n21340),
	.a(n21339),
	.b(n21338));
   na03f04 U25380 (.o(dataOut_E_45_),
	.a(n21345),
	.b(n21344),
	.c(n21343));
   na03f04 U25381 (.o(dataOut_N_45_),
	.a(n21348),
	.b(n21347),
	.c(n21346));
   ao22f01 U25382 (.o(n21352),
	.a(n18077),
	.b(proc_input_NIB_storage_data_f_5__6_),
	.c(FE_OFN20_n17779),
	.d(proc_input_NIB_storage_data_f_7__6_));
   ao22f01 U25383 (.o(n21351),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__6_),
	.c(FE_OCPN25834_n),
	.d(proc_input_NIB_storage_data_f_0__6_));
   ao22f01 U25384 (.o(n21350),
	.a(n24454),
	.b(proc_input_NIB_storage_data_f_13__6_),
	.c(FE_RN_51),
	.d(proc_input_NIB_storage_data_f_1__6_));
   ao22f01 U25385 (.o(n21349),
	.a(n17754),
	.b(proc_input_NIB_storage_data_f_3__6_),
	.c(FE_OCPN25954_n18039),
	.d(proc_input_NIB_storage_data_f_10__6_));
   ao22f01 U25386 (.o(n21356),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__6_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__6_));
   ao22f01 U25387 (.o(n21355),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__6_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__6_));
   ao22f01 U25388 (.o(n21354),
	.a(FE_OFN25635_n19595),
	.b(proc_input_NIB_storage_data_f_15__6_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__6_));
   ao22f01 U25389 (.o(n21353),
	.a(n24060),
	.b(proc_input_NIB_storage_data_f_9__6_),
	.c(FE_OFN25645_n21748),
	.d(proc_input_NIB_storage_data_f_8__6_));
   ao22f01 U25390 (.o(n21360),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__6_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__6_));
   ao22f01 U25391 (.o(n21359),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__6_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__6_));
   na02f02 U25392 (.o(n24010),
	.a(n21360),
	.b(n21359));
   ao22f01 U25393 (.o(n21362),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__6_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__6_));
   ao22f01 U25394 (.o(n21361),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__6_),
	.c(FE_RN_27),
	.d(west_input_NIB_storage_data_f_1__6_));
   na02f02 U25395 (.o(n24011),
	.a(n21362),
	.b(n21361));
   ao22f01 U25396 (.o(n21364),
	.a(FE_OFN24771_n19075),
	.b(north_input_NIB_storage_data_f_0__6_),
	.c(n19220),
	.d(north_input_NIB_storage_data_f_2__6_));
   ao22f01 U25397 (.o(n21363),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__6_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__6_));
   na02f02 U25398 (.o(n24013),
	.a(n21364),
	.b(n21363));
   ao22f01 U25399 (.o(n21367),
	.a(FE_RN_13),
	.b(south_input_NIB_storage_data_f_3__6_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__6_));
   ao22f01 U25400 (.o(n21366),
	.a(n21365),
	.b(south_input_NIB_storage_data_f_2__6_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__6_));
   na02f02 U25401 (.o(n24012),
	.a(n21367),
	.b(n21366));
   na02f02 U25402 (.o(n21370),
	.a(n21369),
	.b(n21368));
   in01f01 U25403 (.o(n21371),
	.a(n21370));
   na03f03 U25405 (.o(dataOut_E_47_),
	.a(n21378),
	.b(n21377),
	.c(n21376));
   no02f01 U25406 (.o(west_input_control_N46),
	.a(FE_OFN25647_reset),
	.b(n21383));
   oa12s01 U25407 (.o(n21389),
	.a(south_input_control_count_f_3_),
	.b(south_input_control_count_f_2_),
	.c(n21384));
   no02s01 U25408 (.o(n21386),
	.a(south_input_control_count_f_3_),
	.b(south_input_control_count_f_2_));
   na02f02 U25409 (.o(n23309),
	.a(n21386),
	.b(n21385));
   in01s01 U25410 (.o(n21387),
	.a(n23309));
   na02s01 U25411 (.o(n21388),
	.a(south_input_control_thanks_all_f),
	.b(n21387));
   ao12s01 U25412 (.o(n21390),
	.a(n25247),
	.b(n21389),
	.c(n21388));
   no02f01 U25413 (.o(south_input_control_N44),
	.a(FE_OFN5_reset),
	.b(n21391));
   na03f03 U25414 (.o(dataOut_N_47_),
	.a(n21394),
	.b(n21393),
	.c(n21392));
   na02f02 U25415 (.o(n21397),
	.a(n21396),
	.b(n21395));
   in01f01 U25417 (.o(n21402),
	.a(n21401));
   na03f06 U25418 (.o(dataOut_E_44_),
	.a(n21406),
	.b(n21405),
	.c(n21404));
   no02f01 U25419 (.o(n21411),
	.a(n21410),
	.b(n21409));
   na03f06 U25420 (.o(dataOut_N_44_),
	.a(n21414),
	.b(n21413),
	.c(n21412));
   oa22f01 U25421 (.o(n21417),
	.a(n21615),
	.b(n21673),
	.c(n23589),
	.d(FE_OFN565_n25385));
   no02f01 U25422 (.o(n21419),
	.a(n21418),
	.b(n21417));
   oa12f02 U25423 (.o(dataOut_E_58_),
	.a(n21419),
	.b(FE_OFN134_n23594),
	.c(FE_OFN25895_n25395));
   oa22f01 U25424 (.o(n21420),
	.a(n21615),
	.b(n21662),
	.c(n23589),
	.d(FE_OFN563_n25120));
   no02f01 U25425 (.o(n21422),
	.a(FE_OFN408_n21421),
	.b(n21420));
   oa12f02 U25426 (.o(dataOut_N_58_),
	.a(n21422),
	.b(FE_OFN134_n23594),
	.c(n21666));
   oa22f01 U25427 (.o(n21423),
	.a(n21615),
	.b(FE_OFN525_n24731),
	.c(n23589),
	.d(n22772));
   no02f01 U25428 (.o(n21425),
	.a(n21424),
	.b(n21423));
   oa12f02 U25429 (.o(dataOut_W_58_),
	.a(n21425),
	.b(FE_OFN134_n23594),
	.c(FE_OFN25878_n19446));
   in01s01 U25430 (.o(n21433),
	.a(n21430));
   oa22f01 U25431 (.o(n21432),
	.a(FE_OFN483_n23987),
	.b(FE_OFN565_n25385),
	.c(n23986),
	.d(n21673));
   oa22f01 U25433 (.o(n21436),
	.a(FE_OFN483_n23987),
	.b(FE_OFN563_n25120),
	.c(n23986),
	.d(n21662));
   no02f01 U25434 (.o(n21438),
	.a(n21437),
	.b(n21436));
   oa12f02 U25435 (.o(dataOut_N_22_),
	.a(n21438),
	.b(FE_OFN144_n23991),
	.c(FE_OFN25869_n21666));
   na03f03 U25436 (.o(dataOut_N_46_),
	.a(n21441),
	.b(n21440),
	.c(n21439));
   na02f01 U25437 (.o(n21447),
	.a(n21446),
	.b(n21445));
   in01s01 U25438 (.o(n21448),
	.a(n21447));
   in01s01 U25439 (.o(n21452),
	.a(n21451));
   no02f01 U25440 (.o(n21455),
	.a(n21454),
	.b(n21453));
   no02f01 U25441 (.o(n21458),
	.a(n21457),
	.b(n21456));
   in01f01 U25442 (.o(n23478),
	.a(n25003));
   ao22f01 U25443 (.o(n21460),
	.a(n19017),
	.b(n23478),
	.c(n19020),
	.d(n23480));
   na03f02 U25444 (.o(dataOut_E_30_),
	.a(n21461),
	.b(n21460),
	.c(n21459));
   na03f02 U25445 (.o(dataOut_N_30_),
	.a(n21464),
	.b(n21463),
	.c(n21462));
   na03f02 U25446 (.o(dataOut_N_53_),
	.a(n21468),
	.b(n21467),
	.c(n21466));
   in01f01 U25447 (.o(n23495),
	.a(n21471));
   na03f01 U25448 (.o(FE_OFN352_dataOut_E_43),
	.a(n21474),
	.b(n21473),
	.c(n21472));
   na03f01 U25449 (.o(FE_OFN288_dataOut_N_43),
	.a(n21477),
	.b(n21476),
	.c(n21475));
   na03f02 U25450 (.o(dataOut_E_55_),
	.a(n21488),
	.b(n21487),
	.c(n21486));
   na03f02 U25451 (.o(dataOut_N_55_),
	.a(n21491),
	.b(n21490),
	.c(n21489));
   no02f01 U25452 (.o(n21499),
	.a(n21497),
	.b(n21496));
   na02f01 U25453 (.o(FE_OFN354_dataOut_E_40),
	.a(n21499),
	.b(n21498));
   no02f01 U25454 (.o(n21503),
	.a(n21501),
	.b(n21500));
   na02f01 U25455 (.o(FE_OFN360_dataOut_S_40),
	.a(n21503),
	.b(n21502));
   no02f01 U25456 (.o(n21507),
	.a(n21505),
	.b(n21504));
   na02f01 U25457 (.o(FE_OFN0_dataOut_N_40),
	.a(n21507),
	.b(n21506));
   no02f01 U25458 (.o(n21512),
	.a(n21511),
	.b(n21510));
   oa12f01 U25459 (.o(dataOut_E_61_),
	.a(n21512),
	.b(n24009),
	.c(FE_OFN25895_n25395));
   no02f01 U25460 (.o(n21515),
	.a(n21514),
	.b(n21513));
   oa12f01 U25461 (.o(dataOut_N_61_),
	.a(n21515),
	.b(n24009),
	.c(n21666));
   ao22f01 U25462 (.o(n21517),
	.a(n19017),
	.b(n23527),
	.c(n19022),
	.d(n23526));
   na03f04 U25463 (.o(dataOut_E_26_),
	.a(n21518),
	.b(n21517),
	.c(n21516));
   na03f04 U25464 (.o(dataOut_N_26_),
	.a(n21521),
	.b(n21520),
	.c(n21519));
   no02f01 U25465 (.o(n21530),
	.a(n21528),
	.b(n21527));
   na02f01 U25466 (.o(dataOut_E_41_),
	.a(n21530),
	.b(n21529));
   no02f01 U25467 (.o(n21534),
	.a(n21532),
	.b(n21531));
   na02f02 U25468 (.o(dataOut_S_41_),
	.a(n21534),
	.b(n21533));
   no04f01 U25469 (.o(n21535),
	.a(west_input_control_count_f_2_),
	.b(west_input_control_count_f_3_),
	.c(west_input_control_count_f_5_),
	.d(west_input_control_count_f_4_));
   in01s01 U25470 (.o(n21536),
	.a(n21535));
   no03s01 U25471 (.o(n21537),
	.a(west_input_control_count_f_7_),
	.b(west_input_control_count_f_6_),
	.c(n21536));
   in01s01 U25472 (.o(n21540),
	.a(n26012));
   no02f01 U25473 (.o(west_input_control_N52),
	.a(FE_OFN91_n21590),
	.b(n21540));
   no02f01 U25474 (.o(n21544),
	.a(n21542),
	.b(n21541));
   na02f02 U25475 (.o(dataOut_N_41_),
	.a(n21544),
	.b(n21543));
   in01f01 U25476 (.o(n21547),
	.a(n21545));
   no02f01 U25477 (.o(n21551),
	.a(n21550),
	.b(n21549));
   no02f01 U25478 (.o(west_input_control_N53),
	.a(reset),
	.b(n25028));
   ao22f01 U25479 (.o(n21553),
	.a(n19017),
	.b(n23534),
	.c(n19020),
	.d(n23535));
   na03f04 U25480 (.o(dataOut_E_25_),
	.a(n21554),
	.b(n21553),
	.c(n21552));
   na03m02 U25481 (.o(FE_OFN312_dataOut_N_25),
	.a(n21557),
	.b(n21556),
	.c(n21555));
   in01f01 U25482 (.o(n23517),
	.a(n21558));
   ao22f01 U25483 (.o(n21561),
	.a(n19019),
	.b(n23517),
	.c(n19020),
	.d(n23516));
   ao22f01 U25484 (.o(n21560),
	.a(n19017),
	.b(n23519),
	.c(n19022),
	.d(n23518));
   na03m02 U25485 (.o(FE_OFN627_dataOut_E_27),
	.a(n21561),
	.b(n21560),
	.c(n21559));
   na03f01 U25486 (.o(FE_OFN595_dataOut_N_27),
	.a(n21564),
	.b(n21563),
	.c(n21562));
   in01s01 U25487 (.o(n21588),
	.a(n21565));
   in01s01 U25488 (.o(n21583),
	.a(east_input_control_count_f_2_));
   in01s01 U25489 (.o(n21566),
	.a(east_input_control_count_f_3_));
   ao12s01 U25490 (.o(n21567),
	.a(n21566),
	.b(n21584),
	.c(n21583));
   no02s01 U25491 (.o(n21568),
	.a(n21577),
	.b(n21567));
   oa22f01 U25492 (.o(east_input_control_N44),
	.a(n21569),
	.b(n21588),
	.c(n21568),
	.d(FE_OFN906_n21586));
   in01s01 U25493 (.o(n21575),
	.a(n23959));
   in01s01 U25494 (.o(n21585),
	.a(n21584));
   na02s01 U25495 (.o(n21571),
	.a(n21902),
	.b(n21570));
   no02s01 U25496 (.o(n21572),
	.a(n21585),
	.b(n21571));
   in01s01 U25497 (.o(n21573),
	.a(n21572));
   in01s01 U25498 (.o(n21901),
	.a(east_input_control_count_f_7_));
   na02s01 U25499 (.o(n21580),
	.a(n21577),
	.b(n21576));
   in01s01 U25500 (.o(n21579),
	.a(n21580));
   in01s01 U25501 (.o(n21578),
	.a(east_input_control_count_f_5_));
   ao22m01 U25502 (.o(n21581),
	.a(east_input_control_count_f_5_),
	.b(n21580),
	.c(n21579),
	.d(n21578));
   oa22f01 U25503 (.o(east_input_control_N46),
	.a(n21582),
	.b(n21588),
	.c(n21581),
	.d(FE_OFN906_n21586));
   ao22s01 U25504 (.o(n21587),
	.a(east_input_control_count_f_2_),
	.b(n21585),
	.c(n21584),
	.d(n21583));
   oa22s01 U25505 (.o(east_input_control_N43),
	.a(n21589),
	.b(n21588),
	.c(n21587),
	.d(FE_OFN906_n21586));
   ao12f01 U25506 (.o(west_input_control_N51),
	.a(n26012),
	.b(FE_OFN91_n21590),
	.c(FE_OFN25598_reset));
   no02f01 U25507 (.o(n21593),
	.a(n21592),
	.b(n21591));
   oa12f01 U25508 (.o(FE_OFN683_dataOut_S_38),
	.a(n21593),
	.b(n18031),
	.c(FE_OFN266_n25499));
   no02f01 U25509 (.o(n21596),
	.a(n21595),
	.b(n21594));
   no02f01 U25510 (.o(n21599),
	.a(n21598),
	.b(n21597));
   no02f01 U25511 (.o(n21608),
	.a(n21607),
	.b(n21606));
   no02f01 U25512 (.o(n21611),
	.a(n21610),
	.b(n21609));
   no02f01 U25513 (.o(n21614),
	.a(n21613),
	.b(n21612));
   no02f01 U25514 (.o(n21619),
	.a(n21618),
	.b(n21617));
   oa12f02 U25515 (.o(dataOut_S_58_),
	.a(n21619),
	.b(FE_OFN134_n23594),
	.c(FE_OFN25652_n25499));
   no02f01 U25516 (.o(n21622),
	.a(n21621),
	.b(n21620));
   no02f02 U25517 (.o(n21625),
	.a(n21624),
	.b(n21623));
   no02f01 U25518 (.o(n21628),
	.a(n21627),
	.b(n21626));
   oa12f02 U25519 (.o(dataOut_S_61_),
	.a(n21628),
	.b(n24009),
	.c(FE_OFN25652_n25499));
   no02f01 U25520 (.o(n21631),
	.a(n21630),
	.b(n21629));
   ao22f01 U25521 (.o(n21632),
	.a(n19493),
	.b(n23984),
	.c(FE_OFN105_n22517),
	.d(n23983));
   in01s01 U25522 (.o(n21634),
	.a(n21632));
   oa12f01 U25523 (.o(FE_OFN709_dataOut_S_22),
	.a(n21635),
	.b(FE_OFN144_n23991),
	.c(FE_OFN25651_n25499));
   no02f01 U25524 (.o(n21683),
	.a(proc_input_control_count_f_0_),
	.b(proc_input_control_count_f_1_));
   in01f01 U25525 (.o(n21677),
	.a(n21683));
   no02f01 U25526 (.o(n21658),
	.a(n21688),
	.b(n21677));
   in01s01 U25527 (.o(n21636),
	.a(proc_input_control_count_f_2_));
   na02f01 U25528 (.o(n21678),
	.a(n21658),
	.b(n21636));
   in01s01 U25529 (.o(n21637),
	.a(proc_input_control_count_f_3_));
   na02f02 U25530 (.o(n21647),
	.a(n21638),
	.b(n21637));
   no02f02 U25531 (.o(n21651),
	.a(proc_input_control_count_f_4_),
	.b(n21647));
   in01s01 U25532 (.o(n21639),
	.a(proc_input_control_count_f_5_));
   ao22f01 U25533 (.o(n21641),
	.a(proc_input_control_count_f_5_),
	.b(n21640),
	.c(n21651),
	.d(n21639));
   na02f01 U25534 (.o(n21643),
	.a(proc_input_control_count_f_3_),
	.b(n21678));
   in01s01 U25535 (.o(n21645),
	.a(n21644));
   ao12f01 U25536 (.o(n21648),
	.a(n21651),
	.b(proc_input_control_count_f_4_),
	.c(n21647));
   na02f01 U25537 (.o(n21654),
	.a(n21651),
	.b(n21650));
   in01f01 U25538 (.o(n21653),
	.a(n21654));
   in01s01 U25539 (.o(n21652),
	.a(proc_input_control_count_f_7_));
   oa22f01 U25540 (.o(proc_input_control_N48),
	.a(n23964),
	.b(n21694),
	.c(n21655),
	.d(n21689));
   in01f01 U25541 (.o(n21656),
	.a(proc_input_control_count_f_1_));
   no02s01 U25542 (.o(n21659),
	.a(n21657),
	.b(n21656));
   oa22f01 U25543 (.o(proc_input_control_N42),
	.a(n23628),
	.b(n21694),
	.c(n22899),
	.d(n21689));
   in01f01 U25544 (.o(n24000),
	.a(n18120));
   no02s01 U25545 (.o(n21665),
	.a(n21664),
	.b(n21663));
   oa12f01 U25546 (.o(dataOut_N_54_),
	.a(n21665),
	.b(n24000),
	.c(FE_OFN25977_n21666));
   no02f01 U25547 (.o(n21670),
	.a(n21669),
	.b(n21668));
   oa12f01 U25548 (.o(dataOut_S_54_),
	.a(n21670),
	.b(n24000),
	.c(FE_OFN25652_n25499));
   no02f01 U25549 (.o(n21676),
	.a(n21675),
	.b(n21674));
   oa12f01 U25550 (.o(dataOut_E_54_),
	.a(n21676),
	.b(n24000),
	.c(FE_OFN25895_n25395));
   oa12f01 U25551 (.o(n21679),
	.a(proc_input_control_count_f_2_),
	.b(n21677),
	.c(n21688));
   no02f01 U25552 (.o(proc_input_control_N43),
	.a(FE_OFN8_reset),
	.b(n21682));
   no04f01 U25553 (.o(n22898),
	.a(proc_input_control_count_f_5_),
	.b(proc_input_control_count_f_4_),
	.c(proc_input_control_count_f_3_),
	.d(proc_input_control_count_f_2_));
   in01s01 U25554 (.o(n21686),
	.a(proc_input_control_count_f_6_));
   na02s01 U25555 (.o(n21684),
	.a(proc_input_control_thanks_all_f),
	.b(FE_OFN574_n25463));
   oa12s01 U25556 (.o(n21691),
	.a(n21685),
	.b(n21687),
	.c(n21686));
   na02s01 U25557 (.o(n21690),
	.a(proc_input_control_count_f_6_),
	.b(n21688));
   in01s01 U25558 (.o(n21693),
	.a(n21692));
   oa12f01 U25559 (.o(proc_input_control_N47),
	.a(n21693),
	.b(n23956),
	.c(n21694));
   na03m02 U25560 (.o(dataOut_W_51_),
	.a(n21699),
	.b(n21698),
	.c(n21697));
   na03f03 U25561 (.o(dataOut_W_47_),
	.a(n21702),
	.b(n21701),
	.c(n21700));
   na03f04 U25562 (.o(dataOut_W_45_),
	.a(n21705),
	.b(n21704),
	.c(n21703));
   na03f02 U25563 (.o(dataOut_W_30_),
	.a(n21708),
	.b(n21707),
	.c(n21706));
   na03f04 U25564 (.o(dataOut_W_44_),
	.a(n21711),
	.b(n21710),
	.c(n21709));
   na03f02 U25565 (.o(dataOut_W_55_),
	.a(n21714),
	.b(n21713),
	.c(n21712));
   na03f02 U25566 (.o(dataOut_W_50_),
	.a(n21717),
	.b(n21716),
	.c(n21715));
   na03m02 U25567 (.o(dataOut_W_63_),
	.a(n21720),
	.b(n21719),
	.c(n21718));
   ao22f01 U25568 (.o(n21722),
	.a(n17755),
	.b(n23535),
	.c(FE_OFN526_n24731),
	.d(n23534));
   na03f02 U25569 (.o(FE_OFN779_dataOut_W_25),
	.a(n21723),
	.b(n21722),
	.c(n21721));
   na03f04 U25570 (.o(dataOut_W_43_),
	.a(n21729),
	.b(n21728),
	.c(n21727));
   ao22f01 U25571 (.o(n21735),
	.a(n17786),
	.b(n23517),
	.c(n17755),
	.d(n23516));
   ao22f01 U25572 (.o(n21734),
	.a(FE_OFN111_n22773),
	.b(n23519),
	.c(FE_OFN94_n21695),
	.d(n23518));
   na03m02 U25573 (.o(FE_OFN775_dataOut_W_27),
	.a(n21735),
	.b(n21734),
	.c(n21733));
   ao22f01 U25574 (.o(n21737),
	.a(FE_OFN111_n22773),
	.b(n23527),
	.c(FE_OFN94_n21695),
	.d(n23526));
   na03f04 U25575 (.o(dataOut_W_26_),
	.a(n21738),
	.b(n21737),
	.c(n21736));
   ao22f01 U25576 (.o(n21744),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__8_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__8_));
   ao22f01 U25577 (.o(n21743),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__8_),
	.c(FE_OCPN25834_n),
	.d(proc_input_NIB_storage_data_f_0__8_));
   ao22f01 U25578 (.o(n21741),
	.a(n20056),
	.b(proc_input_NIB_storage_data_f_9__8_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__8_));
   ao22f01 U25579 (.o(n21753),
	.a(FE_OCPN25814_FE_OFN186_n24453),
	.b(proc_input_NIB_storage_data_f_2__8_),
	.c(FE_OCPN25954_n18039),
	.d(proc_input_NIB_storage_data_f_10__8_));
   ao22f01 U25580 (.o(n21752),
	.a(n18077),
	.b(proc_input_NIB_storage_data_f_5__8_),
	.c(FE_OFN25692_n19503),
	.d(proc_input_NIB_storage_data_f_6__8_));
   ao22f01 U25581 (.o(n21751),
	.a(FE_OFN25635_n19595),
	.b(proc_input_NIB_storage_data_f_15__8_),
	.c(FE_RN_51),
	.d(proc_input_NIB_storage_data_f_1__8_));
   ao22f01 U25582 (.o(n21750),
	.a(FE_OFN168_n24343),
	.b(proc_input_NIB_storage_data_f_8__8_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__8_));
   ao22f01 U25584 (.o(n21756),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__8_),
	.c(FE_RN_27),
	.d(west_input_NIB_storage_data_f_1__8_));
   na02f04 U25585 (.o(n23147),
	.a(n21757),
	.b(n21756));
   ao22f01 U25586 (.o(n21759),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__8_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__8_));
   ao22m02 U25587 (.o(n21758),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__8_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__8_));
   na02f04 U25588 (.o(n23146),
	.a(n21759),
	.b(n21758));
   ao22f01 U25589 (.o(n21761),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__8_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__8_));
   ao22f01 U25590 (.o(n21760),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__8_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__8_));
   na02f02 U25591 (.o(n23148),
	.a(n21761),
	.b(n21760));
   ao22f01 U25592 (.o(n21763),
	.a(n24472),
	.b(south_input_NIB_storage_data_f_0__8_),
	.c(n17782),
	.d(south_input_NIB_storage_data_f_2__8_));
   ao22f01 U25593 (.o(n21762),
	.a(FE_RN_13),
	.b(south_input_NIB_storage_data_f_3__8_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__8_));
   na02f02 U25594 (.o(n23149),
	.a(n21763),
	.b(n21762));
   na02f02 U25595 (.o(n21766),
	.a(n21765),
	.b(n21764));
   in01s01 U25596 (.o(n21767),
	.a(n21766));
   ao22f01 U25597 (.o(n21772),
	.a(n18077),
	.b(proc_input_NIB_storage_data_f_5__10_),
	.c(FE_OFN20_n17779),
	.d(proc_input_NIB_storage_data_f_7__10_));
   ao22m02 U25598 (.o(n21770),
	.a(FE_OFN25691_n19503),
	.b(proc_input_NIB_storage_data_f_6__10_),
	.c(n19709),
	.d(proc_input_NIB_storage_data_f_3__10_));
   ao22f01 U25599 (.o(n21769),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__10_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__10_));
   ao22f01 U25600 (.o(n21776),
	.a(n24454),
	.b(proc_input_NIB_storage_data_f_13__10_),
	.c(FE_OFN25645_n21748),
	.d(proc_input_NIB_storage_data_f_8__10_));
   ao22f01 U25601 (.o(n21775),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__10_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__10_));
   ao22f01 U25602 (.o(n21774),
	.a(FE_OFN25635_n19595),
	.b(proc_input_NIB_storage_data_f_15__10_),
	.c(FE_RN_51),
	.d(proc_input_NIB_storage_data_f_1__10_));
   ao22f01 U25603 (.o(n21773),
	.a(n24060),
	.b(proc_input_NIB_storage_data_f_9__10_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__10_));
   ao22f01 U25604 (.o(n21780),
	.a(FE_OCPN25938_n24965),
	.b(south_input_NIB_storage_data_f_3__10_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__10_));
   ao22f01 U25605 (.o(n21779),
	.a(n21365),
	.b(south_input_NIB_storage_data_f_2__10_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__10_));
   na02m02 U25606 (.o(n23577),
	.a(n21780),
	.b(n21779));
   ao22f01 U25607 (.o(n21782),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__10_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__10_));
   ao22f01 U25608 (.o(n21781),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__10_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__10_));
   na02f02 U25609 (.o(n23578),
	.a(n21782),
	.b(n21781));
   ao22f01 U25610 (.o(n21784),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__10_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__10_));
   ao22f01 U25611 (.o(n21783),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__10_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__10_));
   na02f04 U25612 (.o(n23580),
	.a(n21784),
	.b(n21783));
   ao22f01 U25613 (.o(n21786),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__10_),
	.c(FE_OFN24800_n20506),
	.d(east_input_NIB_storage_data_f_3__10_));
   ao22f01 U25614 (.o(n21785),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__10_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__10_));
   ao22f01 U25615 (.o(n21787),
	.a(n19019),
	.b(n23580),
	.c(n19017),
	.d(n23579));
   in01f01 U25616 (.o(n21790),
	.a(n21789));
   ao22f01 U25617 (.o(n21794),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__9_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__9_));
   ao22m02 U25618 (.o(n21793),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__9_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__9_));
   ao22f01 U25619 (.o(n21792),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__9_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__9_));
   ao22m02 U25620 (.o(n21791),
	.a(FE_OCPN25834_n),
	.b(proc_input_NIB_storage_data_f_0__9_),
	.c(FE_RN_51),
	.d(proc_input_NIB_storage_data_f_1__9_));
   ao22f01 U25621 (.o(n21799),
	.a(FE_OCPN25814_FE_OFN186_n24453),
	.b(proc_input_NIB_storage_data_f_2__9_),
	.c(n17754),
	.d(proc_input_NIB_storage_data_f_3__9_));
   ao22f01 U25622 (.o(n21798),
	.a(n18077),
	.b(proc_input_NIB_storage_data_f_5__9_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__9_));
   ao22f01 U25623 (.o(n21796),
	.a(n20056),
	.b(proc_input_NIB_storage_data_f_9__9_),
	.c(FE_OCPN25954_n18039),
	.d(proc_input_NIB_storage_data_f_10__9_));
   ao22f01 U25624 (.o(n21803),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__9_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__9_));
   ao22f01 U25625 (.o(n21802),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__9_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__9_));
   na02f03 U25626 (.o(n23569),
	.a(n21803),
	.b(n21802));
   ao22f01 U25627 (.o(n21805),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__9_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__9_));
   ao22f01 U25628 (.o(n21804),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__9_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__9_));
   na02f03 U25629 (.o(n23568),
	.a(n21805),
	.b(n21804));
   ao22f01 U25630 (.o(n21808),
	.a(FE_OFN24791_n24965),
	.b(south_input_NIB_storage_data_f_3__9_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__9_));
   ao22f01 U25631 (.o(n21807),
	.a(n24321),
	.b(south_input_NIB_storage_data_f_2__9_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__9_));
   na02f02 U25632 (.o(n23570),
	.a(n21808),
	.b(n21807));
   ao22f01 U25633 (.o(n21810),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__9_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__9_));
   ao22f01 U25634 (.o(n21809),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__9_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__9_));
   na02f04 U25635 (.o(n23571),
	.a(n21810),
	.b(n21809));
   na02f02 U25636 (.o(n21813),
	.a(n21812),
	.b(n21811));
   in01s01 U25637 (.o(n21814),
	.a(n21813));
   ao22f01 U25638 (.o(n21818),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__7_),
	.c(FE_OFN188_n24453),
	.d(proc_input_NIB_storage_data_f_2__7_));
   ao22f01 U25639 (.o(n21817),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__7_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__7_));
   ao22f01 U25640 (.o(n21816),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__7_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__7_));
   ao22f01 U25641 (.o(n21815),
	.a(FE_OCPN25834_n),
	.b(proc_input_NIB_storage_data_f_0__7_),
	.c(FE_OFN25645_n21748),
	.d(proc_input_NIB_storage_data_f_8__7_));
   ao22f01 U25642 (.o(n21822),
	.a(n24454),
	.b(proc_input_NIB_storage_data_f_13__7_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__7_));
   ao22f01 U25643 (.o(n21821),
	.a(n18077),
	.b(proc_input_NIB_storage_data_f_5__7_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__7_));
   ao22f01 U25644 (.o(n21820),
	.a(n17754),
	.b(proc_input_NIB_storage_data_f_3__7_),
	.c(FE_OFN165_n24129),
	.d(proc_input_NIB_storage_data_f_1__7_));
   ao22f01 U25645 (.o(n21819),
	.a(n20056),
	.b(proc_input_NIB_storage_data_f_9__7_),
	.c(FE_OCPN25954_n18039),
	.d(proc_input_NIB_storage_data_f_10__7_));
   ao22f01 U25646 (.o(n21826),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__7_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__7_));
   ao22f01 U25647 (.o(n21825),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__7_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__7_));
   na02f02 U25648 (.o(n23559),
	.a(n21826),
	.b(n21825));
   ao22f01 U25649 (.o(n21828),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__7_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__7_));
   ao22f01 U25650 (.o(n21827),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__7_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__7_));
   ao22f01 U25651 (.o(n21831),
	.a(FE_OFN28_n18974),
	.b(west_input_NIB_storage_data_f_0__7_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__7_));
   ao22f01 U25652 (.o(n21830),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__7_),
	.c(n24466),
	.d(west_input_NIB_storage_data_f_2__7_));
   na02f04 U25653 (.o(n23562),
	.a(n21831),
	.b(n21830));
   ao22f01 U25654 (.o(n21833),
	.a(FE_RN_13),
	.b(south_input_NIB_storage_data_f_3__7_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__7_));
   ao22f01 U25655 (.o(n21832),
	.a(FE_RN_17),
	.b(south_input_NIB_storage_data_f_2__7_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__7_));
   na02f02 U25656 (.o(n23561),
	.a(n21833),
	.b(n21832));
   ao22f01 U25657 (.o(n21834),
	.a(n19019),
	.b(n23562),
	.c(FE_OFN42_n19022),
	.d(n23561));
   na02f02 U25659 (.o(n21840),
	.a(n21839),
	.b(n21838));
   in01s01 U25660 (.o(n21841),
	.a(n21840));
   ao22f01 U25661 (.o(n21842),
	.a(FE_OFN44_n19054),
	.b(FE_OFN116_n23148),
	.c(FE_OFN366_n17753),
	.d(n23149));
   na02f02 U25662 (.o(n21844),
	.a(n21843),
	.b(n21842));
   ao22f01 U25664 (.o(n21850),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__33_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__33_));
   ao22m02 U25665 (.o(n21849),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__33_),
	.c(FE_OCPN25834_n),
	.d(proc_input_NIB_storage_data_f_0__33_));
   ao22f01 U25666 (.o(n21848),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__33_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__33_));
   ao22f01 U25667 (.o(n21847),
	.a(n21768),
	.b(proc_input_NIB_storage_data_f_3__33_),
	.c(n24060),
	.d(proc_input_NIB_storage_data_f_9__33_));
   ao22f01 U25668 (.o(n21853),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__33_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__33_));
   ao22f01 U25669 (.o(n21852),
	.a(FE_OFN25635_n19595),
	.b(proc_input_NIB_storage_data_f_15__33_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__33_));
   ao22f01 U25670 (.o(n21851),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__33_),
	.c(FE_OFN167_n24343),
	.d(proc_input_NIB_storage_data_f_8__33_));
   ao22f01 U25671 (.o(n21860),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__33_),
	.c(FE_OFN24800_n20506),
	.d(east_input_NIB_storage_data_f_3__33_));
   ao22f01 U25672 (.o(n21859),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__33_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__33_));
   ao22f01 U25673 (.o(n21863),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__33_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__33_));
   ao22f01 U25674 (.o(n21862),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__33_),
	.c(FE_RN_27),
	.d(west_input_NIB_storage_data_f_1__33_));
   na02f04 U25675 (.o(n24020),
	.a(n21863),
	.b(n21862));
   ao22f01 U25676 (.o(n21867),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__33_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__33_));
   ao22f01 U25677 (.o(n21866),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__33_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__33_));
   na02f02 U25678 (.o(n24022),
	.a(n21867),
	.b(n21866));
   ao22f01 U25679 (.o(n21869),
	.a(FE_RN_13),
	.b(south_input_NIB_storage_data_f_3__33_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__33_));
   ao22f01 U25680 (.o(n21868),
	.a(FE_RN_17),
	.b(south_input_NIB_storage_data_f_2__33_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__33_));
   na02f02 U25681 (.o(n24021),
	.a(n21869),
	.b(n21868));
   na02f02 U25682 (.o(n21872),
	.a(n21871),
	.b(n21870));
   in01s01 U25683 (.o(n21873),
	.a(n21872));
   ao22f01 U25684 (.o(n21875),
	.a(n19019),
	.b(n24020),
	.c(n19017),
	.d(FE_OFN151_n24019));
   na02f02 U25685 (.o(n21876),
	.a(n21875),
	.b(n21874));
   na02f02 U25687 (.o(n21880),
	.a(n21879),
	.b(n21878));
   ao22f01 U25689 (.o(n21882),
	.a(n19019),
	.b(n23571),
	.c(FE_OFN42_n19022),
	.d(n23570));
   in01f01 U25690 (.o(n21885),
	.a(n21884));
   in01s01 U25691 (.o(n21898),
	.a(n26009));
   no02s01 U25692 (.o(n21889),
	.a(north_input_control_count_f_5_),
	.b(north_input_control_count_f_7_));
   ao22s01 U25693 (.o(n21891),
	.a(n21889),
	.b(n21888),
	.c(n21887),
	.d(n21886));
   in01s01 U25694 (.o(n21909),
	.a(east_input_control_N41));
   ao22f01 U25695 (.o(n21905),
	.a(n21902),
	.b(n21901),
	.c(n21900),
	.d(n21899));
   no02m01 U25696 (.o(east_input_control_N52),
	.a(n21909),
	.b(n22083));
   in01s01 U25697 (.o(n23733),
	.a(proc_input_NIB_tail_ptr_f_2_));
   na02f01 U25698 (.o(n21912),
	.a(proc_input_NIB_storage_data_f_12__46_),
	.b(n21911));
   in01s01 U25699 (.o(n22137),
	.a(proc_input_NIB_tail_ptr_f_1_));
   na02s01 U25700 (.o(n21913),
	.a(proc_input_NIB_tail_ptr_f_0_),
	.b(n22137));
   na02f01 U25701 (.o(n21916),
	.a(proc_input_NIB_storage_data_f_13__59_),
	.b(FE_OFN25781_FE_OFN448_n23236));
   oa12f01 U25702 (.o(n7273),
	.a(n21916),
	.b(FE_OFN25781_FE_OFN448_n23236),
	.c(n23938));
   na02f01 U25703 (.o(n21917),
	.a(proc_input_NIB_storage_data_f_13__54_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   na02f01 U25704 (.o(n21918),
	.a(proc_input_NIB_storage_data_f_13__60_),
	.b(FE_OFN25781_FE_OFN448_n23236));
   oa12f01 U25705 (.o(n7268),
	.a(n21918),
	.b(FE_OFN25781_FE_OFN448_n23236),
	.c(n23926));
   na02f01 U25706 (.o(n21919),
	.a(proc_input_NIB_storage_data_f_13__57_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25707 (.o(n7283),
	.a(n21919),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23932));
   na02f01 U25708 (.o(n21920),
	.a(proc_input_NIB_storage_data_f_13__52_),
	.b(FE_OFN25781_FE_OFN448_n23236));
   oa12f01 U25709 (.o(n7308),
	.a(n21920),
	.b(FE_OFN25781_FE_OFN448_n23236),
	.c(n23890));
   na02f01 U25710 (.o(n21921),
	.a(proc_input_NIB_storage_data_f_13__53_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25711 (.o(n7303),
	.a(n21921),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23922));
   na02f01 U25712 (.o(n21922),
	.a(proc_input_NIB_storage_data_f_13__62_),
	.b(FE_OFN25781_FE_OFN448_n23236));
   oa12f01 U25713 (.o(n7258),
	.a(n21922),
	.b(FE_OFN25781_FE_OFN448_n23236),
	.c(n23810));
   na02f01 U25714 (.o(n21923),
	.a(proc_input_NIB_storage_data_f_13__55_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25715 (.o(n7293),
	.a(n21923),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23910));
   na02f01 U25716 (.o(n21924),
	.a(proc_input_NIB_storage_data_f_13__50_),
	.b(FE_OFN25781_FE_OFN448_n23236));
   na02f01 U25717 (.o(n21925),
	.a(proc_input_NIB_storage_data_f_13__56_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25718 (.o(n7288),
	.a(n21925),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23930));
   na02f01 U25719 (.o(n21926),
	.a(proc_input_NIB_storage_data_f_13__63_),
	.b(FE_OFN25781_FE_OFN448_n23236));
   na02f01 U25720 (.o(n21927),
	.a(proc_input_NIB_storage_data_f_13__58_),
	.b(FE_OFN25781_FE_OFN448_n23236));
   oa12f01 U25721 (.o(n7278),
	.a(n21927),
	.b(FE_OFN25781_FE_OFN448_n23236),
	.c(n23936));
   na02f01 U25722 (.o(n21928),
	.a(proc_input_NIB_storage_data_f_12__37_),
	.b(n21911));
   oa12f01 U25723 (.o(n7063),
	.a(n21928),
	.b(n21911),
	.c(n23796));
   na02f01 U25724 (.o(n21929),
	.a(proc_input_NIB_storage_data_f_13__48_),
	.b(n23236));
   oa12f01 U25725 (.o(n7328),
	.a(n21929),
	.b(n23236),
	.c(n23912));
   oa12f01 U25726 (.o(n7323),
	.a(n21930),
	.b(n23236),
	.c(n23908));
   na02f01 U25727 (.o(n21931),
	.a(proc_input_NIB_storage_data_f_13__61_),
	.b(FE_OFN25781_FE_OFN448_n23236));
   oa12f01 U25728 (.o(n7263),
	.a(n21931),
	.b(FE_OFN25781_FE_OFN448_n23236),
	.c(n23918));
   na02f01 U25729 (.o(n21932),
	.a(proc_input_NIB_storage_data_f_12__45_),
	.b(FE_OFN25627_n21910));
   oa12f01 U25730 (.o(n7023),
	.a(n21932),
	.b(FE_OFN25627_n21910),
	.c(n23942));
   oa12f01 U25731 (.o(n7028),
	.a(n21933),
	.b(FE_OFN25627_n21910),
	.c(n23920));
   na02f01 U25732 (.o(n21934),
	.a(proc_input_NIB_storage_data_f_12__47_),
	.b(FE_OFN914_n23246));
   oa12f01 U25733 (.o(n7013),
	.a(n21934),
	.b(FE_OFN914_n23246),
	.c(n23914));
   na02f01 U25734 (.o(n21935),
	.a(proc_input_NIB_storage_data_f_12__43_),
	.b(FE_OFN913_n23246));
   oa12f01 U25735 (.o(n7033),
	.a(n21935),
	.b(FE_OFN913_n23246),
	.c(n23806));
   na02f01 U25736 (.o(n21936),
	.a(proc_input_NIB_storage_data_f_12__48_),
	.b(n21911));
   oa12f01 U25737 (.o(n7008),
	.a(n21936),
	.b(n21911),
	.c(n23912));
   na02f01 U25738 (.o(n21937),
	.a(proc_input_NIB_storage_data_f_12__22_),
	.b(FE_OFN913_n23246));
   oa12f01 U25739 (.o(n7138),
	.a(n21937),
	.b(FE_OFN913_n23246),
	.c(n23820));
   na02f01 U25740 (.o(n21938),
	.a(proc_input_NIB_storage_data_f_12__49_),
	.b(n21911));
   oa12f01 U25741 (.o(n7003),
	.a(n21938),
	.b(n21911),
	.c(n23908));
   na02f01 U25742 (.o(n21939),
	.a(proc_input_NIB_storage_data_f_12__42_),
	.b(n21911));
   oa12f01 U25743 (.o(n7038),
	.a(n21939),
	.b(n21911),
	.c(n23808));
   na02f01 U25744 (.o(n21940),
	.a(proc_input_NIB_storage_data_f_12__50_),
	.b(FE_OFN25628_n21910));
   oa12f01 U25745 (.o(n6998),
	.a(n21940),
	.b(FE_OFN25628_n21910),
	.c(n23903));
   na02f01 U25746 (.o(n21941),
	.a(proc_input_NIB_storage_data_f_12__52_),
	.b(FE_OFN25628_n21910));
   oa12f01 U25747 (.o(n6988),
	.a(n21941),
	.b(FE_OFN25628_n21910),
	.c(n23890));
   in01s01 U25748 (.o(n25970),
	.a(proc_input_NIB_tail_ptr_f_0_));
   na02s01 U25749 (.o(n21942),
	.a(proc_input_NIB_tail_ptr_f_1_),
	.b(n25970));
   na02f01 U25750 (.o(n21946),
	.a(proc_input_NIB_storage_data_f_14__22_),
	.b(FE_OFN25740_FE_OFN25605_n21944));
   oa12f01 U25751 (.o(n7778),
	.a(n21946),
	.b(FE_OFN25740_FE_OFN25605_n21944),
	.c(n23820));
   na02f01 U25752 (.o(n21947),
	.a(proc_input_NIB_storage_data_f_12__41_),
	.b(FE_OFN914_n23246));
   oa12f01 U25753 (.o(n7043),
	.a(n21947),
	.b(FE_OFN914_n23246),
	.c(n23928));
   na02f01 U25754 (.o(n21948),
	.a(proc_input_NIB_storage_data_f_12__24_),
	.b(FE_OFN25626_n21910));
   na02f01 U25755 (.o(n21949),
	.a(proc_input_NIB_storage_data_f_12__40_),
	.b(FE_OFN25627_n21910));
   oa12f01 U25756 (.o(n7048),
	.a(n21949),
	.b(FE_OFN25627_n21910),
	.c(n23800));
   na02f01 U25757 (.o(n21950),
	.a(proc_input_NIB_storage_data_f_12__53_),
	.b(FE_OFN25628_n21910));
   oa12f01 U25758 (.o(n6983),
	.a(n21950),
	.b(FE_OFN25628_n21910),
	.c(n23922));
   na02f01 U25759 (.o(n21951),
	.a(proc_input_NIB_storage_data_f_12__54_),
	.b(FE_OFN25627_n21910));
   na02f01 U25760 (.o(n21952),
	.a(proc_input_NIB_storage_data_f_12__25_),
	.b(FE_OFN913_n23246));
   oa12f01 U25761 (.o(n7123),
	.a(n21952),
	.b(FE_OFN913_n23246),
	.c(n23802));
   na02f01 U25762 (.o(n21953),
	.a(proc_input_NIB_storage_data_f_12__55_),
	.b(FE_OFN25628_n21910));
   oa12f01 U25763 (.o(n6973),
	.a(n21953),
	.b(FE_OFN25628_n21910),
	.c(n23910));
   na02f01 U25764 (.o(n21954),
	.a(proc_input_NIB_storage_data_f_12__63_),
	.b(FE_OFN25628_n21910));
   na02f01 U25765 (.o(n21955),
	.a(proc_input_NIB_storage_data_f_12__62_),
	.b(FE_OFN25628_n21910));
   oa12f01 U25766 (.o(n6938),
	.a(n21955),
	.b(FE_OFN25628_n21910),
	.c(n23810));
   na02f01 U25767 (.o(n21956),
	.a(proc_input_NIB_storage_data_f_12__26_),
	.b(n21911));
   oa12f01 U25768 (.o(n7118),
	.a(n21956),
	.b(n21911),
	.c(n23818));
   na02f01 U25769 (.o(n21957),
	.a(proc_input_NIB_storage_data_f_12__27_),
	.b(FE_OFN913_n23246));
   oa12f01 U25770 (.o(n7113),
	.a(n21957),
	.b(FE_OFN913_n23246),
	.c(n23822));
   na02f01 U25771 (.o(n21958),
	.a(proc_input_NIB_storage_data_f_12__28_),
	.b(FE_OFN913_n23246));
   oa12f01 U25772 (.o(n7108),
	.a(n21958),
	.b(FE_OFN913_n23246),
	.c(n23814));
   oa12f01 U25773 (.o(n7103),
	.a(n21959),
	.b(FE_OFN25626_n21910),
	.c(n23804));
   na02f01 U25774 (.o(n21960),
	.a(proc_input_NIB_storage_data_f_12__30_),
	.b(n21911));
   oa12f01 U25775 (.o(n7098),
	.a(n21960),
	.b(n21911),
	.c(n23894));
   na02f01 U25776 (.o(n21961),
	.a(proc_input_NIB_storage_data_f_12__39_),
	.b(FE_OFN913_n23246));
   na02f01 U25777 (.o(n21962),
	.a(proc_input_NIB_storage_data_f_12__61_),
	.b(FE_OFN25628_n21910));
   na02f01 U25778 (.o(n21963),
	.a(proc_input_NIB_storage_data_f_12__60_),
	.b(FE_OFN25628_n21910));
   oa12f01 U25779 (.o(n6948),
	.a(n21963),
	.b(FE_OFN25628_n21910),
	.c(n23926));
   oa12f01 U25780 (.o(n6953),
	.a(n21964),
	.b(FE_OFN25628_n21910),
	.c(n23938));
   na02f01 U25781 (.o(n21965),
	.a(proc_input_NIB_storage_data_f_12__31_),
	.b(FE_OFN25627_n21910));
   na02f01 U25782 (.o(n21966),
	.a(proc_input_NIB_storage_data_f_12__58_),
	.b(FE_OFN25628_n21910));
   oa12f01 U25783 (.o(n6958),
	.a(n21966),
	.b(FE_OFN25628_n21910),
	.c(n23936));
   na02f01 U25784 (.o(n21967),
	.a(proc_input_NIB_storage_data_f_12__57_),
	.b(FE_OFN25627_n21910));
   oa12f01 U25785 (.o(n6963),
	.a(n21967),
	.b(FE_OFN25627_n21910),
	.c(n23932));
   na02f01 U25786 (.o(n21968),
	.a(proc_input_NIB_storage_data_f_12__56_),
	.b(FE_OFN25628_n21910));
   oa12f01 U25787 (.o(n6968),
	.a(n21968),
	.b(FE_OFN25628_n21910),
	.c(n23930));
   na02f01 U25788 (.o(n21969),
	.a(proc_input_NIB_storage_data_f_12__32_),
	.b(FE_OFN914_n23246));
   oa12f01 U25789 (.o(n7088),
	.a(n21969),
	.b(FE_OFN914_n23246),
	.c(n23905));
   na02f01 U25790 (.o(n21970),
	.a(proc_input_NIB_storage_data_f_12__34_),
	.b(FE_OFN914_n23246));
   oa12f01 U25791 (.o(n7078),
	.a(n21970),
	.b(FE_OFN914_n23246),
	.c(n23816));
   na02f01 U25792 (.o(n21971),
	.a(proc_input_NIB_storage_data_f_12__35_),
	.b(FE_OFN914_n23246));
   oa12f01 U25793 (.o(n7073),
	.a(n21971),
	.b(FE_OFN914_n23246),
	.c(n23944));
   na02f01 U25794 (.o(n21972),
	.a(proc_input_NIB_storage_data_f_12__36_),
	.b(FE_OFN913_n23246));
   oa12f01 U25795 (.o(n7068),
	.a(n21972),
	.b(FE_OFN913_n23246),
	.c(n23940));
   na02f01 U25796 (.o(n21973),
	.a(proc_input_NIB_storage_data_f_12__38_),
	.b(FE_OFN914_n23246));
   oa12f01 U25797 (.o(n7058),
	.a(n21973),
	.b(FE_OFN914_n23246),
	.c(n23812));
   na02f01 U25798 (.o(n21974),
	.a(proc_input_NIB_storage_data_f_13__47_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25799 (.o(n7333),
	.a(n21974),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23914));
   na02f01 U25800 (.o(n21975),
	.a(proc_input_NIB_storage_data_f_12__23_),
	.b(FE_OFN914_n23246));
   oa12f01 U25801 (.o(n7133),
	.a(n21975),
	.b(FE_OFN914_n23246),
	.c(n23793));
   na02f01 U25802 (.o(n21976),
	.a(proc_input_NIB_storage_data_f_13__46_),
	.b(n23236));
   oa12f01 U25803 (.o(n7338),
	.a(n21976),
	.b(n23236),
	.c(n23916));
   na02f01 U25804 (.o(n21977),
	.a(proc_input_NIB_storage_data_f_14__23_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25805 (.o(n7773),
	.a(n21977),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23793));
   na02f01 U25806 (.o(n21979),
	.a(proc_input_NIB_storage_data_f_14__25_),
	.b(FE_OFN25740_FE_OFN25605_n21944));
   oa12f01 U25807 (.o(n7763),
	.a(n21979),
	.b(FE_OFN25740_FE_OFN25605_n21944),
	.c(n23802));
   na02f01 U25808 (.o(n21980),
	.a(proc_input_NIB_storage_data_f_14__26_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25809 (.o(n7758),
	.a(n21980),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23818));
   na02f01 U25810 (.o(n21981),
	.a(proc_input_NIB_storage_data_f_14__27_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25811 (.o(n7753),
	.a(n21981),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23822));
   na02f01 U25812 (.o(n21982),
	.a(proc_input_NIB_storage_data_f_14__28_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25813 (.o(n7748),
	.a(n21982),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23814));
   na02f01 U25814 (.o(n21983),
	.a(proc_input_NIB_storage_data_f_13__27_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25815 (.o(n7433),
	.a(n21983),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23822));
   na02f01 U25816 (.o(n21984),
	.a(proc_input_NIB_storage_data_f_14__29_),
	.b(FE_OFN25739_FE_OFN25605_n21944));
   oa12f01 U25817 (.o(n7743),
	.a(n21984),
	.b(FE_OFN25739_FE_OFN25605_n21944),
	.c(n23804));
   na02f01 U25818 (.o(n21985),
	.a(proc_input_NIB_storage_data_f_14__30_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25819 (.o(n7738),
	.a(n21985),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23894));
   na02f01 U25820 (.o(n21986),
	.a(proc_input_NIB_storage_data_f_14__31_),
	.b(FE_OFN25605_n21944));
   na02f01 U25821 (.o(n21987),
	.a(proc_input_NIB_storage_data_f_14__32_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25822 (.o(n7728),
	.a(n21987),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23905));
   na02f01 U25823 (.o(n21988),
	.a(proc_input_NIB_storage_data_f_14__34_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25824 (.o(n7718),
	.a(n21988),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23816));
   na02f01 U25825 (.o(n21989),
	.a(proc_input_NIB_storage_data_f_14__35_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25826 (.o(n7713),
	.a(n21989),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23944));
   na02f01 U25827 (.o(n21990),
	.a(proc_input_NIB_storage_data_f_14__36_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25828 (.o(n7708),
	.a(n21990),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23940));
   na02f01 U25829 (.o(n21991),
	.a(proc_input_NIB_storage_data_f_14__37_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25830 (.o(n7703),
	.a(n21991),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23796));
   na02f01 U25831 (.o(n21992),
	.a(proc_input_NIB_storage_data_f_14__38_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25832 (.o(n7698),
	.a(n21992),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23812));
   na02f01 U25833 (.o(n21994),
	.a(proc_input_NIB_storage_data_f_14__40_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25834 (.o(n7688),
	.a(n21994),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23800));
   na02f01 U25835 (.o(n21995),
	.a(proc_input_NIB_storage_data_f_14__41_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25836 (.o(n7683),
	.a(n21995),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23928));
   na02f01 U25837 (.o(n21996),
	.a(proc_input_NIB_storage_data_f_14__42_),
	.b(FE_OFN453_n23262));
   oa12f01 U25838 (.o(n7678),
	.a(n21996),
	.b(FE_OFN453_n23262),
	.c(n23808));
   na02f01 U25839 (.o(n21997),
	.a(proc_input_NIB_storage_data_f_14__43_),
	.b(FE_OFN25740_FE_OFN25605_n21944));
   oa12f01 U25840 (.o(n7673),
	.a(n21997),
	.b(FE_OFN25740_FE_OFN25605_n21944),
	.c(n23806));
   na02f01 U25841 (.o(n21999),
	.a(proc_input_NIB_storage_data_f_14__44_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25842 (.o(n7668),
	.a(n21999),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23920));
   na02f01 U25843 (.o(n22000),
	.a(proc_input_NIB_storage_data_f_14__45_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25844 (.o(n7663),
	.a(n22000),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23942));
   na02f01 U25845 (.o(n22001),
	.a(proc_input_NIB_storage_data_f_14__46_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25846 (.o(n7658),
	.a(n22001),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23916));
   na02f01 U25847 (.o(n22002),
	.a(proc_input_NIB_storage_data_f_13__24_),
	.b(n23236));
   na02f01 U25848 (.o(n22003),
	.a(proc_input_NIB_storage_data_f_13__45_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25849 (.o(n7343),
	.a(n22003),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23942));
   na02f01 U25850 (.o(n22004),
	.a(proc_input_NIB_storage_data_f_13__26_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25851 (.o(n7438),
	.a(n22004),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23818));
   na02f01 U25852 (.o(n22005),
	.a(proc_input_NIB_storage_data_f_14__58_),
	.b(FE_OFN453_n23262));
   oa12f01 U25853 (.o(n7598),
	.a(n22005),
	.b(FE_OFN453_n23262),
	.c(n23936));
   na02f01 U25854 (.o(n22006),
	.a(proc_input_NIB_storage_data_f_14__47_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25855 (.o(n7653),
	.a(n22006),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23914));
   na02f01 U25856 (.o(n22007),
	.a(proc_input_NIB_storage_data_f_14__48_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25857 (.o(n7648),
	.a(n22007),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23912));
   na02f01 U25858 (.o(n22008),
	.a(proc_input_NIB_storage_data_f_14__49_),
	.b(FE_OFN25742_FE_OFN25605_n21944));
   oa12f01 U25859 (.o(n7643),
	.a(n22008),
	.b(FE_OFN25742_FE_OFN25605_n21944),
	.c(n23908));
   na02f01 U25860 (.o(n22009),
	.a(proc_input_NIB_storage_data_f_14__50_),
	.b(FE_OFN25741_FE_OFN25605_n21944));
   oa12f01 U25861 (.o(n7638),
	.a(n22009),
	.b(FE_OFN25741_FE_OFN25605_n21944),
	.c(n23903));
   na02f01 U25862 (.o(n22010),
	.a(proc_input_NIB_storage_data_f_13__40_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25863 (.o(n7368),
	.a(n22010),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23800));
   na02f01 U25864 (.o(n22011),
	.a(proc_input_NIB_storage_data_f_13__39_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   na02f01 U25865 (.o(n22012),
	.a(proc_input_NIB_storage_data_f_13__38_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25866 (.o(n7378),
	.a(n22012),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23812));
   na02f01 U25867 (.o(n22013),
	.a(proc_input_NIB_storage_data_f_14__60_),
	.b(FE_OFN453_n23262));
   oa12f01 U25868 (.o(n7588),
	.a(n22013),
	.b(FE_OFN453_n23262),
	.c(n23926));
   na02f01 U25869 (.o(n22014),
	.a(proc_input_NIB_storage_data_f_14__52_),
	.b(FE_OFN25741_FE_OFN25605_n21944));
   oa12f01 U25870 (.o(n7628),
	.a(n22014),
	.b(FE_OFN25741_FE_OFN25605_n21944),
	.c(n23890));
   na02f01 U25871 (.o(n22015),
	.a(proc_input_NIB_storage_data_f_14__53_),
	.b(FE_OFN25741_FE_OFN25605_n21944));
   oa12f01 U25872 (.o(n7623),
	.a(n22015),
	.b(FE_OFN25741_FE_OFN25605_n21944),
	.c(n23922));
   oa12f01 U25873 (.o(n7398),
	.a(n22016),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23816));
   na02f01 U25874 (.o(n22017),
	.a(proc_input_NIB_storage_data_f_14__55_),
	.b(FE_OFN25741_FE_OFN25605_n21944));
   oa12f01 U25875 (.o(n7613),
	.a(n22017),
	.b(FE_OFN25741_FE_OFN25605_n21944),
	.c(n23910));
   na02f01 U25876 (.o(n22018),
	.a(proc_input_NIB_storage_data_f_14__56_),
	.b(FE_OFN25741_FE_OFN25605_n21944));
   oa12f01 U25877 (.o(n7608),
	.a(n22018),
	.b(FE_OFN25741_FE_OFN25605_n21944),
	.c(n23930));
   na02f01 U25878 (.o(n22019),
	.a(proc_input_NIB_storage_data_f_14__57_),
	.b(FE_OFN25605_n21944));
   oa12f01 U25879 (.o(n7603),
	.a(n22019),
	.b(FE_OFN25605_n21944),
	.c(n23932));
   na02f01 U25880 (.o(n22020),
	.a(proc_input_NIB_storage_data_f_14__62_),
	.b(FE_OFN453_n23262));
   oa12f01 U25881 (.o(n7578),
	.a(n22020),
	.b(FE_OFN453_n23262),
	.c(n23810));
   na02f01 U25882 (.o(n22021),
	.a(proc_input_NIB_storage_data_f_14__63_),
	.b(FE_OFN25741_FE_OFN25605_n21944));
   na02f01 U25883 (.o(n22022),
	.a(proc_input_NIB_storage_data_f_13__29_),
	.b(n23236));
   oa12f01 U25884 (.o(n7423),
	.a(n22022),
	.b(n23236),
	.c(n23804));
   na02f01 U25885 (.o(n22023),
	.a(proc_input_NIB_storage_data_f_13__23_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25886 (.o(n7453),
	.a(n22023),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23793));
   na02f01 U25887 (.o(n22024),
	.a(proc_input_NIB_storage_data_f_13__44_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25888 (.o(n7348),
	.a(n22024),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23920));
   na02f01 U25889 (.o(n22025),
	.a(proc_input_NIB_storage_data_f_13__43_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25890 (.o(n7353),
	.a(n22025),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23806));
   na02f01 U25891 (.o(n22026),
	.a(proc_input_NIB_storage_data_f_13__42_),
	.b(n23236));
   oa12f01 U25892 (.o(n7358),
	.a(n22026),
	.b(n23236),
	.c(n23808));
   na02f01 U25893 (.o(n22027),
	.a(proc_input_NIB_storage_data_f_13__41_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25894 (.o(n7363),
	.a(n22027),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23928));
   na02f01 U25895 (.o(n22028),
	.a(proc_input_NIB_storage_data_f_13__28_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25896 (.o(n7428),
	.a(n22028),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23814));
   na02f01 U25897 (.o(n22029),
	.a(proc_input_NIB_storage_data_f_13__30_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25898 (.o(n7418),
	.a(n22029),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23894));
   na02f01 U25899 (.o(n22030),
	.a(proc_input_NIB_storage_data_f_14__59_),
	.b(FE_OFN453_n23262));
   oa12f01 U25900 (.o(n7593),
	.a(n22030),
	.b(FE_OFN453_n23262),
	.c(n23938));
   na02f01 U25901 (.o(n22031),
	.a(proc_input_NIB_storage_data_f_13__37_),
	.b(n23236));
   oa12f01 U25902 (.o(n7383),
	.a(n22031),
	.b(n23236),
	.c(n23796));
   na02f01 U25903 (.o(n22032),
	.a(proc_input_NIB_storage_data_f_13__36_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25904 (.o(n7388),
	.a(n22032),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23940));
   na02f01 U25905 (.o(n22033),
	.a(proc_input_NIB_storage_data_f_13__35_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   na02f01 U25906 (.o(n22034),
	.a(proc_input_NIB_storage_data_f_13__22_),
	.b(FE_OFN448_n23236));
   oa12f01 U25907 (.o(n7458),
	.a(n22034),
	.b(FE_OFN448_n23236),
	.c(n23820));
   na02f01 U25908 (.o(n22035),
	.a(proc_input_NIB_storage_data_f_13__32_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25909 (.o(n7408),
	.a(n22035),
	.b(FE_OFN25782_FE_OFN448_n23236),
	.c(n23905));
   na02f01 U25910 (.o(n22036),
	.a(proc_input_NIB_storage_data_f_13__31_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   na02f01 U25911 (.o(n22037),
	.a(proc_input_NIB_storage_data_f_13__25_),
	.b(FE_OFN25782_FE_OFN448_n23236));
   oa12f01 U25912 (.o(n7443),
	.a(n22037),
	.b(FE_OFN448_n23236),
	.c(n23802));
   na02f01 U25913 (.o(n22038),
	.a(proc_input_NIB_storage_data_f_14__61_),
	.b(FE_OFN453_n23262));
   oa12f01 U25914 (.o(n7583),
	.a(n22038),
	.b(FE_OFN453_n23262),
	.c(n23918));
   na02f01 U25915 (.o(n22039),
	.a(proc_input_NIB_storage_data_f_12__51_),
	.b(FE_OFN25628_n21910));
   oa12f01 U25916 (.o(n6993),
	.a(n22039),
	.b(FE_OFN25628_n21910),
	.c(n23947));
   na02f01 U25917 (.o(n22040),
	.a(proc_input_NIB_storage_data_f_13__51_),
	.b(FE_OFN25781_FE_OFN448_n23236));
   oa12f01 U25918 (.o(n7313),
	.a(n22040),
	.b(FE_OFN25781_FE_OFN448_n23236),
	.c(n23947));
   na02f01 U25919 (.o(n22041),
	.a(proc_input_NIB_storage_data_f_14__51_),
	.b(FE_OFN453_n23262));
   oa12f01 U25920 (.o(n7633),
	.a(n22041),
	.b(FE_OFN453_n23262),
	.c(n23947));
   in01s01 U25921 (.o(n13043),
	.a(n22042));
   oa22f01 U25922 (.o(n22043),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_9_),
	.c(north_input_NIB_storage_data_f_2__9_),
	.d(n20656));
   in01s01 U25923 (.o(n13013),
	.a(n22043));
   in01s01 U25924 (.o(n13048),
	.a(n22044));
   in01s01 U25925 (.o(n13058),
	.a(n22045));
   in01s01 U25926 (.o(n12988),
	.a(n22046));
   in01s01 U25927 (.o(n12983),
	.a(n22047));
   oa22f01 U25928 (.o(n22048),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_10_),
	.c(north_input_NIB_storage_data_f_2__10_),
	.d(n20656));
   in01s01 U25929 (.o(n13008),
	.a(n22048));
   oa22f01 U25930 (.o(n22049),
	.a(FE_OFN25875_n25842),
	.b(dataIn_N_17_),
	.c(north_input_NIB_storage_data_f_2__17_),
	.d(n20656));
   in01s01 U25931 (.o(n12973),
	.a(n22049));
   in01s01 U25932 (.o(n13038),
	.a(n22050));
   oa22f01 U25933 (.o(n22051),
	.a(FE_OFN25875_n25842),
	.b(dataIn_N_20_),
	.c(north_input_NIB_storage_data_f_2__20_),
	.d(n20656));
   in01s01 U25934 (.o(n12958),
	.a(n22051));
   oa22f01 U25935 (.o(n22052),
	.a(FE_OFN25875_n25842),
	.b(dataIn_N_12_),
	.c(north_input_NIB_storage_data_f_2__12_),
	.d(n20656));
   in01s01 U25936 (.o(n12998),
	.a(n22052));
   oa22f01 U25937 (.o(n22053),
	.a(n25842),
	.b(dataIn_N_33_),
	.c(north_input_NIB_storage_data_f_2__33_),
	.d(n20656));
   in01s01 U25938 (.o(n12893),
	.a(n22053));
   in01s01 U25939 (.o(n13033),
	.a(n22054));
   in01s01 U25940 (.o(n13053),
	.a(n22055));
   oa22f01 U25941 (.o(n22056),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_16_),
	.c(north_input_NIB_storage_data_f_2__16_),
	.d(n20656));
   in01s01 U25942 (.o(n12978),
	.a(n22056));
   oa22f01 U25943 (.o(n22057),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_7_),
	.c(north_input_NIB_storage_data_f_2__7_),
	.d(n20656));
   in01s01 U25944 (.o(n13023),
	.a(n22057));
   oa22f01 U25945 (.o(n22058),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_8_),
	.c(north_input_NIB_storage_data_f_2__8_),
	.d(n20656));
   oa22f01 U25946 (.o(n22059),
	.a(FE_OFN25876_n25842),
	.b(dataIn_N_11_),
	.c(north_input_NIB_storage_data_f_2__11_),
	.d(n20656));
   in01s01 U25947 (.o(n13003),
	.a(n22059));
   in01s01 U25948 (.o(n22067),
	.a(proc_output_space_count_f_1_));
   in01s01 U25949 (.o(n22079),
	.a(proc_output_space_count_f_0_));
   no02m01 U25950 (.o(n22062),
	.a(proc_output_space_count_f_1_),
	.b(n22069));
   no02m01 U25951 (.o(n22063),
	.a(n22071),
	.b(n22062));
   in01s01 U25952 (.o(n22065),
	.a(proc_output_space_count_f_2_));
   oa22f01 U25953 (.o(n22064),
	.a(proc_output_space_count_f_2_),
	.b(n22071),
	.c(n22063),
	.d(n22065));
   na02f01 U25954 (.o(proc_output_space_N44),
	.a(FE_OFN25598_reset),
	.b(n22064));
   no02s01 U25955 (.o(n22076),
	.a(proc_output_space_count_f_1_),
	.b(n22065));
   na02s01 U25956 (.o(n22068),
	.a(n22067),
	.b(n22082));
   na02s01 U25957 (.o(n22070),
	.a(n22069),
	.b(n22068));
   na02f01 U25958 (.o(proc_output_space_N48),
	.a(n22074),
	.b(n25825));
   no02s01 U25959 (.o(n22075),
	.a(proc_output_space_count_f_1_),
	.b(proc_output_space_count_f_2_));
   in01s01 U25960 (.o(n22078),
	.a(n22075));
   no02s01 U25961 (.o(n22077),
	.a(proc_output_space_valid_f),
	.b(n22076));
   ao22s01 U25962 (.o(n22080),
	.a(n22941),
	.b(n22078),
	.c(proc_output_space_yummy_f),
	.d(n22077));
   na02s01 U25963 (.o(n25824),
	.a(n22082),
	.b(n22081));
   ao12m02 U25964 (.o(east_input_control_N51),
	.a(east_input_control_N41),
	.b(FE_OFN575_n25463),
	.c(n22083));
   na02f01 U25965 (.o(n22086),
	.a(proc_input_NIB_storage_data_f_8__60_),
	.b(n23471));
   na02f01 U25966 (.o(n22087),
	.a(proc_input_NIB_storage_data_f_8__59_),
	.b(n23471));
   oa12f01 U25967 (.o(n5673),
	.a(n22087),
	.b(n23471),
	.c(n23938));
   na02f01 U25968 (.o(n22088),
	.a(proc_input_NIB_storage_data_f_8__58_),
	.b(n23471));
   oa12f01 U25969 (.o(n5678),
	.a(n22088),
	.b(n23471),
	.c(n23936));
   na02f01 U25970 (.o(n22089),
	.a(proc_input_NIB_storage_data_f_8__57_),
	.b(n23471));
   oa12f01 U25971 (.o(n5683),
	.a(n22089),
	.b(n23471),
	.c(n23932));
   na02f01 U25972 (.o(n22090),
	.a(proc_input_NIB_storage_data_f_8__61_),
	.b(n23471));
   oa12f01 U25973 (.o(n5663),
	.a(n22090),
	.b(n23471),
	.c(n23918));
   na02f01 U25974 (.o(n22091),
	.a(proc_input_NIB_storage_data_f_8__55_),
	.b(n23471));
   oa12f01 U25975 (.o(n5693),
	.a(n22091),
	.b(n23471),
	.c(n23910));
   na02f01 U25976 (.o(n22092),
	.a(proc_input_NIB_storage_data_f_8__54_),
	.b(n23471));
   na02f01 U25977 (.o(n22093),
	.a(proc_input_NIB_storage_data_f_8__53_),
	.b(n23471));
   oa12f01 U25978 (.o(n5703),
	.a(n22093),
	.b(n23471),
	.c(n23922));
   oa12f01 U25979 (.o(n5708),
	.a(n22094),
	.b(n23471),
	.c(n23890));
   na02f01 U25980 (.o(n22095),
	.a(proc_input_NIB_storage_data_f_8__56_),
	.b(n23471));
   oa12f01 U25981 (.o(n5688),
	.a(n22095),
	.b(n23471),
	.c(n23930));
   no02f01 U25982 (.o(n22096),
	.a(proc_input_NIB_tail_ptr_f_1_),
	.b(n25970));
   na02f01 U25983 (.o(n22099),
	.a(proc_input_NIB_storage_data_f_9__38_),
	.b(FE_OFN101_n22098));
   oa12f01 U25984 (.o(n6098),
	.a(n22099),
	.b(FE_OFN101_n22098),
	.c(n23812));
   na02f01 U25985 (.o(n22100),
	.a(proc_input_NIB_storage_data_f_8__48_),
	.b(n22085));
   oa12f01 U25986 (.o(n5728),
	.a(n22100),
	.b(n22085),
	.c(n23912));
   na02f01 U25987 (.o(n22101),
	.a(proc_input_NIB_storage_data_f_8__47_),
	.b(n22085));
   oa12f01 U25988 (.o(n5733),
	.a(n22101),
	.b(n22085),
	.c(n23914));
   na02f01 U25989 (.o(n22102),
	.a(proc_input_NIB_storage_data_f_8__46_),
	.b(n22085));
   oa12f01 U25990 (.o(n5738),
	.a(n22102),
	.b(n22085),
	.c(n23916));
   na02f01 U25991 (.o(n22103),
	.a(proc_input_NIB_storage_data_f_8__45_),
	.b(n22085));
   na02f01 U25992 (.o(n22104),
	.a(proc_input_NIB_storage_data_f_8__44_),
	.b(n22085));
   oa12f01 U25993 (.o(n5748),
	.a(n22104),
	.b(n22085),
	.c(n23920));
   na02f01 U25994 (.o(n22105),
	.a(proc_input_NIB_storage_data_f_8__43_),
	.b(n22085));
   oa12f01 U25995 (.o(n5753),
	.a(n22105),
	.b(n22085),
	.c(n23806));
   na02f01 U25996 (.o(n22106),
	.a(proc_input_NIB_storage_data_f_8__42_),
	.b(n22085));
   oa12f01 U25997 (.o(n5758),
	.a(n22106),
	.b(n22085),
	.c(n23808));
   na02f01 U25998 (.o(n22107),
	.a(proc_input_NIB_storage_data_f_8__41_),
	.b(n22085));
   oa12f01 U25999 (.o(n5763),
	.a(n22107),
	.b(n22085),
	.c(n23928));
   na02f01 U26000 (.o(n22108),
	.a(proc_input_NIB_storage_data_f_8__40_),
	.b(n23471));
   oa12f01 U26001 (.o(n5768),
	.a(n22108),
	.b(n23471),
	.c(n23800));
   na02f01 U26002 (.o(n22109),
	.a(proc_input_NIB_storage_data_f_8__39_),
	.b(n22085));
   na02f01 U26003 (.o(n22110),
	.a(proc_input_NIB_storage_data_f_8__38_),
	.b(n22085));
   oa12f01 U26004 (.o(n5778),
	.a(n22110),
	.b(n22085),
	.c(n23812));
   na02f01 U26005 (.o(n22111),
	.a(proc_input_NIB_storage_data_f_8__50_),
	.b(n23471));
   oa12f01 U26006 (.o(n5718),
	.a(n22111),
	.b(n23471),
	.c(n23903));
   na02f01 U26007 (.o(n22112),
	.a(proc_input_NIB_storage_data_f_8__49_),
	.b(n22085));
   oa12f01 U26008 (.o(n5723),
	.a(n22112),
	.b(n22085),
	.c(n23908));
   oa12f01 U26009 (.o(n5783),
	.a(n22113),
	.b(n22085),
	.c(n23796));
   na02f01 U26010 (.o(n22114),
	.a(proc_input_NIB_storage_data_f_8__36_),
	.b(n22085));
   oa12f01 U26011 (.o(n5788),
	.a(n22114),
	.b(n22085),
	.c(n23940));
   na02f01 U26012 (.o(n22115),
	.a(proc_input_NIB_storage_data_f_8__35_),
	.b(n22085));
   oa12f01 U26013 (.o(n5793),
	.a(n22115),
	.b(n22085),
	.c(n23944));
   na02f01 U26014 (.o(n22116),
	.a(proc_input_NIB_storage_data_f_8__34_),
	.b(n22085));
   oa12f01 U26015 (.o(n5798),
	.a(n22116),
	.b(n22085),
	.c(n23816));
   na02f01 U26016 (.o(n22117),
	.a(proc_input_NIB_storage_data_f_8__62_),
	.b(n23471));
   oa12f01 U26017 (.o(n5658),
	.a(n22117),
	.b(n23471),
	.c(n23810));
   na02f01 U26018 (.o(n22118),
	.a(proc_input_NIB_storage_data_f_8__32_),
	.b(n22085));
   oa12f01 U26019 (.o(n5808),
	.a(n22118),
	.b(n22085),
	.c(n23905));
   na02f01 U26020 (.o(n22119),
	.a(proc_input_NIB_storage_data_f_8__31_),
	.b(n23471));
   na02f01 U26021 (.o(n22120),
	.a(proc_input_NIB_storage_data_f_8__30_),
	.b(n22085));
   na02f01 U26022 (.o(n22121),
	.a(proc_input_NIB_storage_data_f_8__29_),
	.b(n22085));
   oa12f01 U26023 (.o(n5823),
	.a(n22121),
	.b(n22085),
	.c(n23804));
   na02f01 U26024 (.o(n22122),
	.a(proc_input_NIB_storage_data_f_8__28_),
	.b(n22085));
   oa12f01 U26025 (.o(n5828),
	.a(n22122),
	.b(n22085),
	.c(n23814));
   na02f01 U26026 (.o(n22123),
	.a(proc_input_NIB_storage_data_f_8__27_),
	.b(n22085));
   oa12f01 U26027 (.o(n5833),
	.a(n22123),
	.b(n22085),
	.c(n23822));
   na02f01 U26028 (.o(n22124),
	.a(proc_input_NIB_storage_data_f_8__26_),
	.b(n22085));
   oa12f01 U26029 (.o(n5838),
	.a(n22124),
	.b(n22085),
	.c(n23818));
   na02f01 U26030 (.o(n22125),
	.a(proc_input_NIB_storage_data_f_8__25_),
	.b(n22085));
   oa12f01 U26031 (.o(n5843),
	.a(n22125),
	.b(n22085),
	.c(n23802));
   na02f01 U26032 (.o(n22126),
	.a(proc_input_NIB_storage_data_f_8__24_),
	.b(n22085));
   na02f01 U26033 (.o(n22127),
	.a(proc_input_NIB_storage_data_f_8__23_),
	.b(n22085));
   oa12f01 U26034 (.o(n5853),
	.a(n22127),
	.b(n22085),
	.c(n23793));
   oa12f01 U26035 (.o(n5858),
	.a(n22128),
	.b(n22085),
	.c(n23820));
   na02f01 U26036 (.o(n22129),
	.a(proc_input_NIB_storage_data_f_9__63_),
	.b(FE_OFN465_n23476));
   na02f01 U26037 (.o(n22130),
	.a(proc_input_NIB_storage_data_f_9__62_),
	.b(FE_OFN465_n23476));
   oa12f01 U26038 (.o(n5978),
	.a(n22130),
	.b(FE_OFN465_n23476),
	.c(n23810));
   na02f01 U26039 (.o(n22131),
	.a(proc_input_NIB_storage_data_f_9__61_),
	.b(FE_OFN465_n23476));
   oa12f01 U26040 (.o(n5983),
	.a(n22131),
	.b(FE_OFN465_n23476),
	.c(n23918));
   na02f01 U26041 (.o(n22132),
	.a(proc_input_NIB_storage_data_f_9__60_),
	.b(FE_OFN465_n23476));
   oa12f01 U26042 (.o(n5988),
	.a(n22132),
	.b(FE_OFN465_n23476),
	.c(n23926));
   na02f01 U26043 (.o(n22133),
	.a(proc_input_NIB_storage_data_f_9__59_),
	.b(FE_OFN465_n23476));
   oa12f01 U26044 (.o(n5993),
	.a(n22133),
	.b(FE_OFN465_n23476),
	.c(n23938));
   na02f01 U26045 (.o(n22134),
	.a(proc_input_NIB_storage_data_f_9__58_),
	.b(FE_OFN465_n23476));
   oa12f01 U26046 (.o(n5998),
	.a(n22134),
	.b(FE_OFN465_n23476),
	.c(n23936));
   oa12f01 U26047 (.o(n6003),
	.a(n22135),
	.b(FE_OFN465_n23476),
	.c(n23932));
   na02f01 U26048 (.o(n22136),
	.a(proc_input_NIB_storage_data_f_9__56_),
	.b(FE_OFN465_n23476));
   oa12f01 U26049 (.o(n6008),
	.a(n22136),
	.b(FE_OFN465_n23476),
	.c(n23930));
   no02f01 U26050 (.o(n22138),
	.a(proc_input_NIB_tail_ptr_f_0_),
	.b(n22137));
   na02f01 U26051 (.o(n22141),
	.a(proc_input_NIB_storage_data_f_10__22_),
	.b(FE_OFN103_n22140));
   oa12f01 U26052 (.o(n6498),
	.a(n22141),
	.b(FE_OFN103_n22140),
	.c(n23820));
   na02f01 U26053 (.o(n22142),
	.a(proc_input_NIB_storage_data_f_10__23_),
	.b(FE_OFN103_n22140));
   na02f01 U26054 (.o(n22143),
	.a(proc_input_NIB_storage_data_f_10__24_),
	.b(n23453));
   na02f01 U26055 (.o(n22144),
	.a(proc_input_NIB_storage_data_f_10__25_),
	.b(FE_OFN103_n22140));
   oa12f01 U26056 (.o(n6483),
	.a(n22144),
	.b(FE_OFN103_n22140),
	.c(n23802));
   na02f01 U26057 (.o(n22145),
	.a(proc_input_NIB_storage_data_f_10__26_),
	.b(n23453));
   oa12f01 U26058 (.o(n6478),
	.a(n22145),
	.b(n23453),
	.c(n23818));
   na02f01 U26059 (.o(n22146),
	.a(proc_input_NIB_storage_data_f_10__27_),
	.b(FE_OFN103_n22140));
   oa12f01 U26060 (.o(n6473),
	.a(n22146),
	.b(FE_OFN103_n22140),
	.c(n23822));
   na02f01 U26061 (.o(n22147),
	.a(proc_input_NIB_storage_data_f_10__28_),
	.b(FE_OFN103_n22140));
   oa12f01 U26062 (.o(n6468),
	.a(n22147),
	.b(FE_OFN103_n22140),
	.c(n23814));
   na02f01 U26063 (.o(n22148),
	.a(proc_input_NIB_storage_data_f_10__29_),
	.b(n23453));
   oa12f01 U26064 (.o(n6463),
	.a(n22148),
	.b(n23453),
	.c(n23804));
   na02f01 U26065 (.o(n22149),
	.a(proc_input_NIB_storage_data_f_10__30_),
	.b(n23453));
   oa12f01 U26066 (.o(n6458),
	.a(n22149),
	.b(n23453),
	.c(n23894));
   na02f01 U26067 (.o(n22150),
	.a(proc_input_NIB_storage_data_f_10__31_),
	.b(FE_OFN103_n22140));
   oa12f01 U26068 (.o(n6448),
	.a(n22151),
	.b(FE_OFN103_n22140),
	.c(n23905));
   na02f01 U26069 (.o(n22152),
	.a(proc_input_NIB_storage_data_f_9__55_),
	.b(FE_OFN465_n23476));
   oa12f01 U26070 (.o(n6013),
	.a(n22152),
	.b(FE_OFN465_n23476),
	.c(n23910));
   na02f01 U26071 (.o(n22153),
	.a(proc_input_NIB_storage_data_f_10__34_),
	.b(FE_OFN103_n22140));
   oa12f01 U26072 (.o(n6438),
	.a(n22153),
	.b(FE_OFN103_n22140),
	.c(n23816));
   na02f01 U26073 (.o(n22154),
	.a(proc_input_NIB_storage_data_f_10__35_),
	.b(FE_OFN103_n22140));
   oa12f01 U26074 (.o(n6433),
	.a(n22154),
	.b(FE_OFN103_n22140),
	.c(n23944));
   na02f01 U26075 (.o(n22155),
	.a(proc_input_NIB_storage_data_f_10__36_),
	.b(FE_OFN103_n22140));
   oa12f01 U26076 (.o(n6428),
	.a(n22155),
	.b(FE_OFN103_n22140),
	.c(n23940));
   na02f01 U26077 (.o(n22156),
	.a(proc_input_NIB_storage_data_f_8__63_),
	.b(n23471));
   na02f01 U26078 (.o(n22157),
	.a(proc_input_NIB_storage_data_f_10__37_),
	.b(FE_OFN103_n22140));
   oa12f01 U26079 (.o(n6423),
	.a(n22157),
	.b(FE_OFN103_n22140),
	.c(n23796));
   na02f01 U26080 (.o(n22158),
	.a(proc_input_NIB_storage_data_f_10__38_),
	.b(FE_OFN103_n22140));
   na02f01 U26081 (.o(n22159),
	.a(proc_input_NIB_storage_data_f_10__39_),
	.b(FE_OFN103_n22140));
   na02f01 U26082 (.o(n22160),
	.a(proc_input_NIB_storage_data_f_10__40_),
	.b(FE_OFN103_n22140));
   oa12f01 U26083 (.o(n6408),
	.a(n22160),
	.b(FE_OFN103_n22140),
	.c(n23800));
   na02f01 U26084 (.o(n22161),
	.a(proc_input_NIB_storage_data_f_10__41_),
	.b(FE_OFN103_n22140));
   oa12f01 U26085 (.o(n6403),
	.a(n22161),
	.b(FE_OFN103_n22140),
	.c(n23928));
   na02f01 U26086 (.o(n22162),
	.a(proc_input_NIB_storage_data_f_10__42_),
	.b(n23453));
   oa12f01 U26087 (.o(n6398),
	.a(n22162),
	.b(n23453),
	.c(n23808));
   na02f01 U26088 (.o(n22163),
	.a(proc_input_NIB_storage_data_f_10__43_),
	.b(FE_OFN103_n22140));
   oa12f01 U26089 (.o(n6393),
	.a(n22163),
	.b(FE_OFN103_n22140),
	.c(n23806));
   na02f01 U26090 (.o(n22164),
	.a(proc_input_NIB_storage_data_f_10__44_),
	.b(FE_OFN103_n22140));
   oa12f01 U26091 (.o(n6388),
	.a(n22164),
	.b(FE_OFN103_n22140),
	.c(n23920));
   na02f01 U26092 (.o(n22165),
	.a(proc_input_NIB_storage_data_f_10__45_),
	.b(FE_OFN103_n22140));
   oa12f01 U26093 (.o(n6383),
	.a(n22165),
	.b(FE_OFN103_n22140),
	.c(n23942));
   na02f01 U26094 (.o(n22166),
	.a(proc_input_NIB_storage_data_f_10__46_),
	.b(n23453));
   oa12f01 U26095 (.o(n6378),
	.a(n22166),
	.b(n23453),
	.c(n23916));
   oa12f01 U26096 (.o(n6373),
	.a(n22167),
	.b(FE_OFN103_n22140),
	.c(n23914));
   na02f01 U26097 (.o(n22168),
	.a(proc_input_NIB_storage_data_f_10__48_),
	.b(n23453));
   oa12f01 U26098 (.o(n6368),
	.a(n22168),
	.b(n23453),
	.c(n23912));
   na02f01 U26099 (.o(n22169),
	.a(proc_input_NIB_storage_data_f_10__49_),
	.b(n23453));
   oa12f01 U26100 (.o(n6363),
	.a(n22169),
	.b(n23453),
	.c(n23908));
   na02f01 U26101 (.o(n22170),
	.a(proc_input_NIB_storage_data_f_10__50_),
	.b(n23453));
   oa12f01 U26102 (.o(n6358),
	.a(n22170),
	.b(n23453),
	.c(n23903));
   na02f01 U26103 (.o(n22171),
	.a(proc_input_NIB_storage_data_f_10__51_),
	.b(n23453));
   oa12f01 U26104 (.o(n6353),
	.a(n22171),
	.b(n23453),
	.c(n23947));
   na02f01 U26105 (.o(n22172),
	.a(proc_input_NIB_storage_data_f_10__52_),
	.b(n23453));
   oa12f01 U26106 (.o(n6348),
	.a(n22172),
	.b(n23453),
	.c(n23890));
   na02f01 U26107 (.o(n22173),
	.a(proc_input_NIB_storage_data_f_10__53_),
	.b(FE_OFN103_n22140));
   na02f01 U26108 (.o(n22174),
	.a(proc_input_NIB_storage_data_f_10__54_),
	.b(FE_OFN103_n22140));
   na02f01 U26109 (.o(n22175),
	.a(proc_input_NIB_storage_data_f_10__55_),
	.b(FE_OFN103_n22140));
   oa12f01 U26110 (.o(n6333),
	.a(n22175),
	.b(FE_OFN103_n22140),
	.c(n23910));
   na02f01 U26111 (.o(n22176),
	.a(proc_input_NIB_storage_data_f_10__56_),
	.b(FE_OFN103_n22140));
   oa12f01 U26112 (.o(n6328),
	.a(n22176),
	.b(FE_OFN103_n22140),
	.c(n23930));
   na02f01 U26113 (.o(n22177),
	.a(proc_input_NIB_storage_data_f_10__57_),
	.b(FE_OFN103_n22140));
   oa12f01 U26114 (.o(n6323),
	.a(n22177),
	.b(FE_OFN103_n22140),
	.c(n23932));
   na02f01 U26115 (.o(n22178),
	.a(proc_input_NIB_storage_data_f_10__58_),
	.b(n23453));
   oa12f01 U26116 (.o(n6318),
	.a(n22178),
	.b(n23453),
	.c(n23936));
   na02f01 U26117 (.o(n22179),
	.a(proc_input_NIB_storage_data_f_9__23_),
	.b(FE_OFN101_n22098));
   oa12f01 U26118 (.o(n6173),
	.a(n22179),
	.b(FE_OFN101_n22098),
	.c(n23793));
   na02f01 U26119 (.o(n22180),
	.a(proc_input_NIB_storage_data_f_9__24_),
	.b(FE_OFN101_n22098));
   na02f01 U26120 (.o(n22181),
	.a(proc_input_NIB_storage_data_f_10__59_),
	.b(n23453));
   oa12f01 U26121 (.o(n6313),
	.a(n22181),
	.b(n23453),
	.c(n23938));
   na02f01 U26122 (.o(n22182),
	.a(proc_input_NIB_storage_data_f_10__60_),
	.b(n23453));
   oa12f01 U26123 (.o(n6308),
	.a(n22182),
	.b(n23453),
	.c(n23926));
   na02f01 U26124 (.o(n22183),
	.a(proc_input_NIB_storage_data_f_10__61_),
	.b(n23453));
   oa12f01 U26125 (.o(n6303),
	.a(n22183),
	.b(n23453),
	.c(n23918));
   oa12f01 U26126 (.o(n6298),
	.a(n22184),
	.b(n23453),
	.c(n23810));
   na02f01 U26127 (.o(n22185),
	.a(proc_input_NIB_storage_data_f_10__63_),
	.b(FE_OFN103_n22140));
   na02f01 U26128 (.o(n22186),
	.a(proc_input_NIB_storage_data_f_9__54_),
	.b(FE_OFN465_n23476));
   na02f01 U26129 (.o(n22187),
	.a(proc_input_NIB_storage_data_f_9__53_),
	.b(FE_OFN465_n23476));
   oa12f01 U26130 (.o(n6023),
	.a(n22187),
	.b(FE_OFN465_n23476),
	.c(n23922));
   na02f01 U26131 (.o(n22188),
	.a(proc_input_NIB_storage_data_f_9__52_),
	.b(FE_OFN465_n23476));
   oa12f01 U26132 (.o(n6028),
	.a(n22188),
	.b(FE_OFN465_n23476),
	.c(n23890));
   na02f01 U26133 (.o(n22189),
	.a(proc_input_NIB_storage_data_f_9__51_),
	.b(FE_OFN465_n23476));
   oa12f01 U26134 (.o(n6033),
	.a(n22189),
	.b(FE_OFN465_n23476),
	.c(n23947));
   na02f01 U26135 (.o(n22190),
	.a(proc_input_NIB_storage_data_f_9__50_),
	.b(FE_OFN465_n23476));
   oa12f01 U26136 (.o(n6038),
	.a(n22190),
	.b(FE_OFN465_n23476),
	.c(n23903));
   na02f01 U26137 (.o(n22191),
	.a(proc_input_NIB_storage_data_f_9__49_),
	.b(FE_OFN101_n22098));
   na02f01 U26138 (.o(n22192),
	.a(proc_input_NIB_storage_data_f_9__39_),
	.b(FE_OFN465_n23476));
   na02f01 U26139 (.o(n22193),
	.a(proc_input_NIB_storage_data_f_9__48_),
	.b(FE_OFN101_n22098));
   oa12f01 U26140 (.o(n6048),
	.a(n22193),
	.b(FE_OFN101_n22098),
	.c(n23912));
   na02f01 U26141 (.o(n22194),
	.a(proc_input_NIB_storage_data_f_9__47_),
	.b(FE_OFN101_n22098));
   oa12f01 U26142 (.o(n6053),
	.a(n22194),
	.b(FE_OFN101_n22098),
	.c(n23914));
   na02f01 U26143 (.o(n22195),
	.a(proc_input_NIB_storage_data_f_9__46_),
	.b(FE_OFN101_n22098));
   oa12f01 U26144 (.o(n6058),
	.a(n22195),
	.b(FE_OFN101_n22098),
	.c(n23916));
   na02f01 U26145 (.o(n22196),
	.a(proc_input_NIB_storage_data_f_9__36_),
	.b(FE_OFN101_n22098));
   oa12f01 U26146 (.o(n6108),
	.a(n22196),
	.b(FE_OFN101_n22098),
	.c(n23940));
   na02f01 U26147 (.o(n22197),
	.a(proc_input_NIB_storage_data_f_9__37_),
	.b(FE_OFN101_n22098));
   oa12f01 U26148 (.o(n6103),
	.a(n22197),
	.b(FE_OFN101_n22098),
	.c(n23796));
   na02f01 U26149 (.o(n22198),
	.a(proc_input_NIB_storage_data_f_9__35_),
	.b(FE_OFN101_n22098));
   oa12f01 U26150 (.o(n6113),
	.a(n22198),
	.b(FE_OFN101_n22098),
	.c(n23944));
   na02f01 U26151 (.o(n22199),
	.a(proc_input_NIB_storage_data_f_9__25_),
	.b(FE_OFN101_n22098));
   oa12f01 U26152 (.o(n6163),
	.a(n22199),
	.b(FE_OFN101_n22098),
	.c(n23802));
   oa12f01 U26153 (.o(n6078),
	.a(n22200),
	.b(FE_OFN101_n22098),
	.c(n23808));
   na02f01 U26154 (.o(n22201),
	.a(proc_input_NIB_storage_data_f_9__26_),
	.b(FE_OFN101_n22098));
   oa12f01 U26155 (.o(n6158),
	.a(n22201),
	.b(FE_OFN101_n22098),
	.c(n23818));
   na02f01 U26156 (.o(n22202),
	.a(proc_input_NIB_storage_data_f_9__45_),
	.b(FE_OFN465_n23476));
   oa12f01 U26157 (.o(n6063),
	.a(n22202),
	.b(FE_OFN465_n23476),
	.c(n23942));
   na02f01 U26158 (.o(n22203),
	.a(proc_input_NIB_storage_data_f_9__28_),
	.b(FE_OFN101_n22098));
   oa12f01 U26159 (.o(n6148),
	.a(n22203),
	.b(FE_OFN101_n22098),
	.c(n23814));
   na02f01 U26160 (.o(n22204),
	.a(proc_input_NIB_storage_data_f_9__44_),
	.b(FE_OFN465_n23476));
   oa12f01 U26161 (.o(n6068),
	.a(n22204),
	.b(FE_OFN465_n23476),
	.c(n23920));
   na02f01 U26162 (.o(n22205),
	.a(proc_input_NIB_storage_data_f_9__43_),
	.b(FE_OFN101_n22098));
   oa12f01 U26163 (.o(n6073),
	.a(n22205),
	.b(FE_OFN101_n22098),
	.c(n23806));
   na02f01 U26164 (.o(n22206),
	.a(proc_input_NIB_storage_data_f_9__34_),
	.b(FE_OFN101_n22098));
   na02f01 U26165 (.o(n22207),
	.a(proc_input_NIB_storage_data_f_9__32_),
	.b(FE_OFN101_n22098));
   oa12f01 U26166 (.o(n6128),
	.a(n22207),
	.b(FE_OFN101_n22098),
	.c(n23905));
   na02f01 U26167 (.o(n22208),
	.a(proc_input_NIB_storage_data_f_9__30_),
	.b(FE_OFN101_n22098));
   oa12f01 U26168 (.o(n6138),
	.a(n22208),
	.b(FE_OFN101_n22098),
	.c(n23894));
   na02f01 U26169 (.o(n22209),
	.a(proc_input_NIB_storage_data_f_9__41_),
	.b(FE_OFN101_n22098));
   oa12f01 U26170 (.o(n6083),
	.a(n22209),
	.b(FE_OFN101_n22098),
	.c(n23928));
   na02f01 U26171 (.o(n22210),
	.a(proc_input_NIB_storage_data_f_9__40_),
	.b(FE_OFN465_n23476));
   oa12f01 U26172 (.o(n6088),
	.a(n22210),
	.b(FE_OFN465_n23476),
	.c(n23800));
   na02f01 U26173 (.o(n22211),
	.a(proc_input_NIB_storage_data_f_9__22_),
	.b(FE_OFN465_n23476));
   oa12f01 U26174 (.o(n6178),
	.a(n22211),
	.b(FE_OFN465_n23476),
	.c(n23820));
   na02f01 U26175 (.o(n22212),
	.a(proc_input_NIB_storage_data_f_9__29_),
	.b(FE_OFN101_n22098));
   oa12f01 U26176 (.o(n6143),
	.a(n22212),
	.b(FE_OFN101_n22098),
	.c(n23804));
   na02f01 U26177 (.o(n22213),
	.a(proc_input_NIB_storage_data_f_9__31_),
	.b(FE_OFN465_n23476));
   oa12f01 U26178 (.o(n6153),
	.a(n22214),
	.b(FE_OFN465_n23476),
	.c(n23822));
   na02f01 U26179 (.o(n22215),
	.a(proc_input_NIB_storage_data_f_8__51_),
	.b(n23471));
   oa12f01 U26180 (.o(n5713),
	.a(n22215),
	.b(n23471),
	.c(n23947));
   no02f01 U26181 (.o(north_input_control_N53),
	.a(FE_OFN5_reset),
	.b(n18112));
   na02f01 U26182 (.o(n22219),
	.a(n22218),
	.b(n22217));
   na02f02 U26183 (.o(n22223),
	.a(n22222),
	.b(n22221));
   in01s01 U26184 (.o(n22224),
	.a(n22223));
   na02f02 U26185 (.o(n22227),
	.a(n22226),
	.b(n22225));
   in01s01 U26186 (.o(n22228),
	.a(n22227));
   na02f01 U26187 (.o(n22231),
	.a(n22230),
	.b(n22229));
   in01s01 U26189 (.o(n22236),
	.a(n22235));
   oa22m01 U26190 (.o(n22237),
	.a(FE_OFN25787_n17770),
	.b(dataIn_S_4_),
	.c(south_input_NIB_storage_data_f_1__4_),
	.d(n20797));
   in01s01 U26191 (.o(n10138),
	.a(n22237));
   oa22s01 U26192 (.o(n22238),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_1_),
	.c(south_input_NIB_storage_data_f_0__1_),
	.d(FE_OFN83_n20814));
   in01s01 U26193 (.o(n9833),
	.a(n22238));
   oa22m01 U26194 (.o(n22239),
	.a(FE_OFN25787_n17770),
	.b(dataIn_S_7_),
	.c(south_input_NIB_storage_data_f_1__7_),
	.d(n20797));
   in01s01 U26195 (.o(n10123),
	.a(n22239));
   oa22m01 U26196 (.o(n22240),
	.a(FE_OFN25787_n17770),
	.b(dataIn_S_5_),
	.c(south_input_NIB_storage_data_f_1__5_),
	.d(n20797));
   in01s01 U26197 (.o(n10133),
	.a(n22240));
   oa22m01 U26198 (.o(n22241),
	.a(n17770),
	.b(dataIn_S_1_),
	.c(south_input_NIB_storage_data_f_1__1_),
	.d(n20797));
   in01s01 U26199 (.o(n10153),
	.a(n22241));
   oa22m01 U26200 (.o(n22242),
	.a(FE_OFN25787_n17770),
	.b(dataIn_S_2_),
	.c(south_input_NIB_storage_data_f_1__2_),
	.d(n20797));
   in01s01 U26201 (.o(n10148),
	.a(n22242));
   oa22m01 U26202 (.o(n22243),
	.a(FE_OFN25787_n17770),
	.b(dataIn_S_3_),
	.c(south_input_NIB_storage_data_f_1__3_),
	.d(n20797));
   in01s01 U26203 (.o(n10143),
	.a(n22243));
   oa22s01 U26204 (.o(n22244),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_0_),
	.c(south_input_NIB_storage_data_f_0__0_),
	.d(FE_OFN83_n20814));
   in01s01 U26205 (.o(n9838),
	.a(n22244));
   oa22m01 U26206 (.o(n22245),
	.a(FE_OFN25787_n17770),
	.b(dataIn_S_0_),
	.c(south_input_NIB_storage_data_f_1__0_),
	.d(n20797));
   in01s01 U26207 (.o(n10158),
	.a(n22245));
   oa22m01 U26208 (.o(n22246),
	.a(FE_OFN25787_n17770),
	.b(dataIn_S_6_),
	.c(south_input_NIB_storage_data_f_1__6_),
	.d(n20797));
   in01s01 U26209 (.o(n10128),
	.a(n22246));
   oa22s01 U26210 (.o(n22247),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_5_),
	.c(south_input_NIB_storage_data_f_0__5_),
	.d(FE_OFN83_n20814));
   in01s01 U26211 (.o(n9813),
	.a(n22247));
   oa22m01 U26212 (.o(n22248),
	.a(FE_OFN25787_n17770),
	.b(dataIn_S_9_),
	.c(south_input_NIB_storage_data_f_1__9_),
	.d(n20797));
   in01s01 U26213 (.o(n10113),
	.a(n22248));
   oa22m01 U26214 (.o(n22249),
	.a(FE_OFN25787_n17770),
	.b(dataIn_S_10_),
	.c(south_input_NIB_storage_data_f_1__10_),
	.d(n20797));
   in01s01 U26215 (.o(n10108),
	.a(n22249));
   oa22s01 U26216 (.o(n22250),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_11_),
	.c(south_input_NIB_storage_data_f_0__11_),
	.d(FE_OFN83_n20814));
   in01s01 U26217 (.o(n9783),
	.a(n22250));
   oa22s01 U26218 (.o(n22251),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_4_),
	.c(south_input_NIB_storage_data_f_0__4_),
	.d(FE_OFN83_n20814));
   in01s01 U26219 (.o(n9818),
	.a(n22251));
   oa22s01 U26220 (.o(n22252),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_3_),
	.c(south_input_NIB_storage_data_f_0__3_),
	.d(FE_OFN83_n20814));
   in01s01 U26221 (.o(n9823),
	.a(n22252));
   oa22s01 U26222 (.o(n22253),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_6_),
	.c(south_input_NIB_storage_data_f_0__6_),
	.d(FE_OFN83_n20814));
   in01s01 U26223 (.o(n9808),
	.a(n22253));
   in01s01 U26224 (.o(n9828),
	.a(n22254));
   oa22s01 U26225 (.o(n22255),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_9_),
	.c(south_input_NIB_storage_data_f_0__9_),
	.d(FE_OFN83_n20814));
   oa22s01 U26226 (.o(n22256),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_7_),
	.c(south_input_NIB_storage_data_f_0__7_),
	.d(FE_OFN83_n20814));
   in01s01 U26227 (.o(n9803),
	.a(n22256));
   oa22s01 U26228 (.o(n22257),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_10_),
	.c(south_input_NIB_storage_data_f_0__10_),
	.d(FE_OFN83_n20814));
   in01s01 U26229 (.o(n9788),
	.a(n22257));
   oa22m01 U26230 (.o(n22258),
	.a(FE_OFN25750_FE_OFN24796_n20854),
	.b(dataIn_W_8_),
	.c(west_input_NIB_storage_data_f_0__8_),
	.d(n20855));
   in01s01 U26231 (.o(n8508),
	.a(n22258));
   oa22m01 U26232 (.o(n22259),
	.a(FE_OFN25749_FE_OFN24796_n20854),
	.b(dataIn_W_2_),
	.c(west_input_NIB_storage_data_f_0__2_),
	.d(n20855));
   in01s01 U26233 (.o(n8538),
	.a(n22259));
   oa22m01 U26234 (.o(n22260),
	.a(FE_OFN25750_FE_OFN24796_n20854),
	.b(dataIn_W_6_),
	.c(west_input_NIB_storage_data_f_0__6_),
	.d(n20855));
   oa22m01 U26235 (.o(n22261),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_0_),
	.c(west_input_NIB_storage_data_f_1__0_),
	.d(FE_OFN380_n17772));
   in01s01 U26236 (.o(n8868),
	.a(n22261));
   oa22m01 U26237 (.o(n22262),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_2_),
	.c(west_input_NIB_storage_data_f_1__2_),
	.d(FE_OFN380_n17772));
   in01s01 U26238 (.o(n8858),
	.a(n22262));
   oa22m01 U26239 (.o(n22263),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_6_),
	.c(west_input_NIB_storage_data_f_1__6_),
	.d(FE_OFN380_n17772));
   in01s01 U26240 (.o(n8838),
	.a(n22263));
   oa22m01 U26241 (.o(n22264),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_5_),
	.c(west_input_NIB_storage_data_f_1__5_),
	.d(FE_OFN380_n17772));
   in01s01 U26242 (.o(n8843),
	.a(n22264));
   oa22m01 U26243 (.o(n22265),
	.a(FE_OFN25750_FE_OFN24796_n20854),
	.b(dataIn_W_3_),
	.c(west_input_NIB_storage_data_f_0__3_),
	.d(n20855));
   in01s01 U26244 (.o(n8533),
	.a(n22265));
   in01s01 U26245 (.o(n8853),
	.a(n22266));
   oa22m01 U26246 (.o(n22267),
	.a(FE_OFN25749_FE_OFN24796_n20854),
	.b(dataIn_W_5_),
	.c(west_input_NIB_storage_data_f_0__5_),
	.d(n20855));
   in01s01 U26247 (.o(n8523),
	.a(n22267));
   oa22m01 U26248 (.o(n22268),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_8_),
	.c(west_input_NIB_storage_data_f_1__8_),
	.d(FE_OFN380_n17772));
   in01s01 U26249 (.o(n8828),
	.a(n22268));
   oa22m01 U26250 (.o(n22269),
	.a(FE_OFN25750_FE_OFN24796_n20854),
	.b(dataIn_W_0_),
	.c(west_input_NIB_storage_data_f_0__0_),
	.d(n20855));
   in01s01 U26251 (.o(n8548),
	.a(n22269));
   na02f02 U26252 (.o(n25977),
	.a(proc_input_NIB_tail_ptr_f_2_),
	.b(n25980));
   no02f01 U26253 (.o(east_input_control_N53),
	.a(FE_OFN5_reset),
	.b(n25017));
   na02f01 U26254 (.o(n22285),
	.a(n22284),
	.b(n22283));
   na03m02 U26256 (.o(dataOut_S_50_),
	.a(n22289),
	.b(n22288),
	.c(n22287));
   na03f06 U26257 (.o(dataOut_S_44_),
	.a(n22292),
	.b(n22291),
	.c(n22290));
   na03m02 U26258 (.o(dataOut_S_63_),
	.a(n22296),
	.b(n22295),
	.c(n22294));
   ao22f01 U26259 (.o(n22298),
	.a(n25498),
	.b(n23534),
	.c(FE_OFN93_n21667),
	.d(n23535));
   na03m02 U26260 (.o(FE_OFN703_dataOut_S_25),
	.a(n22299),
	.b(n22298),
	.c(n22297));
   ao22f01 U26261 (.o(n22301),
	.a(n25498),
	.b(n23527),
	.c(FE_OFN105_n22517),
	.d(n23526));
   na03f01 U26262 (.o(FE_OFN701_dataOut_S_26),
	.a(n22302),
	.b(n22301),
	.c(n22300));
   na03f04 U26263 (.o(dataOut_S_45_),
	.a(n22305),
	.b(n22304),
	.c(n22303));
   na03m02 U26264 (.o(dataOut_S_53_),
	.a(n22311),
	.b(n22310),
	.c(n22309));
   na03f01 U26265 (.o(FE_OFN677_dataOut_S_43),
	.a(n22314),
	.b(n22313),
	.c(n22312));
   na03f02 U26266 (.o(dataOut_S_55_),
	.a(n22317),
	.b(n22316),
	.c(n22315));
   na03f03 U26267 (.o(dataOut_S_46_),
	.a(n22320),
	.b(n22319),
	.c(n22318));
   ao22f01 U26268 (.o(n22323),
	.a(FE_OFN105_n22517),
	.b(n23481),
	.c(n25498),
	.d(n23478));
   na03f02 U26269 (.o(dataOut_S_30_),
	.a(n22323),
	.b(n22322),
	.c(n22321));
   ao22f01 U26270 (.o(n22326),
	.a(n19493),
	.b(n23517),
	.c(FE_OFN93_n21667),
	.d(n23516));
   ao22f01 U26271 (.o(n22325),
	.a(n25498),
	.b(n23519),
	.c(FE_OFN105_n22517),
	.d(n23518));
   na03m02 U26272 (.o(dataOut_S_51_),
	.a(n22329),
	.b(n22328),
	.c(n22327));
   na03f03 U26273 (.o(dataOut_S_47_),
	.a(n22332),
	.b(n22331),
	.c(n22330));
   in01s01 U26274 (.o(n12403),
	.a(n22333));
   in01s01 U26275 (.o(n12413),
	.a(n22334));
   in01s01 U26276 (.o(n12383),
	.a(n22335));
   in01s01 U26277 (.o(n12378),
	.a(n22337));
   in01s01 U26278 (.o(n12408),
	.a(n22338));
   in01s01 U26279 (.o(n12368),
	.a(n22339));
   in01s01 U26280 (.o(n12398),
	.a(n22340));
   in01s01 U26281 (.o(n12373),
	.a(n22341));
   in01s01 U26282 (.o(n12393),
	.a(n22342));
   ao22f01 U26283 (.o(n22344),
	.a(n17755),
	.b(FE_OFN473_n23560),
	.c(FE_OFN111_n22773),
	.d(FE_OFN130_n23559));
   in01s01 U26284 (.o(n22346),
	.a(n22345));
   ao22f01 U26285 (.o(n22348),
	.a(n17755),
	.b(n23569),
	.c(FE_OFN111_n22773),
	.d(n23568));
   na02f02 U26286 (.o(n22349),
	.a(n22348),
	.b(n22347));
   in01s01 U26287 (.o(n22350),
	.a(n22349));
   ao22f01 U26288 (.o(n22352),
	.a(FE_OFN389_n17786),
	.b(n24020),
	.c(FE_OFN111_n22773),
	.d(FE_OFN151_n24019));
   na02f02 U26289 (.o(n22353),
	.a(n22352),
	.b(n22351));
   ao22f01 U26291 (.o(n22356),
	.a(FE_OFN389_n17786),
	.b(FE_OFN485_n24011),
	.c(FE_OFN111_n22773),
	.d(FE_OFN146_n24010));
   na02f02 U26292 (.o(n22357),
	.a(n22356),
	.b(n22355));
   ao22m02 U26294 (.o(n22360),
	.a(FE_OFN389_n17786),
	.b(n23147),
	.c(n17755),
	.d(n23146));
   na02f02 U26295 (.o(n22361),
	.a(n22360),
	.b(n22359));
   in01s01 U26296 (.o(n22362),
	.a(n22361));
   ao22f01 U26297 (.o(n22364),
	.a(FE_OFN389_n17786),
	.b(n23975),
	.c(FE_OFN111_n22773),
	.d(n23974));
   na02f02 U26298 (.o(n22365),
	.a(n22364),
	.b(n22363));
   ao22f01 U26300 (.o(n22367),
	.a(n17786),
	.b(n23580),
	.c(FE_OFN111_n22773),
	.d(n23579));
   na02f02 U26301 (.o(n22369),
	.a(n22368),
	.b(n22367));
   in01s01 U26302 (.o(n22370),
	.a(n22369));
   no02f01 U26303 (.o(south_input_control_N53),
	.a(FE_OFN5_reset),
	.b(n25030));
   in01s01 U26304 (.o(n22385),
	.a(east_output_space_count_f_1_));
   no02m01 U26306 (.o(n22389),
	.a(east_output_space_yummy_f),
	.b(n22371));
   na02m01 U26307 (.o(n22377),
	.a(n22389),
	.b(n22388));
   no02m01 U26308 (.o(n22372),
	.a(east_output_space_count_f_1_),
	.b(n22377));
   in01s01 U26309 (.o(n22384),
	.a(east_output_space_count_f_2_));
   na02s01 U26311 (.o(n22375),
	.a(east_output_space_count_f_2_),
	.b(n22385));
   in01s01 U26312 (.o(n22383),
	.a(n22375));
   in01s01 U26313 (.o(n22380),
	.a(n22376));
   na02s01 U26314 (.o(n22378),
	.a(east_output_space_count_f_1_),
	.b(n22377));
   na02s01 U26315 (.o(n22379),
	.a(n22392),
	.b(n22378));
   na02f01 U26316 (.o(east_output_space_N48),
	.a(n22382),
	.b(n25818));
   no02s01 U26317 (.o(n22387),
	.a(east_output_space_valid_f),
	.b(n22383));
   na02s01 U26318 (.o(n22386),
	.a(n22385),
	.b(n22384));
   ao22s01 U26319 (.o(n22390),
	.a(east_output_space_yummy_f),
	.b(n22387),
	.c(n22389),
	.d(n22386));
   na02s01 U26320 (.o(n25817),
	.a(n22392),
	.b(n22391));
   in01s01 U26321 (.o(n10448),
	.a(n22393));
   oa22f01 U26322 (.o(n22394),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_10_),
	.c(south_input_NIB_storage_data_f_2__10_),
	.d(n20972));
   in01s01 U26323 (.o(n10428),
	.a(n22394));
   in01s01 U26324 (.o(n10753),
	.a(n22395));
   in01s01 U26325 (.o(n10793),
	.a(n22396));
   in01s01 U26326 (.o(n10788),
	.a(n22398));
   in01s01 U26327 (.o(n10783),
	.a(n22399));
   oa22f01 U26328 (.o(n22400),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_11_),
	.c(south_input_NIB_storage_data_f_2__11_),
	.d(n20972));
   in01s01 U26329 (.o(n10423),
	.a(n22400));
   in01s01 U26330 (.o(n10743),
	.a(n22401));
   in01s01 U26331 (.o(n10773),
	.a(n22402));
   in01s01 U26332 (.o(n10763),
	.a(n22404));
   in01s01 U26333 (.o(n10798),
	.a(n22405));
   in01s01 U26334 (.o(n10478),
	.a(n22406));
   oa22f01 U26335 (.o(n22407),
	.a(n25905),
	.b(dataIn_S_9_),
	.c(south_input_NIB_storage_data_f_2__9_),
	.d(n20972));
   in01s01 U26336 (.o(n10433),
	.a(n22407));
   in01s01 U26337 (.o(n10458),
	.a(n22408));
   in01s01 U26338 (.o(n10453),
	.a(n22409));
   in01s01 U26339 (.o(n10473),
	.a(n22410));
   in01s01 U26340 (.o(n10748),
	.a(n22411));
   in01s01 U26342 (.o(n10463),
	.a(n22413));
   in01s01 U26343 (.o(n10443),
	.a(n22414));
   oa22f01 U26344 (.o(n22415),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_2_),
	.c(west_input_NIB_storage_data_f_2__2_),
	.d(n25945));
   in01s01 U26345 (.o(n9178),
	.a(n22415));
   oa22f01 U26346 (.o(n22416),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_2_),
	.c(west_input_NIB_storage_data_f_3__2_),
	.d(n21070));
   in01s01 U26347 (.o(n9498),
	.a(n22416));
   in01s01 U26348 (.o(n9468),
	.a(n22417));
   oa22f01 U26349 (.o(n22418),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_3_),
	.c(west_input_NIB_storage_data_f_2__3_),
	.d(n25945));
   in01s01 U26350 (.o(n9173),
	.a(n22418));
   oa22f01 U26351 (.o(n22420),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_6_),
	.c(west_input_NIB_storage_data_f_2__6_),
	.d(n25945));
   in01s01 U26352 (.o(n9158),
	.a(n22420));
   in01s01 U26353 (.o(n9188),
	.a(n22421));
   oa22f01 U26354 (.o(n22422),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_6_),
	.c(west_input_NIB_storage_data_f_3__6_),
	.d(n21070));
   in01s01 U26355 (.o(n9478),
	.a(n22422));
   in01s01 U26356 (.o(n9163),
	.a(n22423));
   oa22f01 U26357 (.o(n22424),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_8_),
	.c(west_input_NIB_storage_data_f_2__8_),
	.d(n25945));
   in01s01 U26358 (.o(n9148),
	.a(n22424));
   in01s01 U26359 (.o(n9508),
	.a(n22425));
   oa22f01 U26360 (.o(n22426),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_5_),
	.c(west_input_NIB_storage_data_f_3__5_),
	.d(n21070));
   in01s01 U26361 (.o(n9483),
	.a(n22426));
   na02s01 U26362 (.o(n22427),
	.a(south_input_NIB_storage_data_f_0__51_),
	.b(FE_OFN403_n20815));
   oa12s01 U26363 (.o(n9583),
	.a(n22427),
	.b(FE_OFN403_n20815),
	.c(n22484));
   na02f01 U26364 (.o(n22428),
	.a(west_input_NIB_storage_data_f_0__53_),
	.b(FE_OFN25748_FE_OFN24796_n20854));
   oa12f01 U26365 (.o(n8283),
	.a(n22428),
	.b(FE_OFN25748_FE_OFN24796_n20854),
	.c(n22488));
   na02m01 U26366 (.o(n22429),
	.a(south_input_NIB_storage_data_f_1__51_),
	.b(FE_OFN899_n17770));
   oa12s01 U26367 (.o(n9903),
	.a(n22429),
	.b(FE_OFN899_n17770),
	.c(n22484));
   na02f01 U26368 (.o(n22430),
	.a(west_input_NIB_storage_data_f_1__53_),
	.b(FE_OFN381_n17772));
   oa12f01 U26369 (.o(n8603),
	.a(n22430),
	.b(FE_OFN381_n17772),
	.c(n22488));
   ao22f01 U26370 (.o(n22432),
	.a(n19493),
	.b(n24020),
	.c(FE_OFN577_n25498),
	.d(FE_OFN151_n24019));
   ao22f01 U26371 (.o(n22431),
	.a(FE_OFN105_n22517),
	.b(n24021),
	.c(FE_OFN93_n21667),
	.d(FE_OFN491_n24022));
   na02f02 U26372 (.o(n22433),
	.a(n22432),
	.b(n22431));
   ao22m01 U26374 (.o(n22435),
	.a(n25498),
	.b(n24030),
	.c(FE_OFN93_n21667),
	.d(n24031));
   na02f02 U26375 (.o(n22437),
	.a(n22436),
	.b(n22435));
   ao22m01 U26376 (.o(n22439),
	.a(n17755),
	.b(n24031),
	.c(FE_OFN111_n22773),
	.d(n24030));
   na02f01 U26377 (.o(n22441),
	.a(n22440),
	.b(n22439));
   in01s01 U26378 (.o(n22442),
	.a(n22441));
   na02s01 U26379 (.o(n22443),
	.a(north_input_NIB_storage_data_f_0__61_),
	.b(n17771));
   oa12s01 U26380 (.o(n12113),
	.a(n22443),
	.b(n17771),
	.c(n22444));
   in01s01 U26381 (.o(n13368),
	.a(n22445));
   in01s01 U26382 (.o(n13363),
	.a(n22446));
   in01s01 U26383 (.o(n13358),
	.a(n22447));
   oa22f01 U26384 (.o(n22448),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_33_),
	.c(north_input_NIB_storage_data_f_3__33_),
	.d(n21175));
   in01s01 U26385 (.o(n13213),
	.a(n22448));
   in01s01 U26386 (.o(n13378),
	.a(n22449));
   in01s01 U26387 (.o(n13328),
	.a(n22450));
   in01s01 U26388 (.o(n13338),
	.a(n22451));
   in01s01 U26389 (.o(n13353),
	.a(n22452));
   in01s01 U26390 (.o(n13373),
	.a(n22453));
   oa22f01 U26391 (.o(n22454),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_20_),
	.c(north_input_NIB_storage_data_f_3__20_),
	.d(n21175));
   in01s01 U26392 (.o(n13278),
	.a(n22454));
   oa22f01 U26393 (.o(n22455),
	.a(n25836),
	.b(dataIn_N_15_),
	.c(north_input_NIB_storage_data_f_3__15_),
	.d(n21175));
   in01s01 U26394 (.o(n13303),
	.a(n22455));
   in01s01 U26395 (.o(n13343),
	.a(n22456));
   in01s01 U26396 (.o(n13333),
	.a(n22457));
   oa22f01 U26397 (.o(n22458),
	.a(n25836),
	.b(dataIn_N_12_),
	.c(north_input_NIB_storage_data_f_3__12_),
	.d(n21175));
   in01s01 U26398 (.o(n13293),
	.a(n22459));
   in01s01 U26399 (.o(n13323),
	.a(n22460));
   oa22f01 U26400 (.o(n22461),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_14_),
	.c(north_input_NIB_storage_data_f_3__14_),
	.d(n21175));
   in01s01 U26401 (.o(n13308),
	.a(n22461));
   oa22f01 U26402 (.o(n22462),
	.a(FE_OFN86_n21175),
	.b(dataIn_N_16_),
	.c(north_input_NIB_storage_data_f_3__16_),
	.d(n21175));
   in01s01 U26403 (.o(n13298),
	.a(n22462));
   oa22f01 U26404 (.o(n22463),
	.a(n25848),
	.b(dataIn_N_16_),
	.c(north_input_NIB_storage_data_f_1__16_),
	.d(n21220));
   in01s01 U26405 (.o(n12658),
	.a(n22463));
   in01s01 U26406 (.o(n12688),
	.a(n22464));
   oa22f01 U26407 (.o(n22465),
	.a(n25848),
	.b(dataIn_N_14_),
	.c(north_input_NIB_storage_data_f_1__14_),
	.d(n21220));
   in01s01 U26408 (.o(n12668),
	.a(n22465));
   oa22f01 U26409 (.o(n22466),
	.a(n25848),
	.b(dataIn_N_17_),
	.c(north_input_NIB_storage_data_f_1__17_),
	.d(n21220));
   in01s01 U26410 (.o(n12653),
	.a(n22466));
   oa22f01 U26411 (.o(n22467),
	.a(n25848),
	.b(dataIn_N_12_),
	.c(north_input_NIB_storage_data_f_1__12_),
	.d(n21220));
   in01s01 U26412 (.o(n12678),
	.a(n22467));
   oa22f01 U26413 (.o(n22469),
	.a(n25848),
	.b(dataIn_N_5_),
	.c(north_input_NIB_storage_data_f_1__5_),
	.d(n21220));
   in01s01 U26414 (.o(n12713),
	.a(n22469));
   in01s01 U26415 (.o(n12693),
	.a(n22470));
   oa22f01 U26416 (.o(n22471),
	.a(n25848),
	.b(dataIn_N_11_),
	.c(north_input_NIB_storage_data_f_1__11_),
	.d(n21220));
   in01s01 U26417 (.o(n12683),
	.a(n22471));
   in01s01 U26418 (.o(n12728),
	.a(n22472));
   oa22f01 U26419 (.o(n22473),
	.a(n25848),
	.b(dataIn_N_33_),
	.c(north_input_NIB_storage_data_f_1__33_),
	.d(n21220));
   in01s01 U26420 (.o(n12573),
	.a(n22473));
   in01s01 U26421 (.o(n12738),
	.a(n22474));
   in01s01 U26422 (.o(n12638),
	.a(n22475));
   in01s01 U26423 (.o(n12733),
	.a(n22476));
   oa22f01 U26424 (.o(n22477),
	.a(n25848),
	.b(dataIn_N_7_),
	.c(north_input_NIB_storage_data_f_1__7_),
	.d(n21220));
   in01s01 U26425 (.o(n12703),
	.a(n22477));
   oa22f01 U26426 (.o(n22478),
	.a(n25848),
	.b(dataIn_N_15_),
	.c(north_input_NIB_storage_data_f_1__15_),
	.d(n21220));
   in01s01 U26427 (.o(n12663),
	.a(n22478));
   in01s01 U26428 (.o(n12723),
	.a(n22479));
   oa22f01 U26429 (.o(n22480),
	.a(n25848),
	.b(dataIn_N_8_),
	.c(north_input_NIB_storage_data_f_1__8_),
	.d(n21220));
   in01s01 U26430 (.o(n12698),
	.a(n22480));
   na02f01 U26431 (.o(n22481),
	.a(south_input_NIB_storage_data_f_2__52_),
	.b(n25905));
   oa12f01 U26432 (.o(n10218),
	.a(n22481),
	.b(n25905),
	.c(n22482));
   na02s01 U26433 (.o(n22483),
	.a(south_input_NIB_storage_data_f_3__51_),
	.b(FE_OFN896_n17769));
   na02f01 U26434 (.o(n22485),
	.a(west_input_NIB_storage_data_f_2__44_),
	.b(FE_OFN25792_n21053));
   na02f01 U26435 (.o(n22487),
	.a(west_input_NIB_storage_data_f_3__53_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U26436 (.o(n9243),
	.a(n22487),
	.b(n22488),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   in01s01 U26437 (.o(n22500),
	.a(south_input_control_count_f_5_));
   na02s01 U26438 (.o(n22495),
	.a(n23553),
	.b(n22912));
   na02s01 U26439 (.o(n22498),
	.a(n23553),
	.b(n23308));
   no02f01 U26440 (.o(n22497),
	.a(FE_OFN5_reset),
	.b(n22496));
   oa12f01 U26441 (.o(n22499),
	.a(n22497),
	.b(n25250),
	.c(n22498));
   ao12f01 U26442 (.o(south_input_control_N46),
	.a(n22499),
	.b(n22911),
	.c(n22500));
   na02f02 U26443 (.o(n22503),
	.a(n22502),
	.b(n22501));
   in01s01 U26444 (.o(n22504),
	.a(n22503));
   ao22m01 U26445 (.o(n22505),
	.a(n25498),
	.b(FE_OFN136_n23623),
	.c(FE_OFN105_n22517),
	.d(n23622));
   na02f02 U26446 (.o(n22507),
	.a(n22506),
	.b(n22505));
   in01s01 U26447 (.o(n22508),
	.a(n22507));
   ao22f01 U26448 (.o(n22509),
	.a(n25498),
	.b(FE_OFN140_n23959),
	.c(FE_OFN105_n22517),
	.d(n23958));
   na02f02 U26449 (.o(n22511),
	.a(n22510),
	.b(n22509));
   in01f01 U26450 (.o(n22512),
	.a(n22511));
   ao22f01 U26451 (.o(n22514),
	.a(FE_OFN105_n22517),
	.b(n23632),
	.c(FE_OFN577_n25498),
	.d(n23629));
   na02f01 U26452 (.o(n22515),
	.a(n22514),
	.b(n22513));
   in01s01 U26453 (.o(n22516),
	.a(n22515));
   no02f01 U26455 (.o(n22522),
	.a(n22521),
	.b(n22520));
   na02f02 U26456 (.o(n22528),
	.a(n22527),
	.b(n22526));
   in01s01 U26457 (.o(n22529),
	.a(n22528));
   oa12f01 U26458 (.o(FE_OFN759_dataOut_W_38),
	.a(n22532),
	.b(n18031),
	.c(FE_OFN25880_n19446));
   no02f02 U26460 (.o(n22536),
	.a(FE_OFN418_n22535),
	.b(n22534));
   in01s01 U26461 (.o(n22704),
	.a(dataIn_S_47_));
   na02s01 U26462 (.o(n22540),
	.a(south_input_NIB_storage_data_f_0__47_),
	.b(FE_OFN952_n25916));
   oa12s01 U26463 (.o(n9603),
	.a(n22540),
	.b(FE_OFN952_n25916),
	.c(n22704));
   na02s01 U26464 (.o(n22541),
	.a(south_input_NIB_storage_data_f_0__63_),
	.b(FE_OFN403_n20815));
   oa12s01 U26465 (.o(n9523),
	.a(n22541),
	.b(FE_OFN403_n20815),
	.c(n22686));
   in01s01 U26466 (.o(n22696),
	.a(dataIn_S_35_));
   na02s01 U26467 (.o(n22542),
	.a(south_input_NIB_storage_data_f_0__35_),
	.b(FE_OFN952_n25916));
   oa12s01 U26468 (.o(n9663),
	.a(n22542),
	.b(FE_OFN952_n25916),
	.c(n22696));
   in01s01 U26469 (.o(n22694),
	.a(dataIn_S_45_));
   na02s01 U26470 (.o(n22543),
	.a(south_input_NIB_storage_data_f_0__45_),
	.b(FE_OFN952_n25916));
   oa12s01 U26471 (.o(n9613),
	.a(n22543),
	.b(FE_OFN952_n25916),
	.c(n22694));
   in01s01 U26472 (.o(n22682),
	.a(dataIn_S_37_));
   na02s01 U26473 (.o(n22544),
	.a(south_input_NIB_storage_data_f_0__37_),
	.b(FE_OFN952_n25916));
   oa12s01 U26474 (.o(n9653),
	.a(n22544),
	.b(FE_OFN952_n25916),
	.c(n22682));
   in01s01 U26475 (.o(n22702),
	.a(dataIn_S_32_));
   na02s01 U26476 (.o(n22545),
	.a(south_input_NIB_storage_data_f_0__32_),
	.b(FE_OFN952_n25916));
   oa12s01 U26477 (.o(n9678),
	.a(n22545),
	.b(FE_OFN952_n25916),
	.c(n22702));
   in01s01 U26478 (.o(n22677),
	.a(dataIn_S_42_));
   na02s01 U26479 (.o(n22546),
	.a(south_input_NIB_storage_data_f_0__42_),
	.b(FE_OFN952_n25916));
   oa12s01 U26480 (.o(n9628),
	.a(n22546),
	.b(FE_OFN952_n25916),
	.c(n22677));
   na02s01 U26481 (.o(n22547),
	.a(south_input_NIB_storage_data_f_0__39_),
	.b(FE_OFN952_n25916));
   in01s01 U26482 (.o(n22692),
	.a(dataIn_S_43_));
   na02s01 U26483 (.o(n22548),
	.a(south_input_NIB_storage_data_f_0__43_),
	.b(FE_OFN952_n25916));
   oa12s01 U26484 (.o(n9623),
	.a(n22548),
	.b(FE_OFN952_n25916),
	.c(n22692));
   in01s01 U26485 (.o(n22700),
	.a(dataIn_S_44_));
   na02s01 U26486 (.o(n22549),
	.a(south_input_NIB_storage_data_f_0__44_),
	.b(FE_OFN952_n25916));
   oa12s01 U26487 (.o(n9618),
	.a(n22549),
	.b(FE_OFN952_n25916),
	.c(n22700));
   in01s01 U26488 (.o(n22706),
	.a(dataIn_S_36_));
   na02s01 U26489 (.o(n22550),
	.a(south_input_NIB_storage_data_f_0__36_),
	.b(FE_OFN953_n25916));
   oa12s01 U26490 (.o(n9658),
	.a(n22550),
	.b(FE_OFN952_n25916),
	.c(n22706));
   in01s01 U26491 (.o(n22698),
	.a(dataIn_S_31_));
   na02s01 U26492 (.o(n22551),
	.a(south_input_NIB_storage_data_f_0__31_),
	.b(FE_OFN953_n25916));
   oa12s01 U26493 (.o(n9683),
	.a(n22551),
	.b(FE_OFN952_n25916),
	.c(n22698));
   na02s01 U26494 (.o(n22552),
	.a(south_input_NIB_storage_data_f_0__34_),
	.b(n20815));
   oa12s01 U26495 (.o(n9668),
	.a(n22552),
	.b(FE_OFN952_n25916),
	.c(n22667));
   in01s01 U26496 (.o(n22684),
	.a(dataIn_S_46_));
   na02s01 U26497 (.o(n22553),
	.a(south_input_NIB_storage_data_f_0__46_),
	.b(FE_OFN82_n20814));
   oa12s01 U26498 (.o(n9608),
	.a(n22553),
	.b(FE_OFN952_n25916),
	.c(n22684));
   in01s01 U26499 (.o(n22745),
	.a(dataIn_W_23_));
   na02s01 U26500 (.o(n22554),
	.a(west_input_NIB_storage_data_f_0__23_),
	.b(FE_OFN1084_n20854));
   oa12s01 U26501 (.o(n8433),
	.a(n22554),
	.b(FE_OFN25751_FE_OFN24796_n20854),
	.c(n22745));
   in01s01 U26502 (.o(n22747),
	.a(dataIn_W_30_));
   na02s01 U26503 (.o(n22555),
	.a(west_input_NIB_storage_data_f_0__30_),
	.b(FE_OFN1084_n20854));
   oa12f01 U26504 (.o(n8398),
	.a(n22555),
	.b(FE_OFN25747_FE_OFN24796_n20854),
	.c(n22747));
   na02s01 U26505 (.o(n22556),
	.a(west_input_NIB_storage_data_f_0__54_),
	.b(FE_OFN1084_n20854));
   oa12f01 U26506 (.o(n8278),
	.a(n22556),
	.b(FE_OFN25748_FE_OFN24796_n20854),
	.c(n22557));
   in01f01 U26507 (.o(n22741),
	.a(dataIn_W_57_));
   na02s01 U26508 (.o(n22558),
	.a(west_input_NIB_storage_data_f_0__57_),
	.b(FE_OFN24795_n20854));
   oa12s01 U26509 (.o(n8263),
	.a(n22558),
	.b(FE_OFN25750_FE_OFN24796_n20854),
	.c(n22741));
   in01s01 U26510 (.o(n22730),
	.a(dataIn_W_58_));
   na02s01 U26511 (.o(n22559),
	.a(west_input_NIB_storage_data_f_0__58_),
	.b(FE_OFN1084_n20854));
   oa12f01 U26512 (.o(n8258),
	.a(n22559),
	.b(FE_OFN25748_FE_OFN24796_n20854),
	.c(n22730));
   in01s01 U26513 (.o(n22734),
	.a(dataIn_W_59_));
   na02s01 U26514 (.o(n22560),
	.a(west_input_NIB_storage_data_f_0__59_),
	.b(FE_OFN1084_n20854));
   oa12f01 U26515 (.o(n8253),
	.a(n22560),
	.b(FE_OFN25748_FE_OFN24796_n20854),
	.c(n22734));
   oa12f01 U26516 (.o(n8423),
	.a(n22561),
	.b(FE_OFN24796_n20854),
	.c(n22726));
   in01s01 U26517 (.o(n22724),
	.a(dataIn_W_55_));
   na02s01 U26518 (.o(n22562),
	.a(west_input_NIB_storage_data_f_0__55_),
	.b(FE_OFN1084_n20854));
   oa12f01 U26519 (.o(n8273),
	.a(n22562),
	.b(FE_OFN25748_FE_OFN24796_n20854),
	.c(n22724));
   in01s01 U26520 (.o(n22732),
	.a(dataIn_W_22_));
   na02s01 U26521 (.o(n22563),
	.a(west_input_NIB_storage_data_f_0__22_),
	.b(FE_OFN1084_n20854));
   oa12s01 U26522 (.o(n8438),
	.a(n22563),
	.b(FE_OFN25747_FE_OFN24796_n20854),
	.c(n22732));
   na02s01 U26523 (.o(n22564),
	.a(west_input_NIB_storage_data_f_0__26_),
	.b(n25965));
   oa12s01 U26524 (.o(n8418),
	.a(n22564),
	.b(FE_OFN24796_n20854),
	.c(n22751));
   in01s01 U26525 (.o(n22712),
	.a(dataIn_W_28_));
   na02s01 U26526 (.o(n22565),
	.a(west_input_NIB_storage_data_f_0__28_),
	.b(FE_OFN1089_n20855));
   oa12s01 U26527 (.o(n8408),
	.a(n22565),
	.b(FE_OFN25749_FE_OFN24796_n20854),
	.c(n22712));
   na02s01 U26528 (.o(n22566),
	.a(west_input_NIB_storage_data_f_0__46_),
	.b(FE_OFN1084_n20854));
   oa12f01 U26529 (.o(n8318),
	.a(n22566),
	.b(FE_OFN25747_FE_OFN24796_n20854),
	.c(n22743));
   na02s01 U26530 (.o(n22567),
	.a(west_input_NIB_storage_data_f_0__24_),
	.b(FE_OFN1083_n20854));
   oa12s01 U26531 (.o(n8428),
	.a(n22567),
	.b(FE_OFN25751_FE_OFN24796_n20854),
	.c(n22736));
   in01s01 U26532 (.o(n22728),
	.a(dataIn_W_27_));
   na02s01 U26533 (.o(n22568),
	.a(west_input_NIB_storage_data_f_0__27_),
	.b(FE_OFN1084_n20854));
   oa12s01 U26534 (.o(n8413),
	.a(n22568),
	.b(FE_OFN25751_FE_OFN24796_n20854),
	.c(n22728));
   na02s01 U26535 (.o(n22569),
	.a(south_input_NIB_storage_data_f_1__47_),
	.b(FE_OFN25785_n17770));
   oa12s01 U26536 (.o(n9923),
	.a(n22569),
	.b(FE_OFN25785_n17770),
	.c(n22704));
   na02f01 U26537 (.o(n22570),
	.a(south_input_NIB_storage_data_f_1__44_),
	.b(FE_OFN25785_n17770));
   oa12s01 U26538 (.o(n9938),
	.a(n22570),
	.b(FE_OFN25785_n17770),
	.c(n22700));
   na02s01 U26539 (.o(n22571),
	.a(south_input_NIB_storage_data_f_1__34_),
	.b(FE_OFN25785_n17770));
   oa12s01 U26540 (.o(n9988),
	.a(n22571),
	.b(FE_OFN25785_n17770),
	.c(n22667));
   na02s01 U26541 (.o(n22572),
	.a(south_input_NIB_storage_data_f_1__46_),
	.b(FE_OFN25785_n17770));
   oa12s01 U26542 (.o(n9928),
	.a(n22572),
	.b(FE_OFN25785_n17770),
	.c(n22684));
   na02f01 U26543 (.o(n22573),
	.a(south_input_NIB_storage_data_f_1__36_),
	.b(FE_OFN25785_n17770));
   oa12s01 U26544 (.o(n9978),
	.a(n22573),
	.b(FE_OFN25785_n17770),
	.c(n22706));
   na02f02 U26545 (.o(n22574),
	.a(south_input_NIB_storage_data_f_1__45_),
	.b(FE_OFN25785_n17770));
   oa12s01 U26546 (.o(n9933),
	.a(n22574),
	.b(FE_OFN25785_n17770),
	.c(n22694));
   na02s01 U26547 (.o(n22575),
	.a(south_input_NIB_storage_data_f_1__63_),
	.b(FE_OFN25849_FE_OFN899_n17770));
   oa12s01 U26548 (.o(n9843),
	.a(n22575),
	.b(FE_OFN25849_FE_OFN899_n17770),
	.c(n22686));
   na02s01 U26549 (.o(n22576),
	.a(south_input_NIB_storage_data_f_1__43_),
	.b(FE_OFN25785_n17770));
   na02f01 U26550 (.o(n22577),
	.a(south_input_NIB_storage_data_f_1__32_),
	.b(FE_OFN25785_n17770));
   oa12s01 U26551 (.o(n9998),
	.a(n22577),
	.b(FE_OFN25785_n17770),
	.c(n22702));
   na02f02 U26552 (.o(n22578),
	.a(south_input_NIB_storage_data_f_1__31_),
	.b(FE_OFN25785_n17770));
   oa12s01 U26553 (.o(n10003),
	.a(n22578),
	.b(FE_OFN25785_n17770),
	.c(n22698));
   na02f01 U26554 (.o(n22579),
	.a(south_input_NIB_storage_data_f_1__35_),
	.b(FE_OFN25785_n17770));
   oa12s01 U26555 (.o(n9983),
	.a(n22579),
	.b(FE_OFN25785_n17770),
	.c(n22696));
   na02f01 U26556 (.o(n22580),
	.a(south_input_NIB_storage_data_f_1__37_),
	.b(FE_OFN25785_n17770));
   oa12s01 U26557 (.o(n9973),
	.a(n22580),
	.b(FE_OFN25785_n17770),
	.c(n22682));
   na02f01 U26558 (.o(n22581),
	.a(south_input_NIB_storage_data_f_1__39_),
	.b(FE_OFN25785_n17770));
   oa12s01 U26559 (.o(n9963),
	.a(n22581),
	.b(FE_OFN25785_n17770),
	.c(n22582));
   na02f01 U26560 (.o(n22583),
	.a(south_input_NIB_storage_data_f_1__42_),
	.b(FE_OFN25785_n17770));
   oa12s01 U26561 (.o(n9948),
	.a(n22583),
	.b(FE_OFN25785_n17770),
	.c(n22677));
   na02f01 U26562 (.o(n22584),
	.a(west_input_NIB_storage_data_f_1__30_),
	.b(FE_OFN381_n17772));
   oa12f01 U26563 (.o(n8718),
	.a(n22584),
	.b(FE_OFN381_n17772),
	.c(n22747));
   oa12f01 U26564 (.o(n8708),
	.a(n22585),
	.b(FE_OFN381_n17772),
	.c(n22749));
   na02f01 U26565 (.o(n22586),
	.a(west_input_NIB_storage_data_f_1__55_),
	.b(FE_OFN381_n17772));
   na02s01 U26566 (.o(n22587),
	.a(west_input_NIB_storage_data_f_1__29_),
	.b(FE_OFN381_n17772));
   oa12s01 U26567 (.o(n8723),
	.a(n22587),
	.b(FE_OFN381_n17772),
	.c(n22739));
   na02s01 U26568 (.o(n22588),
	.a(west_input_NIB_storage_data_f_1__46_),
	.b(FE_OFN381_n17772));
   oa12f01 U26569 (.o(n8638),
	.a(n22588),
	.b(FE_OFN381_n17772),
	.c(n22743));
   na02s01 U26570 (.o(n22589),
	.a(west_input_NIB_storage_data_f_1__24_),
	.b(FE_OFN381_n17772));
   oa12s01 U26571 (.o(n8748),
	.a(n22589),
	.b(FE_OFN381_n17772),
	.c(n22736));
   na02s01 U26572 (.o(n22590),
	.a(west_input_NIB_storage_data_f_1__23_),
	.b(FE_OFN381_n17772));
   oa12s01 U26573 (.o(n8753),
	.a(n22590),
	.b(FE_OFN381_n17772),
	.c(n22745));
   na02s01 U26574 (.o(n22591),
	.a(west_input_NIB_storage_data_f_1__22_),
	.b(FE_OFN381_n17772));
   oa12s01 U26575 (.o(n8758),
	.a(n22591),
	.b(FE_OFN381_n17772),
	.c(n22732));
   na02s01 U26576 (.o(n22592),
	.a(west_input_NIB_storage_data_f_1__28_),
	.b(FE_OFN381_n17772));
   oa12s01 U26577 (.o(n8728),
	.a(n22592),
	.b(FE_OFN381_n17772),
	.c(n22712));
   na02s01 U26578 (.o(n22593),
	.a(west_input_NIB_storage_data_f_1__27_),
	.b(FE_OFN381_n17772));
   oa12s01 U26579 (.o(n8733),
	.a(n22593),
	.b(FE_OFN381_n17772),
	.c(n22728));
   na02s01 U26580 (.o(n22594),
	.a(west_input_NIB_storage_data_f_1__26_),
	.b(FE_OFN381_n17772));
   oa12s01 U26581 (.o(n8738),
	.a(n22594),
	.b(FE_OFN381_n17772),
	.c(n22751));
   na02s01 U26582 (.o(n22595),
	.a(west_input_NIB_storage_data_f_1__57_),
	.b(FE_OFN382_n17772));
   oa12s01 U26583 (.o(n8583),
	.a(n22595),
	.b(FE_OFN382_n17772),
	.c(n22741));
   na02f01 U26584 (.o(n22596),
	.a(west_input_NIB_storage_data_f_1__59_),
	.b(FE_OFN381_n17772));
   oa12f01 U26585 (.o(n8573),
	.a(n22596),
	.b(FE_OFN381_n17772),
	.c(n22734));
   na02f01 U26586 (.o(n22597),
	.a(west_input_NIB_storage_data_f_1__58_),
	.b(FE_OFN381_n17772));
   oa12f01 U26587 (.o(n8578),
	.a(n22597),
	.b(FE_OFN381_n17772),
	.c(n22730));
   ao22f01 U26588 (.o(n22599),
	.a(n19493),
	.b(n23975),
	.c(FE_OFN577_n25498),
	.d(n23974));
   ao22f01 U26589 (.o(n22598),
	.a(FE_OFN105_n22517),
	.b(n23976),
	.c(FE_OFN93_n21667),
	.d(n23977));
   ao22f01 U26591 (.o(n22603),
	.a(n19493),
	.b(n23147),
	.c(FE_OFN93_n21667),
	.d(n23146));
   ao22f01 U26592 (.o(n22602),
	.a(FE_OFN105_n22517),
	.b(n23149),
	.c(n25498),
	.d(FE_OFN116_n23148));
   na02f02 U26593 (.o(n22604),
	.a(n22603),
	.b(n22602));
   ao22f01 U26595 (.o(n22607),
	.a(FE_OFN577_n25498),
	.b(FE_OFN130_n23559),
	.c(FE_OFN93_n21667),
	.d(FE_OFN473_n23560));
   ao22f01 U26596 (.o(n22606),
	.a(n19493),
	.b(n23562),
	.c(FE_OFN105_n22517),
	.d(n23561));
   na02f02 U26597 (.o(n22608),
	.a(n22607),
	.b(n22606));
   in01s01 U26598 (.o(n22609),
	.a(n22608));
   ao22f01 U26599 (.o(n22611),
	.a(FE_OFN577_n25498),
	.b(n23568),
	.c(FE_OFN93_n21667),
	.d(n23569));
   ao22f01 U26600 (.o(n22610),
	.a(n19493),
	.b(n23571),
	.c(FE_OFN105_n22517),
	.d(n23570));
   na02f02 U26601 (.o(n22612),
	.a(n22611),
	.b(n22610));
   ao22f01 U26602 (.o(n22615),
	.a(n19493),
	.b(FE_OFN485_n24011),
	.c(FE_OFN577_n25498),
	.d(FE_OFN146_n24010));
   ao22f01 U26603 (.o(n22614),
	.a(FE_OFN105_n22517),
	.b(n24012),
	.c(FE_OFN93_n21667),
	.d(FE_OFN487_n24013));
   na02f02 U26604 (.o(n22616),
	.a(n22615),
	.b(n22614));
   ao22f01 U26606 (.o(n22619),
	.a(FE_OFN105_n22517),
	.b(n23577),
	.c(FE_OFN93_n21667),
	.d(FE_OFN477_n23578));
   ao22f01 U26607 (.o(n22618),
	.a(n19493),
	.b(n23580),
	.c(n25498),
	.d(n23579));
   na02f02 U26608 (.o(n22620),
	.a(n22619),
	.b(n22618));
   in01s01 U26609 (.o(n22621),
	.a(n22620));
   na02f01 U26610 (.o(n22624),
	.a(n22623),
	.b(n22622));
   in01s01 U26611 (.o(n22625),
	.a(n22624));
   na02s01 U26612 (.o(n22629),
	.a(north_input_NIB_storage_data_f_0__43_),
	.b(n20934));
   oa12s01 U26613 (.o(n12203),
	.a(n22629),
	.b(n20934),
	.c(n22630));
   na02s01 U26614 (.o(n22631),
	.a(north_input_NIB_storage_data_f_0__45_),
	.b(n20934));
   na02s01 U26615 (.o(n22633),
	.a(north_input_NIB_storage_data_f_0__49_),
	.b(n20934));
   oa12s01 U26616 (.o(n12173),
	.a(n22633),
	.b(n20934),
	.c(n22634));
   na02s01 U26617 (.o(n22635),
	.a(north_input_NIB_storage_data_f_0__46_),
	.b(n20934));
   oa12s01 U26618 (.o(n12188),
	.a(n22635),
	.b(n20934),
	.c(n22636));
   na02s01 U26619 (.o(n22637),
	.a(north_input_NIB_storage_data_f_0__38_),
	.b(n20934));
   oa12s01 U26620 (.o(n12228),
	.a(n22637),
	.b(n20934),
	.c(n22638));
   oa12s01 U26621 (.o(n12258),
	.a(n22639),
	.b(n20934),
	.c(n22640));
   na02s01 U26622 (.o(n22641),
	.a(north_input_NIB_storage_data_f_0__59_),
	.b(n17771));
   oa12s01 U26623 (.o(n12123),
	.a(n22641),
	.b(n17771),
	.c(n22642));
   na02s01 U26624 (.o(n22643),
	.a(north_input_NIB_storage_data_f_0__35_),
	.b(n20934));
   oa12s01 U26625 (.o(n12243),
	.a(n22643),
	.b(n20934),
	.c(n22644));
   na02s01 U26626 (.o(n22645),
	.a(north_input_NIB_storage_data_f_0__39_),
	.b(n20934));
   oa12s01 U26627 (.o(n12223),
	.a(n22645),
	.b(n20934),
	.c(n22646));
   na02s01 U26628 (.o(n22647),
	.a(north_input_NIB_storage_data_f_0__34_),
	.b(n20934));
   oa12s01 U26629 (.o(n12248),
	.a(n22647),
	.b(n20934),
	.c(n22648));
   na02s01 U26630 (.o(n22649),
	.a(north_input_NIB_storage_data_f_0__42_),
	.b(n20934));
   oa12s01 U26631 (.o(n12208),
	.a(n22649),
	.b(n20934),
	.c(n22650));
   na02s01 U26632 (.o(n22651),
	.a(north_input_NIB_storage_data_f_0__48_),
	.b(n20934));
   oa12s01 U26633 (.o(n12178),
	.a(n22651),
	.b(n20934),
	.c(n22652));
   na02s01 U26634 (.o(n22653),
	.a(north_input_NIB_storage_data_f_0__37_),
	.b(n20934));
   oa12s01 U26635 (.o(n12233),
	.a(n22653),
	.b(n20934),
	.c(n22654));
   na02s01 U26636 (.o(n22655),
	.a(north_input_NIB_storage_data_f_0__36_),
	.b(n20934));
   oa12s01 U26637 (.o(n12238),
	.a(n22655),
	.b(n20934),
	.c(n22656));
   na02s01 U26638 (.o(n22663),
	.a(south_input_NIB_storage_data_f_3__37_),
	.b(n17769));
   oa12s01 U26639 (.o(n10613),
	.a(n22663),
	.b(n22682),
	.c(n17769));
   na02s01 U26640 (.o(n22664),
	.a(south_input_NIB_storage_data_f_3__31_),
	.b(n17769));
   oa12s01 U26641 (.o(n10643),
	.a(n22664),
	.b(n22698),
	.c(n17769));
   na02s01 U26642 (.o(n22665),
	.a(south_input_NIB_storage_data_f_3__32_),
	.b(n17769));
   oa12s01 U26643 (.o(n10638),
	.a(n22665),
	.b(n22702),
	.c(n17769));
   na02s01 U26644 (.o(n22666),
	.a(south_input_NIB_storage_data_f_3__34_),
	.b(n17769));
   oa12s01 U26645 (.o(n10628),
	.a(n22666),
	.b(n22667),
	.c(n17769));
   na02s01 U26646 (.o(n22668),
	.a(south_input_NIB_storage_data_f_3__35_),
	.b(n17769));
   oa12s01 U26647 (.o(n10623),
	.a(n22668),
	.b(n22696),
	.c(n17769));
   na02s01 U26648 (.o(n22669),
	.a(south_input_NIB_storage_data_f_3__36_),
	.b(n17769));
   na02s01 U26649 (.o(n22670),
	.a(south_input_NIB_storage_data_f_3__44_),
	.b(n17769));
   oa12s01 U26650 (.o(n10578),
	.a(n22670),
	.b(n22700),
	.c(n17769));
   na02s01 U26651 (.o(n22671),
	.a(south_input_NIB_storage_data_f_3__45_),
	.b(n17769));
   oa12s01 U26652 (.o(n10573),
	.a(n22671),
	.b(n22694),
	.c(n17769));
   na02s01 U26653 (.o(n22672),
	.a(south_input_NIB_storage_data_f_3__38_),
	.b(n17769));
   oa12s01 U26654 (.o(n10608),
	.a(n22672),
	.b(n22690),
	.c(n17769));
   na02s01 U26655 (.o(n22673),
	.a(south_input_NIB_storage_data_f_3__46_),
	.b(n17769));
   oa12s01 U26656 (.o(n10568),
	.a(n22673),
	.b(n22684),
	.c(n17769));
   na02s01 U26657 (.o(n22674),
	.a(south_input_NIB_storage_data_f_3__42_),
	.b(n17769));
   oa12s01 U26658 (.o(n10588),
	.a(n22674),
	.b(n22677),
	.c(n17769));
   na02s01 U26659 (.o(n22675),
	.a(south_input_NIB_storage_data_f_3__43_),
	.b(n17769));
   oa12s01 U26660 (.o(n10583),
	.a(n22675),
	.b(n22692),
	.c(n17769));
   na02f01 U26661 (.o(n22676),
	.a(south_input_NIB_storage_data_f_2__42_),
	.b(FE_OFN84_n20972));
   oa12f01 U26662 (.o(n10268),
	.a(n22676),
	.b(FE_OFN84_n20972),
	.c(n22677));
   na02f01 U26663 (.o(n22678),
	.a(south_input_NIB_storage_data_f_2__48_),
	.b(FE_OFN84_n20972));
   na02s01 U26664 (.o(n22680),
	.a(south_input_NIB_storage_data_f_3__47_),
	.b(n17769));
   oa12s01 U26665 (.o(n10563),
	.a(n22680),
	.b(n17769),
	.c(n22704));
   na02f01 U26666 (.o(n22681),
	.a(south_input_NIB_storage_data_f_2__37_),
	.b(FE_OFN84_n20972));
   oa12f01 U26667 (.o(n10293),
	.a(n22681),
	.b(FE_OFN84_n20972),
	.c(n22682));
   na02f01 U26668 (.o(n22683),
	.a(south_input_NIB_storage_data_f_2__46_),
	.b(FE_OFN84_n20972));
   oa12f01 U26669 (.o(n10248),
	.a(n22683),
	.b(FE_OFN84_n20972),
	.c(n22684));
   na02s01 U26670 (.o(n22685),
	.a(south_input_NIB_storage_data_f_3__63_),
	.b(FE_OFN896_n17769));
   oa12s01 U26671 (.o(n10483),
	.a(n22685),
	.b(FE_OFN896_n17769),
	.c(n22686));
   na02f01 U26672 (.o(n22687),
	.a(south_input_NIB_storage_data_f_2__41_),
	.b(FE_OFN84_n20972));
   oa12f01 U26673 (.o(n10273),
	.a(n22687),
	.b(FE_OFN84_n20972),
	.c(n22688));
   na02f01 U26674 (.o(n22689),
	.a(south_input_NIB_storage_data_f_2__38_),
	.b(FE_OFN84_n20972));
   oa12f01 U26675 (.o(n10288),
	.a(n22689),
	.b(FE_OFN84_n20972),
	.c(n22690));
   na02f01 U26676 (.o(n22691),
	.a(south_input_NIB_storage_data_f_2__43_),
	.b(FE_OFN84_n20972));
   oa12f01 U26677 (.o(n10263),
	.a(n22691),
	.b(FE_OFN84_n20972),
	.c(n22692));
   na02f01 U26678 (.o(n22693),
	.a(south_input_NIB_storage_data_f_2__45_),
	.b(FE_OFN84_n20972));
   oa12f01 U26679 (.o(n10253),
	.a(n22693),
	.b(FE_OFN84_n20972),
	.c(n22694));
   na02f01 U26680 (.o(n22695),
	.a(south_input_NIB_storage_data_f_2__35_),
	.b(FE_OFN84_n20972));
   oa12f01 U26681 (.o(n10303),
	.a(n22695),
	.b(FE_OFN84_n20972),
	.c(n22696));
   na02f01 U26682 (.o(n22697),
	.a(south_input_NIB_storage_data_f_2__31_),
	.b(FE_OFN84_n20972));
   oa12f01 U26683 (.o(n10323),
	.a(n22697),
	.b(FE_OFN84_n20972),
	.c(n22698));
   na02f01 U26684 (.o(n22699),
	.a(south_input_NIB_storage_data_f_2__44_),
	.b(FE_OFN84_n20972));
   oa12f01 U26685 (.o(n10258),
	.a(n22699),
	.b(FE_OFN84_n20972),
	.c(n22700));
   na02f01 U26686 (.o(n22701),
	.a(south_input_NIB_storage_data_f_2__32_),
	.b(FE_OFN84_n20972));
   na02f01 U26687 (.o(n22703),
	.a(south_input_NIB_storage_data_f_2__47_),
	.b(FE_OFN84_n20972));
   na02f01 U26688 (.o(n22705),
	.a(south_input_NIB_storage_data_f_2__36_),
	.b(FE_OFN84_n20972));
   oa12f01 U26689 (.o(n10298),
	.a(n22705),
	.b(FE_OFN84_n20972),
	.c(n22706));
   na02f01 U26690 (.o(n22707),
	.a(west_input_NIB_storage_data_f_2__27_),
	.b(n21053));
   na02f01 U26691 (.o(n22709),
	.a(west_input_NIB_storage_data_f_2__32_),
	.b(FE_OFN25792_n21053));
   na02f01 U26692 (.o(n22710),
	.a(west_input_NIB_storage_data_f_3__28_),
	.b(FE_OFN25862_FE_OFN24766_n21069));
   na02f01 U26693 (.o(n22711),
	.a(west_input_NIB_storage_data_f_2__28_),
	.b(n21053));
   na02f01 U26694 (.o(n22713),
	.a(west_input_NIB_storage_data_f_2__31_),
	.b(FE_OFN25792_n21053));
   na02f01 U26695 (.o(n22715),
	.a(west_input_NIB_storage_data_f_2__24_),
	.b(n21053));
   na02f01 U26696 (.o(n22716),
	.a(west_input_NIB_storage_data_f_2__52_),
	.b(FE_OFN25791_n21053));
   oa12f01 U26697 (.o(n8928),
	.a(n22716),
	.b(FE_OFN25791_n21053),
	.c(n22717));
   na02f01 U26698 (.o(n22718),
	.a(west_input_NIB_storage_data_f_3__55_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U26699 (.o(n9233),
	.a(n22718),
	.b(n22724),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U26700 (.o(n22719),
	.a(west_input_NIB_storage_data_f_3__59_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U26701 (.o(n9213),
	.a(n22719),
	.b(FE_OFN25866_FE_OFN24766_n21069),
	.c(n22734));
   na02f01 U26702 (.o(n22720),
	.a(west_input_NIB_storage_data_f_2__58_),
	.b(FE_OFN25792_n21053));
   oa12f01 U26703 (.o(n8898),
	.a(n22720),
	.b(FE_OFN25792_n21053),
	.c(n22730));
   na02f01 U26704 (.o(n22721),
	.a(west_input_NIB_storage_data_f_2__22_),
	.b(FE_OFN25792_n21053));
   na02f01 U26705 (.o(n22722),
	.a(west_input_NIB_storage_data_f_3__57_),
	.b(FE_OFN24767_n21069));
   oa12f01 U26706 (.o(n9223),
	.a(n22722),
	.b(n22741),
	.c(FE_OFN24767_n21069));
   na02f01 U26707 (.o(n22723),
	.a(west_input_NIB_storage_data_f_2__55_),
	.b(FE_OFN25792_n21053));
   oa12f01 U26708 (.o(n8913),
	.a(n22723),
	.b(FE_OFN25792_n21053),
	.c(n22724));
   na02f01 U26709 (.o(n22725),
	.a(west_input_NIB_storage_data_f_2__25_),
	.b(n21053));
   na02f01 U26710 (.o(n22727),
	.a(west_input_NIB_storage_data_f_3__27_),
	.b(FE_OFN25865_FE_OFN24766_n21069));
   na02f01 U26711 (.o(n22729),
	.a(west_input_NIB_storage_data_f_3__58_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   oa12f01 U26712 (.o(n9218),
	.a(n22729),
	.b(n22730),
	.c(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U26713 (.o(n22731),
	.a(west_input_NIB_storage_data_f_3__22_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U26714 (.o(n22733),
	.a(west_input_NIB_storage_data_f_2__59_),
	.b(FE_OFN25792_n21053));
   na02s01 U26715 (.o(n22735),
	.a(west_input_NIB_storage_data_f_3__24_),
	.b(FE_OFN1098_n25937));
   na02f01 U26716 (.o(n22737),
	.a(west_input_NIB_storage_data_f_3__30_),
	.b(n25937));
   na02s01 U26717 (.o(n22738),
	.a(west_input_NIB_storage_data_f_3__29_),
	.b(FE_OFN1100_n25937));
   na02f01 U26718 (.o(n22740),
	.a(west_input_NIB_storage_data_f_2__57_),
	.b(FE_OFN25791_n21053));
   oa12f01 U26719 (.o(n8903),
	.a(n22740),
	.b(FE_OFN25791_n21053),
	.c(n22741));
   na02s01 U26720 (.o(n22742),
	.a(west_input_NIB_storage_data_f_3__46_),
	.b(n25937));
   oa12f01 U26721 (.o(n9278),
	.a(n22742),
	.b(FE_OFN25866_FE_OFN24766_n21069),
	.c(n22743));
   na02s01 U26722 (.o(n22744),
	.a(west_input_NIB_storage_data_f_3__23_),
	.b(FE_OFN1099_n25937));
   na02f01 U26723 (.o(n22746),
	.a(west_input_NIB_storage_data_f_2__30_),
	.b(FE_OFN25792_n21053));
   na02f01 U26724 (.o(n22748),
	.a(west_input_NIB_storage_data_f_3__32_),
	.b(FE_OFN25866_FE_OFN24766_n21069));
   na02f01 U26725 (.o(n22750),
	.a(west_input_NIB_storage_data_f_3__26_),
	.b(FE_OFN24766_n21069));
   in01s01 U26726 (.o(n6828),
	.a(n22780));
   in01s01 U26727 (.o(n6898),
	.a(n22781));
   in01s01 U26728 (.o(n6838),
	.a(n22782));
   in01s01 U26729 (.o(n6903),
	.a(n22783));
   in01s01 U26730 (.o(n6878),
	.a(n22784));
   in01s01 U26731 (.o(n6843),
	.a(n22785));
   in01s01 U26732 (.o(n6913),
	.a(n22786));
   in01s01 U26733 (.o(n6873),
	.a(n22787));
   in01s01 U26734 (.o(n6888),
	.a(n22788));
   in01s01 U26735 (.o(n6823),
	.a(n22789));
   in01s01 U26736 (.o(n6848),
	.a(n22790));
   in01s01 U26737 (.o(n6918),
	.a(n22791));
   in01s01 U26738 (.o(n6908),
	.a(n22792));
   in01s01 U26739 (.o(n6863),
	.a(n22794));
   in01s01 U26740 (.o(n6763),
	.a(n22795));
   in01s01 U26741 (.o(n6858),
	.a(n22796));
   in01s01 U26742 (.o(n6883),
	.a(n22797));
   in01s01 U26743 (.o(n6833),
	.a(n22798));
   in01s01 U26744 (.o(n6923),
	.a(n22799));
   in01s01 U26745 (.o(n6893),
	.a(n22800));
   in01s01 U26746 (.o(n6853),
	.a(n22801));
   in01s01 U26747 (.o(n6928),
	.a(n22802));
   no02f01 U26748 (.o(n22825),
	.a(n22824),
	.b(n22823));
   no02f01 U26749 (.o(n22833),
	.a(n22832),
	.b(n22831));
   no02f02 U26750 (.o(n22841),
	.a(n22840),
	.b(n22839));
   no02f01 U26751 (.o(n22856),
	.a(n22855),
	.b(n22854));
   no02f01 U26752 (.o(n22864),
	.a(n22863),
	.b(n22862));
   no02f01 U26753 (.o(n22872),
	.a(n22871),
	.b(n22870));
   no02f01 U26754 (.o(n22880),
	.a(n22879),
	.b(n22878));
   no02f01 U26755 (.o(n22887),
	.a(n22886),
	.b(n22885));
   oa12f01 U26756 (.o(FE_OFN833_dataOut_P_38),
	.a(n22887),
	.b(n18031),
	.c(n24728));
   no02s01 U26757 (.o(n22897),
	.a(proc_input_control_count_f_7_),
	.b(proc_input_control_count_f_6_));
   na02f01 U26758 (.o(n22905),
	.a(FE_OFN251_n25152),
	.b(n18092));
   na03f02 U26759 (.o(dataOut_W_59_),
	.a(n22907),
	.b(n22906),
	.c(n22905));
   na03f02 U26760 (.o(dataOut_W_53_),
	.a(n22910),
	.b(n22909),
	.c(n22908));
   ao22m01 U26761 (.o(n22917),
	.a(n25247),
	.b(n23958),
	.c(south_input_control_count_f_7_),
	.d(n22911));
   na02s01 U26762 (.o(n22913),
	.a(south_input_control_count_f_7_),
	.b(n22912));
   na02s01 U26763 (.o(n22914),
	.a(south_input_control_count_f_6_),
	.b(n22913));
   oa12s01 U26764 (.o(n22916),
	.a(n22914),
	.b(south_input_control_count_f_6_),
	.c(n22915));
   ao12f01 U26765 (.o(south_input_control_N48),
	.a(FE_OFN5_reset),
	.b(n22917),
	.c(n22916));
   no02f01 U26766 (.o(n22933),
	.a(n22930),
	.b(n22929));
   na02f02 U26767 (.o(dataOut_P_41_),
	.a(n22933),
	.b(n22932));
   no02f01 U26768 (.o(n22935),
	.a(FE_OFN8_reset),
	.b(n22934));
   in01s01 U26769 (.o(n22936),
	.a(north_output_space_valid_f));
   no02s01 U26770 (.o(n22937),
	.a(north_output_space_is_one_f),
	.b(north_output_space_yummy_f));
   no02s01 U26771 (.o(n22938),
	.a(n25370),
	.b(n22937));
   no02s01 U26772 (.o(n22940),
	.a(proc_output_space_is_one_f),
	.b(proc_output_space_yummy_f));
   no02s01 U26773 (.o(n22942),
	.a(n22941),
	.b(n22940));
   no03m02 U26774 (.o(proc_output_control_N72),
	.a(proc_output_space_is_two_or_more_f),
	.b(n22943),
	.c(n22942));
   na02f04 U26775 (.o(n22945),
	.a(n22957),
	.b(n22944));
   in01s01 U26776 (.o(n24927),
	.a(dataIn_E_48_));
   na02f01 U26777 (.o(n22947),
	.a(east_input_NIB_storage_data_f_0__48_),
	.b(FE_OFN433_n22945));
   oa12f01 U26778 (.o(n10888),
	.a(n22947),
	.b(n22945),
	.c(n24927));
   in01s01 U26779 (.o(n24935),
	.a(dataIn_E_49_));
   na02f01 U26780 (.o(n22948),
	.a(east_input_NIB_storage_data_f_0__49_),
	.b(FE_OFN24837_n22945));
   oa12f01 U26781 (.o(n10883),
	.a(n22948),
	.b(n22946),
	.c(n24935));
   in01s01 U26782 (.o(n25206),
	.a(dataIn_E_57_));
   na02f01 U26783 (.o(n22949),
	.a(east_input_NIB_storage_data_f_0__57_),
	.b(FE_OFN432_n22945));
   oa12f01 U26784 (.o(n10843),
	.a(n22949),
	.b(FE_OFN432_n22945),
	.c(n25206));
   in01s01 U26785 (.o(n25202),
	.a(dataIn_E_60_));
   na02f01 U26786 (.o(n22950),
	.a(east_input_NIB_storage_data_f_0__60_),
	.b(FE_OFN432_n22945));
   oa12f01 U26787 (.o(n10828),
	.a(n22950),
	.b(FE_OFN432_n22945),
	.c(n25202));
   in01s01 U26788 (.o(n25204),
	.a(dataIn_E_53_));
   na02f01 U26789 (.o(n22951),
	.a(east_input_NIB_storage_data_f_0__53_),
	.b(FE_OFN432_n22945));
   oa12f01 U26790 (.o(n10863),
	.a(n22951),
	.b(FE_OFN432_n22945),
	.c(n25204));
   in01s01 U26791 (.o(n25220),
	.a(dataIn_E_30_));
   na02f01 U26792 (.o(n22952),
	.a(east_input_NIB_storage_data_f_0__30_),
	.b(n22945));
   oa12f01 U26793 (.o(n10978),
	.a(n22952),
	.b(n22945),
	.c(n25220));
   in01s01 U26794 (.o(n24923),
	.a(dataIn_E_43_));
   na02f01 U26795 (.o(n22953),
	.a(east_input_NIB_storage_data_f_0__43_),
	.b(FE_OFN24846_n22945));
   in01s01 U26796 (.o(n24937),
	.a(dataIn_E_42_));
   na02f01 U26797 (.o(n22954),
	.a(east_input_NIB_storage_data_f_0__42_),
	.b(FE_OFN24849_n22945));
   na02s01 U26798 (.o(n22955),
	.a(validIn_E),
	.b(east_input_NIB_tail_ptr_f_1_));
   na02f10 U26799 (.o(n22958),
	.a(n22957),
	.b(n22956));
   na02f01 U26800 (.o(n22960),
	.a(east_input_NIB_storage_data_f_2__42_),
	.b(n22958));
   oa12f01 U26801 (.o(n11558),
	.a(n22960),
	.b(n24937),
	.c(n22958));
   na02f01 U26802 (.o(n22961),
	.a(east_input_NIB_storage_data_f_2__43_),
	.b(n22958));
   oa12f01 U26803 (.o(n11553),
	.a(n22961),
	.b(n22958),
	.c(n24923));
   na02f01 U26804 (.o(n22962),
	.a(east_input_NIB_storage_data_f_0__32_),
	.b(n22945));
   oa12f01 U26805 (.o(n10968),
	.a(n22962),
	.b(n22945),
	.c(n25222));
   na02f01 U26806 (.o(n22963),
	.a(east_input_NIB_storage_data_f_2__48_),
	.b(n22958));
   oa12f01 U26807 (.o(n11528),
	.a(n22963),
	.b(n24927),
	.c(n22958));
   na02f01 U26808 (.o(n22964),
	.a(east_input_NIB_storage_data_f_2__49_),
	.b(n22958));
   oa12f01 U26809 (.o(n11523),
	.a(n22964),
	.b(n24935),
	.c(n22958));
   in01s01 U26810 (.o(n25190),
	.a(dataIn_E_41_));
   na02f01 U26811 (.o(n22965),
	.a(east_input_NIB_storage_data_f_0__41_),
	.b(FE_OFN24838_n22945));
   oa12f01 U26812 (.o(n10923),
	.a(n22965),
	.b(FE_OFN24839_n22945),
	.c(n25190));
   na02f01 U26813 (.o(n22966),
	.a(east_input_NIB_storage_data_f_2__60_),
	.b(FE_OFN436_n22958));
   oa12f01 U26814 (.o(n11468),
	.a(n22966),
	.b(n25202),
	.c(FE_OFN436_n22958));
   na02f01 U26815 (.o(n22967),
	.a(east_input_NIB_storage_data_f_0__40_),
	.b(FE_OFN24840_n22945));
   oa12f01 U26816 (.o(n10928),
	.a(n22967),
	.b(FE_OFN24841_n22945),
	.c(n24931));
   na02f01 U26817 (.o(n22968),
	.a(east_input_NIB_storage_data_f_2__32_),
	.b(n22958));
   oa12f01 U26818 (.o(n11608),
	.a(n22968),
	.b(n25222),
	.c(n22958));
   na02f01 U26819 (.o(n22969),
	.a(east_input_NIB_storage_data_f_2__53_),
	.b(FE_OFN436_n22958));
   oa12f01 U26820 (.o(n11503),
	.a(n22969),
	.b(n25204),
	.c(FE_OFN436_n22958));
   in01s01 U26821 (.o(n24933),
	.a(dataIn_E_39_));
   na02f01 U26822 (.o(n22970),
	.a(east_input_NIB_storage_data_f_0__39_),
	.b(FE_OFN24844_n22945));
   oa12f01 U26823 (.o(n10933),
	.a(n22970),
	.b(FE_OFN24845_n22945),
	.c(n24933));
   in01s01 U26824 (.o(n25210),
	.a(dataIn_E_54_));
   na02f01 U26825 (.o(n22971),
	.a(east_input_NIB_storage_data_f_2__54_),
	.b(FE_OFN436_n22958));
   oa12f01 U26826 (.o(n11498),
	.a(n22971),
	.b(n25210),
	.c(FE_OFN436_n22958));
   in01s01 U26827 (.o(n24929),
	.a(dataIn_E_38_));
   na02f01 U26828 (.o(n22972),
	.a(east_input_NIB_storage_data_f_0__38_),
	.b(FE_OFN24843_n22945));
   oa12f01 U26829 (.o(n10938),
	.a(n22972),
	.b(FE_OFN24842_n22945),
	.c(n24929));
   na02f01 U26830 (.o(n22973),
	.a(east_input_NIB_storage_data_f_2__57_),
	.b(FE_OFN436_n22958));
   oa12f01 U26831 (.o(n11483),
	.a(n22973),
	.b(n25206),
	.c(FE_OFN436_n22958));
   na02f01 U26832 (.o(n22974),
	.a(east_input_NIB_storage_data_f_2__38_),
	.b(n22958));
   oa12f01 U26833 (.o(n11578),
	.a(n22974),
	.b(n24929),
	.c(n22958));
   na02f01 U26834 (.o(n22975),
	.a(east_input_NIB_storage_data_f_2__41_),
	.b(n22958));
   oa12f01 U26835 (.o(n11563),
	.a(n22975),
	.b(n22958),
	.c(n25190));
   oa12f01 U26836 (.o(n11568),
	.a(n22976),
	.b(n24931),
	.c(n22958));
   in01s01 U26837 (.o(n25218),
	.a(dataIn_E_62_));
   na02f01 U26838 (.o(n22977),
	.a(east_input_NIB_storage_data_f_2__62_),
	.b(FE_OFN436_n22958));
   oa12f01 U26839 (.o(n11458),
	.a(n22977),
	.b(n25218),
	.c(FE_OFN436_n22958));
   in01s01 U26840 (.o(n24925),
	.a(dataIn_E_34_));
   na02f01 U26841 (.o(n22978),
	.a(east_input_NIB_storage_data_f_2__34_),
	.b(n22958));
   oa12f01 U26842 (.o(n11598),
	.a(n22978),
	.b(n24925),
	.c(n22958));
   na02f01 U26843 (.o(n22979),
	.a(east_input_NIB_storage_data_f_2__39_),
	.b(n22958));
   oa12f01 U26844 (.o(n11573),
	.a(n22979),
	.b(n24933),
	.c(n22958));
   na02f01 U26845 (.o(n22980),
	.a(east_input_NIB_storage_data_f_2__30_),
	.b(n22958));
   oa12f01 U26846 (.o(n11618),
	.a(n22980),
	.b(n25220),
	.c(n22958));
   in01s01 U26847 (.o(n25257),
	.a(dataIn_E_26_));
   na02f01 U26848 (.o(n22981),
	.a(east_input_NIB_storage_data_f_0__26_),
	.b(FE_OFN24856_n22945));
   in01s01 U26849 (.o(n25212),
	.a(dataIn_E_50_));
   na02f01 U26850 (.o(n22982),
	.a(east_input_NIB_storage_data_f_2__50_),
	.b(FE_OFN436_n22958));
   oa12f01 U26851 (.o(n11518),
	.a(n22982),
	.b(FE_OFN436_n22958),
	.c(n25212));
   in01s01 U26852 (.o(n25208),
	.a(dataIn_E_61_));
   na02f01 U26853 (.o(n22983),
	.a(east_input_NIB_storage_data_f_2__61_),
	.b(FE_OFN436_n22958));
   oa12f01 U26854 (.o(n11463),
	.a(n22983),
	.b(n25208),
	.c(FE_OFN436_n22958));
   in01s01 U26855 (.o(n25194),
	.a(dataIn_E_58_));
   na02f01 U26856 (.o(n22984),
	.a(east_input_NIB_storage_data_f_2__58_),
	.b(FE_OFN436_n22958));
   oa12f01 U26857 (.o(n11478),
	.a(n22984),
	.b(n25194),
	.c(FE_OFN436_n22958));
   in01s01 U26858 (.o(n24941),
	.a(dataIn_E_37_));
   na02f01 U26859 (.o(n22985),
	.a(east_input_NIB_storage_data_f_2__37_),
	.b(n22958));
   oa12f01 U26860 (.o(n11583),
	.a(n22985),
	.b(n24941),
	.c(n22958));
   in01s01 U26861 (.o(n24939),
	.a(dataIn_E_35_));
   na02f01 U26862 (.o(n22986),
	.a(east_input_NIB_storage_data_f_2__35_),
	.b(n22958));
   in01s01 U26863 (.o(n25198),
	.a(dataIn_E_63_));
   na02f01 U26864 (.o(n22987),
	.a(east_input_NIB_storage_data_f_2__63_),
	.b(FE_OFN436_n22958));
   oa12f01 U26865 (.o(n11453),
	.a(n22987),
	.b(FE_OFN436_n22958),
	.c(n25198));
   in01s01 U26866 (.o(n25200),
	.a(dataIn_E_52_));
   na02f01 U26867 (.o(n22988),
	.a(east_input_NIB_storage_data_f_2__52_),
	.b(FE_OFN436_n22958));
   oa12f01 U26868 (.o(n11508),
	.a(n22988),
	.b(n25200),
	.c(FE_OFN436_n22958));
   in01s01 U26869 (.o(n24943),
	.a(dataIn_E_36_));
   na02f01 U26870 (.o(n22989),
	.a(east_input_NIB_storage_data_f_2__36_),
	.b(n22958));
   in01s01 U26871 (.o(n25224),
	.a(dataIn_E_31_));
   na02f01 U26872 (.o(n22990),
	.a(east_input_NIB_storage_data_f_2__31_),
	.b(n22958));
   oa12f01 U26873 (.o(n11613),
	.a(n22990),
	.b(n22958),
	.c(n25224));
   in01s01 U26874 (.o(n24947),
	.a(dataIn_E_44_));
   na02f01 U26875 (.o(n22991),
	.a(east_input_NIB_storage_data_f_2__44_),
	.b(n22958));
   oa12f01 U26876 (.o(n11548),
	.a(n22991),
	.b(n24947),
	.c(n22958));
   in01s01 U26877 (.o(n25259),
	.a(dataIn_E_29_));
   na02f01 U26878 (.o(n22992),
	.a(east_input_NIB_storage_data_f_2__29_),
	.b(n22958));
   oa12f01 U26879 (.o(n11623),
	.a(n22992),
	.b(n22958),
	.c(n25259));
   in01s01 U26880 (.o(n25267),
	.a(dataIn_E_28_));
   na02f01 U26881 (.o(n22993),
	.a(east_input_NIB_storage_data_f_2__28_),
	.b(n22958));
   oa12f01 U26882 (.o(n11628),
	.a(n22993),
	.b(n25267),
	.c(n22958));
   in01s01 U26883 (.o(n25265),
	.a(dataIn_E_27_));
   na02f01 U26884 (.o(n22994),
	.a(east_input_NIB_storage_data_f_2__27_),
	.b(FE_OFN436_n22958));
   oa12f01 U26885 (.o(n11633),
	.a(n22994),
	.b(n25265),
	.c(FE_OFN436_n22958));
   na02f01 U26886 (.o(n22995),
	.a(east_input_NIB_storage_data_f_2__26_),
	.b(n22958));
   in01s01 U26887 (.o(n25263),
	.a(dataIn_E_25_));
   in01s01 U26888 (.o(n25261),
	.a(dataIn_E_24_));
   na02f01 U26889 (.o(n22997),
	.a(east_input_NIB_storage_data_f_2__24_),
	.b(n22958));
   na02f01 U26890 (.o(n22998),
	.a(east_input_NIB_storage_data_f_0__62_),
	.b(FE_OFN432_n22945));
   oa12f01 U26891 (.o(n10818),
	.a(n22998),
	.b(FE_OFN432_n22945),
	.c(n25218));
   oa12f01 U26892 (.o(n10823),
	.a(n22999),
	.b(FE_OFN432_n22945),
	.c(n25208));
   in01s01 U26893 (.o(n25255),
	.a(dataIn_E_23_));
   na02f01 U26894 (.o(n23000),
	.a(east_input_NIB_storage_data_f_2__23_),
	.b(n22958));
   na02f01 U26895 (.o(n23001),
	.a(east_input_NIB_storage_data_f_0__58_),
	.b(FE_OFN432_n22945));
   oa12f01 U26896 (.o(n10838),
	.a(n23001),
	.b(FE_OFN432_n22945),
	.c(n25194));
   in01s01 U26897 (.o(n25253),
	.a(dataIn_E_22_));
   na02f01 U26898 (.o(n23002),
	.a(east_input_NIB_storage_data_f_2__22_),
	.b(n22958));
   na02f01 U26899 (.o(n23003),
	.a(east_input_NIB_storage_data_f_0__63_),
	.b(FE_OFN432_n22945));
   oa12f01 U26900 (.o(n10813),
	.a(n23003),
	.b(n25198),
	.c(FE_OFN432_n22945));
   in01s01 U26901 (.o(n24945),
	.a(dataIn_E_45_));
   na02f01 U26902 (.o(n23004),
	.a(east_input_NIB_storage_data_f_0__45_),
	.b(FE_OFN24861_n22945));
   oa12f01 U26903 (.o(n10903),
	.a(n23004),
	.b(FE_OFN24861_n22945),
	.c(n24945));
   in01s01 U26904 (.o(n25214),
	.a(dataIn_E_51_));
   na02f01 U26905 (.o(n23005),
	.a(east_input_NIB_storage_data_f_0__51_),
	.b(FE_OFN432_n22945));
   oa12f01 U26906 (.o(n10873),
	.a(n23005),
	.b(FE_OFN432_n22945),
	.c(n25214));
   na02f01 U26907 (.o(n23006),
	.a(east_input_NIB_storage_data_f_0__50_),
	.b(FE_OFN432_n22945));
   oa12f01 U26908 (.o(n10878),
	.a(n23006),
	.b(n25212),
	.c(FE_OFN432_n22945));
   na02f01 U26909 (.o(n23007),
	.a(east_input_NIB_storage_data_f_0__36_),
	.b(FE_OFN24850_n22945));
   oa12f01 U26910 (.o(n10948),
	.a(n23007),
	.b(FE_OFN24850_n22945),
	.c(n24943));
   oa12f01 U26911 (.o(n10973),
	.a(n23008),
	.b(n25224),
	.c(FE_OFN24844_n22945));
   na02f01 U26912 (.o(n23009),
	.a(east_input_NIB_storage_data_f_0__37_),
	.b(FE_OFN24844_n22945));
   oa12f01 U26913 (.o(n10943),
	.a(n23009),
	.b(FE_OFN24844_n22945),
	.c(n24941));
   na02f01 U26914 (.o(n23010),
	.a(east_input_NIB_storage_data_f_0__44_),
	.b(FE_OFN24858_n22945));
   oa12f01 U26915 (.o(n10908),
	.a(n23010),
	.b(FE_OFN24859_n22945),
	.c(n24947));
   na02f01 U26916 (.o(n23011),
	.a(east_input_NIB_storage_data_f_0__25_),
	.b(FE_OFN24860_n22945));
   na02f01 U26917 (.o(n23012),
	.a(east_input_NIB_storage_data_f_0__35_),
	.b(FE_OFN24844_n22945));
   oa12f01 U26918 (.o(n10953),
	.a(n23012),
	.b(n24939),
	.c(FE_OFN24844_n22945));
   na02f01 U26919 (.o(n23013),
	.a(east_input_NIB_storage_data_f_0__34_),
	.b(FE_OFN24854_n22945));
   oa12f01 U26920 (.o(n10958),
	.a(n23013),
	.b(FE_OFN24853_n22945),
	.c(n24925));
   na02f01 U26921 (.o(n23014),
	.a(east_input_NIB_storage_data_f_0__22_),
	.b(FE_OFN24844_n22945));
   na02f01 U26922 (.o(n23015),
	.a(east_input_NIB_storage_data_f_0__23_),
	.b(FE_OFN24844_n22945));
   na02f01 U26923 (.o(n23016),
	.a(east_input_NIB_storage_data_f_0__24_),
	.b(FE_OFN24844_n22945));
   in01s01 U26924 (.o(n24949),
	.a(dataIn_E_47_));
   na02f01 U26925 (.o(n23017),
	.a(east_input_NIB_storage_data_f_0__47_),
	.b(FE_OFN24855_n22945));
   oa12f01 U26926 (.o(n10893),
	.a(n23017),
	.b(FE_OFN24855_n22945),
	.c(n24949));
   na02f01 U26927 (.o(n23018),
	.a(east_input_NIB_storage_data_f_0__28_),
	.b(FE_OFN24844_n22945));
   oa12f01 U26928 (.o(n10988),
	.a(n23018),
	.b(FE_OFN24844_n22945),
	.c(n25267));
   na02f01 U26929 (.o(n23019),
	.a(east_input_NIB_storage_data_f_0__29_),
	.b(FE_OFN24844_n22945));
   oa12f01 U26930 (.o(n10983),
	.a(n23019),
	.b(n25259),
	.c(FE_OFN24844_n22945));
   in01s01 U26931 (.o(n24951),
	.a(dataIn_E_46_));
   oa12f01 U26932 (.o(n10898),
	.a(n23020),
	.b(FE_OFN24852_n22945),
	.c(n24951));
   na02f01 U26933 (.o(n23021),
	.a(east_input_NIB_storage_data_f_0__27_),
	.b(FE_OFN432_n22945));
   oa12f01 U26934 (.o(n10993),
	.a(n23021),
	.b(FE_OFN432_n22945),
	.c(n25265));
   oa12f01 U26935 (.o(n11493),
	.a(n23022),
	.b(n25196),
	.c(FE_OFN436_n22958));
   na02f01 U26936 (.o(n23023),
	.a(east_input_NIB_storage_data_f_0__55_),
	.b(FE_OFN432_n22945));
   oa12f01 U26937 (.o(n10853),
	.a(n23023),
	.b(FE_OFN432_n22945),
	.c(n25196));
   na02f01 U26938 (.o(n23024),
	.a(east_input_NIB_storage_data_f_2__51_),
	.b(FE_OFN436_n22958));
   oa12f01 U26939 (.o(n11513),
	.a(n23024),
	.b(n25214),
	.c(FE_OFN436_n22958));
   in01s01 U26940 (.o(n25192),
	.a(dataIn_E_59_));
   na02f01 U26941 (.o(n23025),
	.a(east_input_NIB_storage_data_f_2__59_),
	.b(FE_OFN436_n22958));
   oa12f01 U26942 (.o(n11473),
	.a(n23025),
	.b(n25192),
	.c(FE_OFN436_n22958));
   na02f01 U26943 (.o(n23026),
	.a(east_input_NIB_storage_data_f_2__47_),
	.b(n22958));
   oa12f01 U26944 (.o(n11533),
	.a(n23026),
	.b(n24949),
	.c(n22958));
   na02f01 U26945 (.o(n23027),
	.a(east_input_NIB_storage_data_f_0__52_),
	.b(FE_OFN432_n22945));
   oa12f01 U26946 (.o(n10868),
	.a(n23027),
	.b(FE_OFN432_n22945),
	.c(n25200));
   na02f01 U26947 (.o(n23028),
	.a(east_input_NIB_storage_data_f_2__46_),
	.b(n22958));
   oa12f01 U26948 (.o(n11538),
	.a(n23028),
	.b(n24951),
	.c(n22958));
   na02f01 U26949 (.o(n23029),
	.a(east_input_NIB_storage_data_f_0__59_),
	.b(FE_OFN432_n22945));
   oa12f01 U26950 (.o(n10833),
	.a(n23029),
	.b(FE_OFN432_n22945),
	.c(n25192));
   in01s01 U26951 (.o(n25216),
	.a(dataIn_E_56_));
   na02f01 U26952 (.o(n23030),
	.a(east_input_NIB_storage_data_f_2__56_),
	.b(FE_OFN436_n22958));
   oa12f01 U26953 (.o(n11488),
	.a(n23030),
	.b(n25216),
	.c(FE_OFN436_n22958));
   na02f01 U26954 (.o(n23031),
	.a(east_input_NIB_storage_data_f_0__56_),
	.b(FE_OFN432_n22945));
   oa12f01 U26955 (.o(n10848),
	.a(n23031),
	.b(FE_OFN432_n22945),
	.c(n25216));
   na02f01 U26956 (.o(n23032),
	.a(east_input_NIB_storage_data_f_0__54_),
	.b(FE_OFN432_n22945));
   oa12f01 U26957 (.o(n10858),
	.a(n23032),
	.b(FE_OFN432_n22945),
	.c(n25210));
   na02f01 U26958 (.o(n23033),
	.a(east_input_NIB_storage_data_f_2__45_),
	.b(n22958));
   oa12f01 U26959 (.o(n11543),
	.a(n23033),
	.b(n24945),
	.c(n22958));
   in01s01 U26960 (.o(n23040),
	.a(n25227));
   in01s01 U26961 (.o(n25225),
	.a(west_input_control_count_f_6_));
   na02s01 U26962 (.o(n23042),
	.a(n23041),
	.b(n24970));
   ao12f01 U26963 (.o(west_input_control_N47),
	.a(FE_OFN25647_reset),
	.b(n23043),
	.c(n23042));
   in01s01 U26964 (.o(n5613),
	.a(n23047));
   in01s01 U26965 (.o(n5598),
	.a(n23048));
   in01s01 U26966 (.o(n5623),
	.a(n23049));
   in01s01 U26967 (.o(n5323),
	.a(n23052));
   in01s01 U26968 (.o(n5583),
	.a(n23053));
   in01s01 U26970 (.o(n5608),
	.a(n23055));
   in01s01 U26971 (.o(n5303),
	.a(n23057));
   in01s01 U26972 (.o(n5603),
	.a(n23058));
   in01s01 U26973 (.o(n5588),
	.a(n23059));
   in01s01 U26974 (.o(n5288),
	.a(n23060));
   in01s01 U26975 (.o(n5628),
	.a(n23061));
   in01s01 U26976 (.o(n5633),
	.a(n23062));
   in01s01 U26977 (.o(n5313),
	.a(n23063));
   in01s01 U26978 (.o(n5643),
	.a(n23064));
   in01s01 U26979 (.o(n5268),
	.a(n23065));
   in01s01 U26980 (.o(n5578),
	.a(n23066));
   in01s01 U26981 (.o(n5573),
	.a(n23067));
   in01s01 U26982 (.o(n5568),
	.a(n23069));
   in01s01 U26983 (.o(n5563),
	.a(n23070));
   in01s01 U26984 (.o(n5283),
	.a(n23071));
   in01s01 U26985 (.o(n5278),
	.a(n23072));
   in01s01 U26986 (.o(n5273),
	.a(n23073));
   in01s01 U26987 (.o(n5553),
	.a(n23074));
   in01s01 U26988 (.o(n5248),
	.a(n23075));
   in01s01 U26989 (.o(n5328),
	.a(n23076));
   in01s01 U26990 (.o(n5548),
	.a(n23077));
   in01s01 U26991 (.o(n5638),
	.a(n23078));
   in01s01 U26992 (.o(n5558),
	.a(n23079));
   in01s01 U26993 (.o(n5648),
	.a(n23080));
   in01s01 U26994 (.o(n5263),
	.a(n23081));
   in01s01 U26995 (.o(n5318),
	.a(n23082));
   in01s01 U26996 (.o(n5543),
	.a(n23083));
   in01s01 U26997 (.o(n5258),
	.a(n23084));
   in01s01 U26998 (.o(n5308),
	.a(n23085));
   in01s01 U26999 (.o(n5253),
	.a(n23086));
   in01s01 U27000 (.o(n5298),
	.a(n23087));
   in01s01 U27001 (.o(n5243),
	.a(n23088));
   oa22m01 U27002 (.o(n23091),
	.a(FE_OFN25766_FE_OFN1077_n17766),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_4__33_),
	.d(n23090));
   in01s01 U27003 (.o(n4523),
	.a(n23091));
   in01s01 U27004 (.o(n5238),
	.a(n23092));
   in01s01 U27005 (.o(n5233),
	.a(n23093));
   in01s01 U27006 (.o(n5228),
	.a(n23094));
   in01s01 U27007 (.o(n5223),
	.a(n23095));
   in01s01 U27008 (.o(n5163),
	.a(n23096));
   oa22m01 U27009 (.o(n23097),
	.a(FE_OFN25763_FE_OFN1077_n17766),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_4__21_),
	.d(n23090));
   in01s01 U27010 (.o(n4583),
	.a(n23097));
   oa22m01 U27011 (.o(n23098),
	.a(FE_OFN25761_FE_OFN1077_n17766),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_4__20_),
	.d(n23090));
   in01s01 U27012 (.o(n4588),
	.a(n23098));
   oa22m01 U27013 (.o(n23099),
	.a(FE_OFN1077_n17766),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_4__19_),
	.d(n23090));
   in01s01 U27014 (.o(n4593),
	.a(n23099));
   in01s01 U27015 (.o(n5008),
	.a(n23103));
   oa22m01 U27016 (.o(n23104),
	.a(FE_OFN1077_n17766),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_4__18_),
	.d(n23090));
   in01s01 U27017 (.o(n4598),
	.a(n23104));
   in01s01 U27018 (.o(n5003),
	.a(n23105));
   in01s01 U27019 (.o(n4998),
	.a(n23106));
   in01s01 U27020 (.o(n4988),
	.a(n23108));
   in01s01 U27021 (.o(n4983),
	.a(n23109));
   in01s01 U27022 (.o(n4978),
	.a(n23110));
   in01s01 U27023 (.o(n4973),
	.a(n23111));
   in01s01 U27024 (.o(n4968),
	.a(n23112));
   in01s01 U27025 (.o(n4963),
	.a(n23113));
   oa22m01 U27026 (.o(n23114),
	.a(FE_OFN1077_n17766),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_4__17_),
	.d(n23090));
   in01s01 U27027 (.o(n4603),
	.a(n23114));
   in01s01 U27028 (.o(n4958),
	.a(n23115));
   oa22m01 U27029 (.o(n23116),
	.a(FE_OFN25763_FE_OFN1077_n17766),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_4__16_),
	.d(n23090));
   in01s01 U27030 (.o(n4608),
	.a(n23116));
   in01s01 U27031 (.o(n4953),
	.a(n23117));
   in01s01 U27032 (.o(n4948),
	.a(n23118));
   oa22m01 U27033 (.o(n23119),
	.a(FE_OFN25761_FE_OFN1077_n17766),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_4__15_),
	.d(n23090));
   in01s01 U27034 (.o(n4613),
	.a(n23119));
   in01s01 U27035 (.o(n4943),
	.a(n23120));
   in01s01 U27036 (.o(n4938),
	.a(n23122));
   in01s01 U27037 (.o(n4623),
	.a(n23123));
   in01s01 U27038 (.o(n4933),
	.a(n23124));
   in01s01 U27039 (.o(n4928),
	.a(n23125));
   in01s01 U27040 (.o(n4923),
	.a(n23126));
   oa22m01 U27041 (.o(n23128),
	.a(FE_OFN25761_FE_OFN1077_n17766),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_4__5_),
	.d(n23090));
   in01s01 U27042 (.o(n4663),
	.a(n23128));
   oa22m01 U27043 (.o(n23129),
	.a(FE_OFN1077_n17766),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_4__12_),
	.d(n23090));
   in01s01 U27044 (.o(n4628),
	.a(n23129));
   in01s01 U27046 (.o(n4908),
	.a(n23131));
   in01s01 U27047 (.o(n4903),
	.a(n23132));
   oa22m01 U27048 (.o(n23134),
	.a(FE_OFN1077_n17766),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_4__11_),
	.d(n23090));
   in01s01 U27049 (.o(n4633),
	.a(n23134));
   in01s01 U27050 (.o(n4688),
	.a(n23135));
   oa22m01 U27051 (.o(n23136),
	.a(FE_OFN25761_FE_OFN1077_n17766),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_4__10_),
	.d(n23090));
   in01s01 U27052 (.o(n4638),
	.a(n23136));
   oa22m01 U27053 (.o(n23137),
	.a(FE_OFN1077_n17766),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_4__9_),
	.d(n23090));
   in01s01 U27054 (.o(n4643),
	.a(n23137));
   oa22m01 U27055 (.o(n23138),
	.a(FE_OFN1077_n17766),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_4__4_),
	.d(n23090));
   in01s01 U27056 (.o(n4668),
	.a(n23138));
   oa22m01 U27057 (.o(n23139),
	.a(FE_OFN1077_n17766),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_4__8_),
	.d(n23090));
   in01s01 U27058 (.o(n4648),
	.a(n23139));
   oa22m01 U27059 (.o(n23140),
	.a(FE_OFN25762_FE_OFN1077_n17766),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_4__7_),
	.d(n23090));
   in01s01 U27060 (.o(n4653),
	.a(n23140));
   oa22m01 U27061 (.o(n23141),
	.a(FE_OFN1077_n17766),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_4__6_),
	.d(n23090));
   in01s01 U27062 (.o(n4658),
	.a(n23141));
   in01s01 U27063 (.o(n5483),
	.a(n23142));
   oa22m01 U27064 (.o(n23143),
	.a(FE_OFN25762_FE_OFN1077_n17766),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_4__3_),
	.d(n23090));
   in01s01 U27065 (.o(n4673),
	.a(n23143));
   in01s01 U27066 (.o(n4683),
	.a(n23144));
   in01s01 U27067 (.o(n4678),
	.a(n23145));
   ao22f01 U27068 (.o(n23151),
	.a(n25295),
	.b(n23147),
	.c(n25294),
	.d(n23146));
   na02f02 U27069 (.o(n23152),
	.a(n23151),
	.b(n23150));
   in01s01 U27070 (.o(n23153),
	.a(n23152));
   na02f01 U27071 (.o(n23155),
	.a(proc_input_NIB_storage_data_f_6__38_),
	.b(FE_OFN25801_n23051));
   na02s01 U27072 (.o(n23156),
	.a(proc_input_NIB_storage_data_f_5__41_),
	.b(FE_OFN369_n17761));
   na02s01 U27073 (.o(n23157),
	.a(proc_input_NIB_storage_data_f_7__38_),
	.b(n17767));
   na02s01 U27074 (.o(n23158),
	.a(proc_input_NIB_storage_data_f_7__35_),
	.b(n17767));
   na02f01 U27075 (.o(n23159),
	.a(proc_input_NIB_storage_data_f_4__37_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02f01 U27076 (.o(n23160),
	.a(proc_input_NIB_storage_data_f_5__44_),
	.b(FE_OFN368_n17761));
   na02f01 U27077 (.o(n23161),
	.a(proc_input_NIB_storage_data_f_4__42_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27078 (.o(n23162),
	.a(proc_input_NIB_storage_data_f_7__34_),
	.b(n17767));
   na02s01 U27079 (.o(n23163),
	.a(proc_input_NIB_storage_data_f_7__31_),
	.b(FE_OFN1081_n17767));
   na02s01 U27080 (.o(n23164),
	.a(proc_input_NIB_storage_data_f_7__30_),
	.b(n17767));
   na02s01 U27081 (.o(n23166),
	.a(proc_input_NIB_storage_data_f_4__47_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27082 (.o(n23168),
	.a(proc_input_NIB_storage_data_f_5__43_),
	.b(FE_OFN369_n17761));
   na02s01 U27083 (.o(n23169),
	.a(proc_input_NIB_storage_data_f_7__39_),
	.b(FE_OFN1081_n17767));
   na02f01 U27084 (.o(n23170),
	.a(proc_input_NIB_storage_data_f_6__30_),
	.b(FE_OFN25806_n23051));
   na02f01 U27085 (.o(n23171),
	.a(proc_input_NIB_storage_data_f_5__40_),
	.b(FE_OFN368_n17761));
   na02f01 U27086 (.o(n23172),
	.a(proc_input_NIB_storage_data_f_4__43_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27087 (.o(n23173),
	.a(proc_input_NIB_storage_data_f_5__42_),
	.b(FE_OFN369_n17761));
   na02f01 U27088 (.o(n23174),
	.a(proc_input_NIB_storage_data_f_6__35_),
	.b(FE_OFN25801_n23051));
   na02f01 U27089 (.o(n23175),
	.a(proc_input_NIB_storage_data_f_6__34_),
	.b(FE_OFN25801_n23051));
   na02s01 U27090 (.o(n23176),
	.a(proc_input_NIB_storage_data_f_4__40_),
	.b(FE_OFN1077_n17766));
   na02s01 U27091 (.o(n23177),
	.a(proc_input_NIB_storage_data_f_4__44_),
	.b(FE_OFN25767_FE_OFN1077_n17766));
   na02f01 U27092 (.o(n23178),
	.a(proc_input_NIB_storage_data_f_5__45_),
	.b(FE_OFN368_n17761));
   na02s01 U27093 (.o(n23179),
	.a(proc_input_NIB_storage_data_f_6__39_),
	.b(FE_OFN25801_n23051));
   na02s01 U27094 (.o(n23180),
	.a(proc_input_NIB_storage_data_f_4__45_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27095 (.o(n23181),
	.a(proc_input_NIB_storage_data_f_6__31_),
	.b(FE_OFN25798_n23051));
   na02s01 U27096 (.o(n23182),
	.a(proc_input_NIB_storage_data_f_5__37_),
	.b(FE_OFN369_n17761));
   no02f01 U27097 (.o(n23191),
	.a(n23188),
	.b(n23187));
   na02f01 U27098 (.o(FE_OFN364_dataOut_P_40),
	.a(n23191),
	.b(n23190));
   oa22f01 U27099 (.o(n23192),
	.a(FE_OFN25628_n21910),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_12__17_),
	.d(FE_OFN912_n23246));
   in01s01 U27100 (.o(n7163),
	.a(n23192));
   in01s01 U27101 (.o(n7178),
	.a(n23193));
   oa22f01 U27102 (.o(n23194),
	.a(FE_OFN913_n23246),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_12__20_),
	.d(n23246));
   in01s01 U27103 (.o(n7148),
	.a(n23194));
   oa22f01 U27104 (.o(n23195),
	.a(FE_OFN25626_n21910),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_12__10_),
	.d(FE_OFN912_n23246));
   in01s01 U27105 (.o(n7198),
	.a(n23195));
   oa22f01 U27106 (.o(n23196),
	.a(FE_OFN25628_n21910),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_12__21_),
	.d(FE_OFN912_n23246));
   in01s01 U27107 (.o(n7143),
	.a(n23196));
   oa22f01 U27108 (.o(n23197),
	.a(FE_OFN25626_n21910),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_12__13_),
	.d(FE_OFN912_n23246));
   in01s01 U27109 (.o(n7183),
	.a(n23197));
   in01s01 U27110 (.o(n7223),
	.a(n23198));
   oa22f01 U27111 (.o(n23199),
	.a(FE_OFN25629_n21910),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_12__19_),
	.d(FE_OFN912_n23246));
   in01s01 U27112 (.o(n7153),
	.a(n23199));
   oa22f01 U27113 (.o(n23200),
	.a(FE_OFN25627_n21910),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_12__12_),
	.d(FE_OFN912_n23246));
   in01s01 U27114 (.o(n7188),
	.a(n23200));
   in01s01 U27115 (.o(n7233),
	.a(n23201));
   in01s01 U27116 (.o(n7228),
	.a(n23202));
   oa22f01 U27117 (.o(n23203),
	.a(FE_OFN25628_n21910),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_12__7_),
	.d(FE_OFN912_n23246));
   in01s01 U27118 (.o(n7213),
	.a(n23203));
   in01s01 U27119 (.o(n7173),
	.a(n23204));
   in01s01 U27120 (.o(n7403),
	.a(n23206));
   in01s01 U27121 (.o(n7463),
	.a(n23207));
   oa22f01 U27122 (.o(n23209),
	.a(FE_OFN25629_n21910),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_12__9_),
	.d(FE_OFN912_n23246));
   in01s01 U27123 (.o(n7203),
	.a(n23209));
   in01s01 U27124 (.o(n7238),
	.a(n23210));
   in01s01 U27125 (.o(n7218),
	.a(n23211));
   oa22f01 U27126 (.o(n23212),
	.a(FE_OFN448_n23236),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_13__16_),
	.d(n21915));
   in01s01 U27127 (.o(n7488),
	.a(n23212));
   oa22f01 U27128 (.o(n23213),
	.a(n23236),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_13__15_),
	.d(n21915));
   in01s01 U27129 (.o(n7493),
	.a(n23213));
   oa22f01 U27130 (.o(n23214),
	.a(FE_OFN448_n23236),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_13__14_),
	.d(n21915));
   in01s01 U27131 (.o(n7498),
	.a(n23214));
   oa22f01 U27132 (.o(n23215),
	.a(FE_OFN25627_n21910),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_12__11_),
	.d(FE_OFN912_n23246));
   in01s01 U27133 (.o(n7193),
	.a(n23215));
   oa22f01 U27134 (.o(n23216),
	.a(FE_OFN25627_n21910),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_12__18_),
	.d(FE_OFN912_n23246));
   in01s01 U27135 (.o(n7158),
	.a(n23216));
   oa22f01 U27136 (.o(n23217),
	.a(n23236),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_13__13_),
	.d(n21915));
   in01s01 U27137 (.o(n7503),
	.a(n23217));
   oa22f01 U27138 (.o(n23218),
	.a(FE_OFN448_n23236),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_13__12_),
	.d(n21915));
   in01s01 U27139 (.o(n7508),
	.a(n23218));
   oa22f01 U27140 (.o(n23219),
	.a(FE_OFN448_n23236),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_13__11_),
	.d(n21915));
   in01s01 U27141 (.o(n7513),
	.a(n23219));
   in01s01 U27142 (.o(n7248),
	.a(n23221));
   oa22f01 U27143 (.o(n23222),
	.a(n23236),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_13__10_),
	.d(n21915));
   in01s01 U27144 (.o(n7518),
	.a(n23222));
   oa22f01 U27145 (.o(n23223),
	.a(n23236),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_13__9_),
	.d(n21915));
   in01s01 U27146 (.o(n7523),
	.a(n23223));
   oa22f01 U27147 (.o(n23224),
	.a(n23236),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_13__8_),
	.d(n21915));
   in01s01 U27148 (.o(n7528),
	.a(n23224));
   in01s01 U27149 (.o(n7473),
	.a(n23225));
   oa22f01 U27150 (.o(n23226),
	.a(FE_OFN448_n23236),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_13__18_),
	.d(n21915));
   in01s01 U27151 (.o(n7478),
	.a(n23226));
   oa22f01 U27152 (.o(n23227),
	.a(n23236),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_13__17_),
	.d(n21915));
   in01s01 U27153 (.o(n7483),
	.a(n23227));
   oa22f01 U27154 (.o(n23228),
	.a(FE_OFN448_n23236),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_13__7_),
	.d(n21915));
   in01s01 U27155 (.o(n7533),
	.a(n23228));
   in01s01 U27156 (.o(n7538),
	.a(n23229));
   oa22f01 U27157 (.o(n23231),
	.a(FE_OFN25629_n21910),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_12__8_),
	.d(FE_OFN912_n23246));
   in01s01 U27158 (.o(n7208),
	.a(n23231));
   in01s01 U27159 (.o(n7548),
	.a(n23232));
   in01s01 U27160 (.o(n7553),
	.a(n23233));
   in01s01 U27161 (.o(n7558),
	.a(n23234));
   in01s01 U27162 (.o(n7563),
	.a(n23235));
   in01s01 U27163 (.o(n7568),
	.a(n23237));
   oa22f01 U27164 (.o(n23238),
	.a(FE_OFN25605_n21944),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_14__33_),
	.d(n23262));
   in01s01 U27165 (.o(n7723),
	.a(n23238));
   oa22f01 U27166 (.o(n23239),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_14__21_),
	.d(n21945));
   in01s01 U27167 (.o(n7783),
	.a(n23239));
   oa22f01 U27168 (.o(n23240),
	.a(FE_OFN25605_n21944),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_14__20_),
	.d(n23262));
   in01s01 U27169 (.o(n7788),
	.a(n23240));
   oa22f01 U27170 (.o(n23241),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_14__19_),
	.d(n21945));
   in01s01 U27171 (.o(n7793),
	.a(n23241));
   oa22f01 U27172 (.o(n23242),
	.a(FE_OFN25605_n21944),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_14__18_),
	.d(n23262));
   in01s01 U27173 (.o(n7798),
	.a(n23242));
   oa22f01 U27174 (.o(n23243),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_14__17_),
	.d(n21945));
   in01s01 U27175 (.o(n7803),
	.a(n23243));
   oa22f01 U27176 (.o(n23244),
	.a(FE_OFN25739_FE_OFN25605_n21944),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_14__15_),
	.d(n21945));
   in01s01 U27177 (.o(n7813),
	.a(n23244));
   oa22f01 U27178 (.o(n23245),
	.a(FE_OFN25605_n21944),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_14__16_),
	.d(n23262));
   in01s01 U27179 (.o(n7808),
	.a(n23245));
   oa22f01 U27180 (.o(n23247),
	.a(FE_OFN25626_n21910),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_12__33_),
	.d(FE_OFN912_n23246));
   in01s01 U27181 (.o(n7083),
	.a(n23247));
   in01s01 U27182 (.o(n7888),
	.a(n23248));
   oa22f01 U27183 (.o(n23249),
	.a(FE_OFN25605_n21944),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_14__14_),
	.d(n23262));
   in01s01 U27184 (.o(n7818),
	.a(n23249));
   oa22f01 U27185 (.o(n23250),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_14__13_),
	.d(n21945));
   in01s01 U27186 (.o(n7823),
	.a(n23250));
   oa22f01 U27187 (.o(n23251),
	.a(FE_OFN25605_n21944),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_14__12_),
	.d(n23262));
   in01s01 U27188 (.o(n7828),
	.a(n23251));
   in01s01 U27189 (.o(n7833),
	.a(n23252));
   oa22f01 U27191 (.o(n23255),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_14__8_),
	.d(n21945));
   in01s01 U27192 (.o(n7848),
	.a(n23255));
   oa22f01 U27193 (.o(n23256),
	.a(FE_OFN453_n23262),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_14__7_),
	.d(n21945));
   in01s01 U27194 (.o(n7853),
	.a(n23256));
   in01s01 U27195 (.o(n7858),
	.a(n23257));
   in01s01 U27196 (.o(n7863),
	.a(n23258));
   in01s01 U27197 (.o(n7868),
	.a(n23259));
   in01s01 U27198 (.o(n7873),
	.a(n23260));
   in01s01 U27199 (.o(n7878),
	.a(n23261));
   in01s01 U27200 (.o(n7883),
	.a(n23263));
   ao12s01 U27201 (.o(n23310),
	.a(n23308),
	.b(south_input_control_count_f_4_),
	.c(n23309));
   no02s01 U27202 (.o(n23314),
	.a(n23310),
	.b(n25250));
   in01f01 U27203 (.o(n23313),
	.a(n23311));
   in01s01 U27204 (.o(n25240),
	.a(south_input_control_count_f_4_));
   no02s01 U27205 (.o(n23312),
	.a(n23550),
	.b(n25240));
   no02f01 U27206 (.o(south_input_control_N45),
	.a(FE_OFN5_reset),
	.b(n23315));
   na02f01 U27207 (.o(n23348),
	.a(FE_OFN262_n25301),
	.b(n18092));
   na02s01 U27208 (.o(n23351),
	.a(proc_input_NIB_storage_data_f_4__35_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27209 (.o(n23352),
	.a(proc_input_NIB_storage_data_f_4__36_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02f02 U27210 (.o(n23353),
	.a(proc_input_NIB_storage_data_f_5__39_),
	.b(FE_OFN368_n17761));
   na02s01 U27211 (.o(n23354),
	.a(proc_input_NIB_storage_data_f_4__30_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27212 (.o(n23355),
	.a(proc_input_NIB_storage_data_f_4__38_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27213 (.o(n23356),
	.a(proc_input_NIB_storage_data_f_5__38_),
	.b(FE_OFN369_n17761));
   na02s01 U27214 (.o(n23357),
	.a(proc_input_NIB_storage_data_f_4__31_),
	.b(FE_OFN25765_FE_OFN1077_n17766));
   na02s01 U27215 (.o(n23358),
	.a(proc_input_NIB_storage_data_f_6__42_),
	.b(FE_OFN25798_n23051));
   na02s01 U27216 (.o(n23359),
	.a(proc_input_NIB_storage_data_f_4__34_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02f01 U27217 (.o(n23360),
	.a(proc_input_NIB_storage_data_f_6__37_),
	.b(FE_OFN25802_n23051));
   na02s01 U27218 (.o(n23361),
	.a(proc_input_NIB_storage_data_f_6__45_),
	.b(FE_OFN25798_n23051));
   na02s01 U27219 (.o(n23363),
	.a(proc_input_NIB_storage_data_f_5__35_),
	.b(FE_OFN369_n17761));
   na02s01 U27220 (.o(n23364),
	.a(proc_input_NIB_storage_data_f_5__34_),
	.b(FE_OFN369_n17761));
   na02f01 U27221 (.o(n23365),
	.a(proc_input_NIB_storage_data_f_6__47_),
	.b(FE_OFN25801_n23051));
   na02f01 U27222 (.o(n23366),
	.a(proc_input_NIB_storage_data_f_5__31_),
	.b(FE_OFN368_n17761));
   na02s01 U27223 (.o(n23367),
	.a(proc_input_NIB_storage_data_f_5__30_),
	.b(FE_OFN369_n17761));
   na02s01 U27224 (.o(n23368),
	.a(proc_input_NIB_storage_data_f_6__44_),
	.b(FE_OFN25798_n23051));
   na02f01 U27225 (.o(n23369),
	.a(proc_input_NIB_storage_data_f_6__41_),
	.b(FE_OFN25802_n23051));
   na02f01 U27226 (.o(n23370),
	.a(proc_input_NIB_storage_data_f_6__43_),
	.b(FE_OFN25801_n23051));
   na02s01 U27227 (.o(n23371),
	.a(proc_input_NIB_storage_data_f_7__47_),
	.b(n17767));
   na02s01 U27228 (.o(n23372),
	.a(proc_input_NIB_storage_data_f_7__37_),
	.b(n17767));
   na02s01 U27229 (.o(n23373),
	.a(proc_input_NIB_storage_data_f_7__45_),
	.b(FE_OFN1081_n17767));
   na02s01 U27230 (.o(n23374),
	.a(proc_input_NIB_storage_data_f_7__41_),
	.b(n17767));
   na02s01 U27231 (.o(n23375),
	.a(proc_input_NIB_storage_data_f_7__44_),
	.b(FE_OFN1081_n17767));
   na02s01 U27232 (.o(n23376),
	.a(proc_input_NIB_storage_data_f_7__43_),
	.b(n17767));
   na02s01 U27233 (.o(n23377),
	.a(proc_input_NIB_storage_data_f_7__42_),
	.b(n17767));
   na02s01 U27234 (.o(n23378),
	.a(proc_input_NIB_storage_data_f_7__40_),
	.b(FE_OFN1081_n17767));
   na02s01 U27235 (.o(n23393),
	.a(proc_input_NIB_storage_data_f_11__61_),
	.b(n22923));
   na02s01 U27236 (.o(n23394),
	.a(proc_input_NIB_storage_data_f_11__62_),
	.b(n22923));
   na02s01 U27237 (.o(n23395),
	.a(proc_input_NIB_storage_data_f_11__54_),
	.b(n22923));
   na02s01 U27238 (.o(n23396),
	.a(proc_input_NIB_storage_data_f_11__59_),
	.b(n22923));
   na02s01 U27239 (.o(n23399),
	.a(n23398),
	.b(n23397));
   no02f02 U27240 (.o(east_output_control_N72),
	.a(n23400),
	.b(n23399));
   oa22f01 U27241 (.o(n23406),
	.a(n23453),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_10__13_),
	.d(n22140));
   in01s01 U27242 (.o(n6543),
	.a(n23406));
   oa22f01 U27243 (.o(n23407),
	.a(FE_OFN103_n22140),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_10__14_),
	.d(FE_OFN104_n22140));
   in01s01 U27244 (.o(n6538),
	.a(n23407));
   oa22f01 U27245 (.o(n23408),
	.a(FE_OFN103_n22140),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_10__16_),
	.d(FE_OFN104_n22140));
   in01s01 U27246 (.o(n6528),
	.a(n23408));
   oa22f01 U27247 (.o(n23409),
	.a(n23453),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_10__10_),
	.d(n22140));
   in01s01 U27248 (.o(n6558),
	.a(n23409));
   oa22f01 U27249 (.o(n23410),
	.a(n23453),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_10__9_),
	.d(n22140));
   in01s01 U27250 (.o(n6563),
	.a(n23410));
   oa22f01 U27251 (.o(n23411),
	.a(FE_OFN103_n22140),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_10__12_),
	.d(FE_OFN104_n22140));
   in01s01 U27252 (.o(n6548),
	.a(n23411));
   oa22f01 U27253 (.o(n23412),
	.a(FE_OFN103_n22140),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_10__20_),
	.d(FE_OFN104_n22140));
   in01s01 U27254 (.o(n6508),
	.a(n23412));
   oa22f01 U27255 (.o(n23413),
	.a(FE_OFN103_n22140),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_10__21_),
	.d(FE_OFN104_n22140));
   in01s01 U27256 (.o(n6503),
	.a(n23413));
   oa22f01 U27257 (.o(n23414),
	.a(n23453),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_10__15_),
	.d(n22140));
   in01s01 U27258 (.o(n6533),
	.a(n23414));
   in01s01 U27259 (.o(n6593),
	.a(n23415));
   oa22f01 U27260 (.o(n23416),
	.a(n23453),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_10__17_),
	.d(n22140));
   in01s01 U27261 (.o(n6523),
	.a(n23416));
   in01s01 U27262 (.o(n6288),
	.a(n23417));
   in01s01 U27263 (.o(n6283),
	.a(n23418));
   oa22f01 U27264 (.o(n23419),
	.a(FE_OFN103_n22140),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_10__11_),
	.d(FE_OFN104_n22140));
   in01s01 U27265 (.o(n6553),
	.a(n23419));
   in01s01 U27266 (.o(n6273),
	.a(n23420));
   in01s01 U27267 (.o(n6598),
	.a(n23422));
   in01s01 U27268 (.o(n6263),
	.a(n23423));
   in01s01 U27269 (.o(n6603),
	.a(n23424));
   in01s01 U27270 (.o(n6608),
	.a(n23425));
   in01s01 U27271 (.o(n6518),
	.a(n23426));
   in01s01 U27272 (.o(n6513),
	.a(n23427));
   in01s01 U27273 (.o(n6258),
	.a(n23428));
   oa22f01 U27274 (.o(n23429),
	.a(FE_OFN465_n23476),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_9__7_),
	.d(n22098));
   in01s01 U27275 (.o(n6253),
	.a(n23429));
   in01s01 U27276 (.o(n6588),
	.a(n23430));
   oa22f01 U27277 (.o(n23431),
	.a(FE_OFN101_n22098),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_9__8_),
	.d(n22098));
   in01s01 U27278 (.o(n6248),
	.a(n23431));
   oa22f01 U27279 (.o(n23432),
	.a(FE_OFN465_n23476),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_9__9_),
	.d(n22098));
   in01s01 U27280 (.o(n6243),
	.a(n23432));
   oa22f01 U27281 (.o(n23433),
	.a(FE_OFN101_n22098),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_9__10_),
	.d(n22098));
   in01s01 U27282 (.o(n6238),
	.a(n23433));
   in01s01 U27283 (.o(n6583),
	.a(n23434));
   in01s01 U27284 (.o(n6278),
	.a(n23435));
   oa22f01 U27285 (.o(n23436),
	.a(n23453),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_10__7_),
	.d(n22140));
   in01s01 U27286 (.o(n6573),
	.a(n23436));
   oa22f01 U27287 (.o(n23437),
	.a(n23453),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_10__8_),
	.d(n22140));
   oa22f01 U27288 (.o(n23438),
	.a(FE_OFN101_n22098),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_9__15_),
	.d(n22098));
   in01s01 U27289 (.o(n6213),
	.a(n23438));
   oa22f01 U27290 (.o(n23439),
	.a(FE_OFN465_n23476),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_9__16_),
	.d(n22098));
   in01s01 U27291 (.o(n6208),
	.a(n23439));
   oa22f01 U27292 (.o(n23440),
	.a(FE_OFN101_n22098),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_9__17_),
	.d(n22098));
   in01s01 U27293 (.o(n6203),
	.a(n23440));
   oa22f01 U27294 (.o(n23441),
	.a(FE_OFN465_n23476),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_9__18_),
	.d(n22098));
   in01s01 U27295 (.o(n6198),
	.a(n23441));
   oa22f01 U27296 (.o(n23442),
	.a(FE_OFN101_n22098),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_9__19_),
	.d(n22098));
   oa22f01 U27297 (.o(n23443),
	.a(FE_OFN465_n23476),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_9__20_),
	.d(n22098));
   in01s01 U27298 (.o(n6188),
	.a(n23443));
   oa22f01 U27299 (.o(n23444),
	.a(FE_OFN465_n23476),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_9__21_),
	.d(n22098));
   in01s01 U27300 (.o(n6183),
	.a(n23444));
   oa22f01 U27301 (.o(n23445),
	.a(FE_OFN101_n22098),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_9__33_),
	.d(n22098));
   in01s01 U27302 (.o(n6123),
	.a(n23445));
   in01s01 U27303 (.o(n5963),
	.a(n23447));
   in01s01 U27304 (.o(n5958),
	.a(n23448));
   in01s01 U27305 (.o(n5953),
	.a(n23449));
   in01s01 U27306 (.o(n5948),
	.a(n23450));
   in01s01 U27307 (.o(n6578),
	.a(n23451));
   in01s01 U27308 (.o(n5938),
	.a(n23452));
   oa22f01 U27309 (.o(n23454),
	.a(FE_OFN103_n22140),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_10__33_),
	.d(FE_OFN104_n22140));
   in01s01 U27310 (.o(n6443),
	.a(n23454));
   oa22f01 U27311 (.o(n23455),
	.a(n23471),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_8__7_),
	.d(FE_OFN416_n22085));
   in01s01 U27312 (.o(n5933),
	.a(n23455));
   in01s01 U27313 (.o(n5928),
	.a(n23456));
   in01s01 U27314 (.o(n5923),
	.a(n23457));
   oa22f01 U27315 (.o(n23458),
	.a(n22085),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_8__10_),
	.d(FE_OFN416_n22085));
   in01s01 U27316 (.o(n5918),
	.a(n23458));
   oa22f01 U27317 (.o(n23459),
	.a(n23471),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_8__11_),
	.d(FE_OFN416_n22085));
   in01s01 U27318 (.o(n5913),
	.a(n23459));
   oa22f01 U27319 (.o(n23460),
	.a(n23471),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_8__12_),
	.d(FE_OFN416_n22085));
   in01s01 U27320 (.o(n5908),
	.a(n23460));
   oa22f01 U27321 (.o(n23461),
	.a(n22085),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_8__13_),
	.d(FE_OFN416_n22085));
   in01s01 U27322 (.o(n5903),
	.a(n23461));
   oa22f01 U27323 (.o(n23462),
	.a(n22085),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_8__14_),
	.d(FE_OFN416_n22085));
   in01s01 U27324 (.o(n5898),
	.a(n23462));
   oa22f01 U27325 (.o(n23463),
	.a(n22085),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_8__15_),
	.d(FE_OFN416_n22085));
   oa22f01 U27326 (.o(n23464),
	.a(n23471),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_8__16_),
	.d(FE_OFN416_n22085));
   in01s01 U27327 (.o(n5888),
	.a(n23464));
   oa22f01 U27328 (.o(n23465),
	.a(n23471),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_8__17_),
	.d(FE_OFN416_n22085));
   in01s01 U27329 (.o(n5883),
	.a(n23465));
   oa22f01 U27330 (.o(n23466),
	.a(n23471),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_8__18_),
	.d(FE_OFN416_n22085));
   in01s01 U27331 (.o(n5878),
	.a(n23466));
   oa22f01 U27332 (.o(n23467),
	.a(n23471),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_8__19_),
	.d(FE_OFN416_n22085));
   in01s01 U27333 (.o(n5873),
	.a(n23467));
   in01s01 U27334 (.o(n5943),
	.a(n23468));
   oa22f01 U27335 (.o(n23469),
	.a(n22085),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_8__20_),
	.d(FE_OFN416_n22085));
   in01s01 U27336 (.o(n5868),
	.a(n23469));
   oa22f01 U27337 (.o(n23470),
	.a(n23471),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_8__21_),
	.d(FE_OFN416_n22085));
   in01s01 U27338 (.o(n5863),
	.a(n23470));
   oa22f01 U27339 (.o(n23472),
	.a(n23471),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_8__33_),
	.d(FE_OFN416_n22085));
   in01s01 U27340 (.o(n5803),
	.a(n23472));
   oa22f01 U27341 (.o(n23473),
	.a(FE_OFN465_n23476),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_9__11_),
	.d(n22098));
   in01s01 U27342 (.o(n6233),
	.a(n23473));
   oa22f01 U27343 (.o(n23474),
	.a(FE_OFN465_n23476),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_9__12_),
	.d(n22098));
   in01s01 U27344 (.o(n6228),
	.a(n23474));
   in01s01 U27345 (.o(n6223),
	.a(n23475));
   in01s01 U27346 (.o(n6218),
	.a(n23477));
   ao22f01 U27347 (.o(n23491),
	.a(FE_OFN259_n25295),
	.b(n23487),
	.c(FE_OFN79_n20501),
	.d(n23486));
   ao22f01 U27348 (.o(n23523),
	.a(FE_OFN259_n25295),
	.b(n23517),
	.c(n25294),
	.d(n23516));
   ao22f01 U27349 (.o(n23522),
	.a(FE_OFN79_n20501),
	.b(n23519),
	.c(n17787),
	.d(n23518));
   ao22f01 U27350 (.o(n23530),
	.a(FE_OFN79_n20501),
	.b(n23527),
	.c(n17787),
	.d(n23526));
   ao22f01 U27351 (.o(n23538),
	.a(n25294),
	.b(n23535),
	.c(FE_OFN79_n20501),
	.d(n23534));
   no02f01 U27353 (.o(n23547),
	.a(n23546),
	.b(n23545));
   in01f01 U27354 (.o(proc_output_space_N46),
	.a(n23549));
   no02f01 U27355 (.o(proc_input_control_N53),
	.a(reset),
	.b(n25026));
   in01s01 U27356 (.o(n25245),
	.a(n23550));
   ao22f01 U27357 (.o(n23557),
	.a(n25247),
	.b(n23950),
	.c(n25245),
	.d(south_input_control_count_f_6_));
   in01s01 U27358 (.o(n23555),
	.a(n25250));
   in01s01 U27359 (.o(n23552),
	.a(n23553));
   in01s01 U27360 (.o(n23551),
	.a(south_input_control_count_f_6_));
   in01s01 U27361 (.o(n23554),
	.a(n25237));
   na02s01 U27362 (.o(n23556),
	.a(n23555),
	.b(n23554));
   ao12f01 U27363 (.o(south_input_control_N47),
	.a(FE_OFN5_reset),
	.b(n23557),
	.c(n23556));
   ao22f01 U27365 (.o(n23563),
	.a(n25295),
	.b(n23562),
	.c(n17787),
	.d(n23561));
   na02f02 U27366 (.o(n23565),
	.a(n23564),
	.b(n23563));
   in01s01 U27367 (.o(n23566),
	.a(n23565));
   ao22f01 U27368 (.o(n23572),
	.a(n25295),
	.b(n23571),
	.c(n17787),
	.d(n23570));
   na02f02 U27369 (.o(n23574),
	.a(n23573),
	.b(n23572));
   in01f01 U27370 (.o(n23575),
	.a(n23574));
   ao22f01 U27371 (.o(n23582),
	.a(n25294),
	.b(FE_OFN477_n23578),
	.c(n17787),
	.d(n23577));
   na02f02 U27372 (.o(n23583),
	.a(n23582),
	.b(n23581));
   in01s01 U27373 (.o(n23584),
	.a(n23583));
   in01s01 U27374 (.o(n23592),
	.a(n23588));
   na02s01 U27375 (.o(n23595),
	.a(proc_input_NIB_storage_data_f_4__57_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02s01 U27376 (.o(n23596),
	.a(proc_input_NIB_storage_data_f_4__32_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27377 (.o(n23597),
	.a(proc_input_NIB_storage_data_f_4__50_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02s01 U27378 (.o(n23598),
	.a(proc_input_NIB_storage_data_f_7__50_),
	.b(FE_OFN1081_n17767));
   na02s01 U27379 (.o(n23599),
	.a(proc_input_NIB_storage_data_f_7__51_),
	.b(n17767));
   na02s01 U27380 (.o(n23600),
	.a(proc_input_NIB_storage_data_f_7__32_),
	.b(n17767));
   na02s01 U27381 (.o(n23601),
	.a(proc_input_NIB_storage_data_f_7__57_),
	.b(FE_OFN1081_n17767));
   na02f01 U27382 (.o(n23602),
	.a(proc_input_NIB_storage_data_f_4__49_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02m01 U27383 (.o(n23603),
	.a(proc_input_NIB_storage_data_f_6__32_),
	.b(FE_OFN25802_n23051));
   na02m01 U27384 (.o(n23604),
	.a(proc_input_NIB_storage_data_f_6__50_),
	.b(FE_OFN442_n23051));
   na02m01 U27385 (.o(n23605),
	.a(proc_input_NIB_storage_data_f_6__51_),
	.b(FE_OFN442_n23051));
   na02s01 U27386 (.o(n23606),
	.a(proc_input_NIB_storage_data_f_5__50_),
	.b(FE_OFN368_n17761));
   na02s01 U27387 (.o(n23607),
	.a(proc_input_NIB_storage_data_f_5__49_),
	.b(FE_OFN369_n17761));
   na02f01 U27388 (.o(n23608),
	.a(proc_input_NIB_storage_data_f_5__57_),
	.b(FE_OFN368_n17761));
   na02s01 U27389 (.o(n23609),
	.a(proc_input_NIB_storage_data_f_5__32_),
	.b(FE_OFN369_n17761));
   na02m01 U27390 (.o(n23610),
	.a(proc_input_NIB_storage_data_f_6__57_),
	.b(FE_OFN442_n23051));
   na02f01 U27391 (.o(n23617),
	.a(n23616),
	.b(n23615));
   in01s01 U27392 (.o(n23618),
	.a(n23617));
   na02f02 U27393 (.o(n23626),
	.a(n23625),
	.b(n23624));
   in01s01 U27394 (.o(n23627),
	.a(n23626));
   ao22f01 U27395 (.o(n23633),
	.a(FE_OFN25_n17787),
	.b(n23632),
	.c(n25294),
	.d(FE_OFN479_n23631));
   in01s01 U27396 (.o(n23636),
	.a(n23635));
   na02s01 U27397 (.o(n23639),
	.a(proc_input_NIB_storage_data_f_4__25_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27398 (.o(n23641),
	.a(proc_input_NIB_storage_data_f_4__27_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27399 (.o(n23642),
	.a(proc_input_NIB_storage_data_f_4__22_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27400 (.o(n23643),
	.a(proc_input_NIB_storage_data_f_5__59_),
	.b(FE_OFN368_n17761));
   na02f01 U27401 (.o(n23644),
	.a(proc_input_NIB_storage_data_f_4__24_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27402 (.o(n23645),
	.a(proc_input_NIB_storage_data_f_5__60_),
	.b(FE_OFN368_n17761));
   na02s01 U27403 (.o(n23646),
	.a(proc_input_NIB_storage_data_f_5__54_),
	.b(FE_OFN368_n17761));
   na02s01 U27404 (.o(n23647),
	.a(proc_input_NIB_storage_data_f_5__63_),
	.b(FE_OFN368_n17761));
   na02s01 U27405 (.o(n23649),
	.a(proc_input_NIB_storage_data_f_5__61_),
	.b(FE_OFN368_n17761));
   na02s01 U27406 (.o(n23650),
	.a(proc_input_NIB_storage_data_f_5__52_),
	.b(FE_OFN368_n17761));
   na02f01 U27407 (.o(n23651),
	.a(proc_input_NIB_storage_data_f_4__28_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27408 (.o(n23652),
	.a(proc_input_NIB_storage_data_f_5__48_),
	.b(FE_OFN369_n17761));
   na02s01 U27409 (.o(n23653),
	.a(proc_input_NIB_storage_data_f_5__46_),
	.b(FE_OFN369_n17761));
   na02s01 U27410 (.o(n23654),
	.a(proc_input_NIB_storage_data_f_4__63_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02s01 U27411 (.o(n23655),
	.a(proc_input_NIB_storage_data_f_4__62_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02s01 U27412 (.o(n23656),
	.a(proc_input_NIB_storage_data_f_4__61_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02s01 U27413 (.o(n23657),
	.a(proc_input_NIB_storage_data_f_4__23_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27414 (.o(n23658),
	.a(proc_input_NIB_storage_data_f_5__29_),
	.b(FE_OFN369_n17761));
   na02s01 U27415 (.o(n23659),
	.a(proc_input_NIB_storage_data_f_4__60_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02s01 U27416 (.o(n23660),
	.a(proc_input_NIB_storage_data_f_4__59_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02f01 U27417 (.o(n23661),
	.a(proc_input_NIB_storage_data_f_5__28_),
	.b(FE_OFN368_n17761));
   na02s01 U27418 (.o(n23662),
	.a(proc_input_NIB_storage_data_f_4__56_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02s01 U27419 (.o(n23663),
	.a(proc_input_NIB_storage_data_f_4__54_),
	.b(FE_OFN25765_FE_OFN1077_n17766));
   na02f01 U27420 (.o(n23664),
	.a(proc_input_NIB_storage_data_f_5__27_),
	.b(FE_OFN368_n17761));
   na02s01 U27421 (.o(n23665),
	.a(proc_input_NIB_storage_data_f_5__56_),
	.b(FE_OFN368_n17761));
   na02s01 U27422 (.o(n23666),
	.a(proc_input_NIB_storage_data_f_4__52_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02s01 U27423 (.o(n23667),
	.a(proc_input_NIB_storage_data_f_5__26_),
	.b(FE_OFN369_n17761));
   na02s01 U27424 (.o(n23668),
	.a(proc_input_NIB_storage_data_f_5__25_),
	.b(FE_OFN369_n17761));
   na02f01 U27425 (.o(n23669),
	.a(proc_input_NIB_storage_data_f_4__29_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02f01 U27426 (.o(n23670),
	.a(proc_input_NIB_storage_data_f_4__46_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27427 (.o(n23671),
	.a(proc_input_NIB_storage_data_f_7__22_),
	.b(n17767));
   na02s01 U27428 (.o(n23672),
	.a(proc_input_NIB_storage_data_f_5__24_),
	.b(FE_OFN369_n17761));
   na02s01 U27429 (.o(n23673),
	.a(proc_input_NIB_storage_data_f_7__23_),
	.b(n17767));
   na02s01 U27430 (.o(n23674),
	.a(proc_input_NIB_storage_data_f_7__24_),
	.b(n17767));
   na02s01 U27431 (.o(n23675),
	.a(proc_input_NIB_storage_data_f_7__25_),
	.b(n17767));
   na02s01 U27432 (.o(n23676),
	.a(proc_input_NIB_storage_data_f_7__26_),
	.b(n17767));
   na02f02 U27433 (.o(n23677),
	.a(proc_input_NIB_storage_data_f_4__48_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02s01 U27434 (.o(n23678),
	.a(proc_input_NIB_storage_data_f_7__27_),
	.b(FE_OFN1081_n17767));
   na02s01 U27435 (.o(n23679),
	.a(proc_input_NIB_storage_data_f_7__28_),
	.b(FE_OFN1081_n17767));
   na02s01 U27436 (.o(n23680),
	.a(proc_input_NIB_storage_data_f_5__23_),
	.b(FE_OFN369_n17761));
   na02s01 U27437 (.o(n23681),
	.a(proc_input_NIB_storage_data_f_7__29_),
	.b(n17767));
   na02s01 U27438 (.o(n23683),
	.a(proc_input_NIB_storage_data_f_5__22_),
	.b(FE_OFN369_n17761));
   na02s01 U27439 (.o(n23687),
	.a(proc_input_NIB_storage_data_f_7__63_),
	.b(FE_OFN1081_n17767));
   na02s01 U27440 (.o(n23689),
	.a(proc_input_NIB_storage_data_f_7__48_),
	.b(n17767));
   na02s01 U27441 (.o(n23690),
	.a(proc_input_NIB_storage_data_f_7__49_),
	.b(n17767));
   na02s01 U27442 (.o(n23695),
	.a(proc_input_NIB_storage_data_f_7__60_),
	.b(n17767));
   na02s01 U27443 (.o(n23697),
	.a(proc_input_NIB_storage_data_f_7__53_),
	.b(FE_OFN1081_n17767));
   na02s01 U27444 (.o(n23699),
	.a(proc_input_NIB_storage_data_f_7__55_),
	.b(FE_OFN1081_n17767));
   na02s01 U27445 (.o(n23700),
	.a(proc_input_NIB_storage_data_f_7__56_),
	.b(FE_OFN1081_n17767));
   na02s01 U27446 (.o(n23703),
	.a(proc_input_NIB_storage_data_f_7__58_),
	.b(n17767));
   na02s01 U27447 (.o(n23708),
	.a(proc_input_NIB_storage_data_f_7__62_),
	.b(n17767));
   no02f01 U27448 (.o(south_output_control_N72),
	.a(n18443),
	.b(n23712));
   na02s01 U27449 (.o(n23713),
	.a(proc_input_NIB_storage_data_f_5__58_),
	.b(FE_OFN368_n17761));
   na02s01 U27450 (.o(n23714),
	.a(proc_input_NIB_storage_data_f_5__55_),
	.b(FE_OFN368_n17761));
   na02s01 U27451 (.o(n23715),
	.a(proc_input_NIB_storage_data_f_4__39_),
	.b(FE_OFN25768_FE_OFN1077_n17766));
   na02m01 U27452 (.o(n23716),
	.a(proc_input_NIB_storage_data_f_6__46_),
	.b(FE_OFN25806_n23051));
   na02m01 U27453 (.o(n23717),
	.a(proc_input_NIB_storage_data_f_6__36_),
	.b(FE_OFN25801_n23051));
   na02m01 U27454 (.o(n23718),
	.a(proc_input_NIB_storage_data_f_6__52_),
	.b(FE_OFN442_n23051));
   na02s01 U27455 (.o(n23719),
	.a(proc_input_NIB_storage_data_f_5__51_),
	.b(FE_OFN368_n17761));
   na02m01 U27456 (.o(n23720),
	.a(proc_input_NIB_storage_data_f_6__59_),
	.b(FE_OFN442_n23051));
   na02f01 U27457 (.o(n23721),
	.a(proc_input_NIB_storage_data_f_5__53_),
	.b(FE_OFN368_n17761));
   na02m01 U27458 (.o(n23722),
	.a(proc_input_NIB_storage_data_f_6__54_),
	.b(FE_OFN442_n23051));
   na02s01 U27459 (.o(n23724),
	.a(proc_input_NIB_storage_data_f_4__53_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02s01 U27460 (.o(n23725),
	.a(proc_input_NIB_storage_data_f_4__51_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02s01 U27461 (.o(n23726),
	.a(proc_input_NIB_storage_data_f_4__58_),
	.b(FE_OFN25763_FE_OFN1077_n17766));
   na02f01 U27462 (.o(n23727),
	.a(proc_input_NIB_storage_data_f_5__36_),
	.b(FE_OFN368_n17761));
   na02s01 U27463 (.o(n23729),
	.a(proc_input_NIB_storage_data_f_7__52_),
	.b(FE_OFN1081_n17767));
   na02s01 U27464 (.o(n23730),
	.a(proc_input_NIB_storage_data_f_7__59_),
	.b(FE_OFN1081_n17767));
   na02s01 U27465 (.o(n23731),
	.a(proc_input_NIB_storage_data_f_7__54_),
	.b(FE_OFN1081_n17767));
   na02s01 U27466 (.o(n23732),
	.a(proc_input_NIB_storage_data_f_7__36_),
	.b(FE_OFN1081_n17767));
   na02m01 U27467 (.o(n23762),
	.a(proc_input_NIB_storage_data_f_1__22_),
	.b(FE_OFN373_n17762));
   oa12m01 U27468 (.o(n3618),
	.a(n23762),
	.b(FE_OFN373_n17762),
	.c(n23820));
   oa12m01 U27469 (.o(n3613),
	.a(n23763),
	.b(FE_OFN373_n17762),
	.c(n23793));
   na02m01 U27470 (.o(n23764),
	.a(proc_input_NIB_storage_data_f_1__24_),
	.b(FE_OFN373_n17762));
   oa12m01 U27471 (.o(n3608),
	.a(n23764),
	.b(FE_OFN373_n17762),
	.c(n23798));
   na02m01 U27472 (.o(n23765),
	.a(proc_input_NIB_storage_data_f_1__25_),
	.b(FE_OFN373_n17762));
   oa12m01 U27473 (.o(n3603),
	.a(n23765),
	.b(FE_OFN373_n17762),
	.c(n23802));
   na02m01 U27474 (.o(n23766),
	.a(proc_input_NIB_storage_data_f_1__26_),
	.b(FE_OFN373_n17762));
   oa12m01 U27475 (.o(n3598),
	.a(n23766),
	.b(FE_OFN373_n17762),
	.c(n23818));
   na02m01 U27476 (.o(n23767),
	.a(proc_input_NIB_storage_data_f_1__27_),
	.b(FE_OFN373_n17762));
   oa12m01 U27477 (.o(n3593),
	.a(n23767),
	.b(FE_OFN373_n17762),
	.c(n23822));
   na02m01 U27478 (.o(n23768),
	.a(proc_input_NIB_storage_data_f_1__28_),
	.b(FE_OFN373_n17762));
   oa12m01 U27479 (.o(n3588),
	.a(n23768),
	.b(FE_OFN373_n17762),
	.c(n23814));
   na02m01 U27480 (.o(n23769),
	.a(proc_input_NIB_storage_data_f_1__29_),
	.b(FE_OFN373_n17762));
   oa12m01 U27481 (.o(n3583),
	.a(n23769),
	.b(FE_OFN373_n17762),
	.c(n23804));
   na02m01 U27482 (.o(n23770),
	.a(proc_input_NIB_storage_data_f_1__31_),
	.b(FE_OFN373_n17762));
   oa12m01 U27483 (.o(n3573),
	.a(n23770),
	.b(FE_OFN373_n17762),
	.c(n23791));
   na02m01 U27484 (.o(n23771),
	.a(proc_input_NIB_storage_data_f_1__34_),
	.b(FE_OFN373_n17762));
   oa12m01 U27485 (.o(n3558),
	.a(n23771),
	.b(FE_OFN373_n17762),
	.c(n23816));
   oa12m01 U27486 (.o(n3543),
	.a(n23775),
	.b(FE_OFN373_n17762),
	.c(n23796));
   na02m01 U27487 (.o(n23776),
	.a(proc_input_NIB_storage_data_f_1__38_),
	.b(FE_OFN373_n17762));
   oa12m01 U27488 (.o(n3538),
	.a(n23776),
	.b(FE_OFN373_n17762),
	.c(n23812));
   na02m01 U27489 (.o(n23777),
	.a(proc_input_NIB_storage_data_f_1__40_),
	.b(FE_OFN373_n17762));
   oa12m01 U27490 (.o(n3528),
	.a(n23777),
	.b(FE_OFN373_n17762),
	.c(n23800));
   na02m01 U27491 (.o(n23784),
	.a(proc_input_NIB_storage_data_f_1__42_),
	.b(FE_OFN373_n17762));
   oa12m01 U27492 (.o(n3518),
	.a(n23784),
	.b(FE_OFN373_n17762),
	.c(n23808));
   na02m01 U27493 (.o(n23785),
	.a(proc_input_NIB_storage_data_f_1__43_),
	.b(FE_OFN373_n17762));
   oa12m01 U27494 (.o(n3513),
	.a(n23785),
	.b(FE_OFN373_n17762),
	.c(n23806));
   na02m01 U27495 (.o(n23809),
	.a(proc_input_NIB_storage_data_f_1__62_),
	.b(FE_OFN374_n17762));
   oa12m01 U27496 (.o(n3418),
	.a(n23809),
	.b(FE_OFN374_n17762),
	.c(n23810));
   na02m01 U27497 (.o(n23823),
	.a(proc_input_NIB_storage_data_f_1__63_),
	.b(FE_OFN374_n17762));
   oa12m01 U27498 (.o(n3413),
	.a(n23823),
	.b(FE_OFN374_n17762),
	.c(n23827));
   oa12m01 U27499 (.o(n3468),
	.a(n23831),
	.b(FE_OFN374_n17762),
	.c(n23890));
   na02m01 U27500 (.o(n23893),
	.a(proc_input_NIB_storage_data_f_1__30_),
	.b(FE_OFN373_n17762));
   oa12m01 U27501 (.o(n3578),
	.a(n23893),
	.b(FE_OFN373_n17762),
	.c(n23894));
   na02m01 U27502 (.o(n23900),
	.a(proc_input_NIB_storage_data_f_1__61_),
	.b(FE_OFN374_n17762));
   oa12m01 U27503 (.o(n3423),
	.a(n23900),
	.b(FE_OFN374_n17762),
	.c(n23918));
   na02m01 U27504 (.o(n23902),
	.a(proc_input_NIB_storage_data_f_1__50_),
	.b(FE_OFN374_n17762));
   oa12m01 U27505 (.o(n3478),
	.a(n23902),
	.b(FE_OFN374_n17762),
	.c(n23903));
   na02m01 U27506 (.o(n23904),
	.a(proc_input_NIB_storage_data_f_1__32_),
	.b(FE_OFN373_n17762));
   oa12m01 U27507 (.o(n3568),
	.a(n23904),
	.b(FE_OFN373_n17762),
	.c(n23905));
   na02m01 U27508 (.o(n23907),
	.a(proc_input_NIB_storage_data_f_1__49_),
	.b(FE_OFN373_n17762));
   oa12m01 U27509 (.o(n3483),
	.a(n23907),
	.b(FE_OFN373_n17762),
	.c(n23908));
   na02m01 U27510 (.o(n23909),
	.a(proc_input_NIB_storage_data_f_1__55_),
	.b(FE_OFN374_n17762));
   oa12m01 U27511 (.o(n3453),
	.a(n23909),
	.b(FE_OFN374_n17762),
	.c(n23910));
   na02m01 U27512 (.o(n23911),
	.a(proc_input_NIB_storage_data_f_1__48_),
	.b(FE_OFN373_n17762));
   oa12m01 U27513 (.o(n3488),
	.a(n23911),
	.b(FE_OFN373_n17762),
	.c(n23912));
   na02m01 U27514 (.o(n23913),
	.a(proc_input_NIB_storage_data_f_1__47_),
	.b(FE_OFN373_n17762));
   oa12m01 U27515 (.o(n3493),
	.a(n23913),
	.b(FE_OFN373_n17762),
	.c(n23914));
   na02m01 U27516 (.o(n23915),
	.a(proc_input_NIB_storage_data_f_1__46_),
	.b(FE_OFN373_n17762));
   oa12m01 U27517 (.o(n3498),
	.a(n23915),
	.b(FE_OFN373_n17762),
	.c(n23916));
   na02m01 U27518 (.o(n23919),
	.a(proc_input_NIB_storage_data_f_1__44_),
	.b(FE_OFN373_n17762));
   oa12m01 U27519 (.o(n3508),
	.a(n23919),
	.b(FE_OFN373_n17762),
	.c(n23920));
   na02m01 U27520 (.o(n23921),
	.a(proc_input_NIB_storage_data_f_1__53_),
	.b(FE_OFN373_n17762));
   oa12m01 U27521 (.o(n3463),
	.a(n23921),
	.b(FE_OFN373_n17762),
	.c(n23922));
   na02m01 U27522 (.o(n23923),
	.a(proc_input_NIB_storage_data_f_1__54_),
	.b(FE_OFN374_n17762));
   oa12m01 U27523 (.o(n3458),
	.a(n23923),
	.b(FE_OFN374_n17762),
	.c(n23924));
   na02m01 U27524 (.o(n23925),
	.a(proc_input_NIB_storage_data_f_1__60_),
	.b(FE_OFN374_n17762));
   oa12m01 U27525 (.o(n3428),
	.a(n23925),
	.b(FE_OFN374_n17762),
	.c(n23926));
   na02m01 U27526 (.o(n23927),
	.a(proc_input_NIB_storage_data_f_1__41_),
	.b(FE_OFN373_n17762));
   oa12m01 U27527 (.o(n3523),
	.a(n23927),
	.b(FE_OFN373_n17762),
	.c(n23928));
   na02m01 U27528 (.o(n23929),
	.a(proc_input_NIB_storage_data_f_1__56_),
	.b(FE_OFN374_n17762));
   oa12m01 U27529 (.o(n3448),
	.a(n23929),
	.b(FE_OFN374_n17762),
	.c(n23930));
   na02m01 U27530 (.o(n23931),
	.a(proc_input_NIB_storage_data_f_1__57_),
	.b(FE_OFN373_n17762));
   oa12m01 U27531 (.o(n3443),
	.a(n23931),
	.b(FE_OFN373_n17762),
	.c(n23932));
   na02m01 U27532 (.o(n23933),
	.a(proc_input_NIB_storage_data_f_1__39_),
	.b(FE_OFN373_n17762));
   oa12m01 U27533 (.o(n3533),
	.a(n23933),
	.b(FE_OFN373_n17762),
	.c(n23934));
   na02m01 U27534 (.o(n23935),
	.a(proc_input_NIB_storage_data_f_1__58_),
	.b(FE_OFN374_n17762));
   oa12m01 U27535 (.o(n3438),
	.a(n23935),
	.b(FE_OFN374_n17762),
	.c(n23936));
   na02m01 U27536 (.o(n23937),
	.a(proc_input_NIB_storage_data_f_1__59_),
	.b(FE_OFN374_n17762));
   oa12m01 U27537 (.o(n3433),
	.a(n23937),
	.b(FE_OFN374_n17762),
	.c(n23938));
   na02m01 U27538 (.o(n23939),
	.a(proc_input_NIB_storage_data_f_1__36_),
	.b(FE_OFN373_n17762));
   oa12m01 U27539 (.o(n3548),
	.a(n23939),
	.b(FE_OFN373_n17762),
	.c(n23940));
   na02m01 U27540 (.o(n23941),
	.a(proc_input_NIB_storage_data_f_1__45_),
	.b(FE_OFN373_n17762));
   oa12m01 U27541 (.o(n3503),
	.a(n23941),
	.b(FE_OFN373_n17762),
	.c(n23942));
   na02m01 U27542 (.o(n23943),
	.a(proc_input_NIB_storage_data_f_1__35_),
	.b(FE_OFN373_n17762));
   oa12m01 U27543 (.o(n3553),
	.a(n23943),
	.b(FE_OFN373_n17762),
	.c(n23944));
   na02m01 U27544 (.o(n23945),
	.a(proc_input_NIB_storage_data_f_1__51_),
	.b(FE_OFN374_n17762));
   oa12m01 U27545 (.o(n3473),
	.a(n23945),
	.b(FE_OFN374_n17762),
	.c(n23947));
   in01s01 U27546 (.o(n23955),
	.a(n23954));
   na02f02 U27547 (.o(n23962),
	.a(n23961),
	.b(n23960));
   in01s01 U27548 (.o(n23963),
	.a(n23962));
   na02f02 U27549 (.o(n23971),
	.a(n23970),
	.b(n23969));
   in01s01 U27551 (.o(n23981),
	.a(n23980));
   ao22m01 U27552 (.o(n23985),
	.a(FE_OFN259_n25295),
	.b(n23984),
	.c(n17787),
	.d(n23983));
   in01s01 U27553 (.o(n23989),
	.a(n23985));
   oa12f02 U27554 (.o(dataOut_P_22_),
	.a(n23990),
	.b(FE_OFN144_n23991),
	.c(n24728));
   in01s01 U27555 (.o(n23997),
	.a(n23996));
   no02f01 U27556 (.o(n23999),
	.a(n23998),
	.b(n23997));
   oa12f02 U27557 (.o(dataOut_P_54_),
	.a(n23999),
	.b(n24000),
	.c(FE_OFN524_n24728));
   in01s01 U27558 (.o(n24006),
	.a(n24005));
   ao22f01 U27559 (.o(n24014),
	.a(FE_OFN257_n25294),
	.b(FE_OFN487_n24013),
	.c(n17787),
	.d(n24012));
   na02f02 U27560 (.o(n24016),
	.a(n24015),
	.b(n24014));
   ao22f01 U27562 (.o(n24023),
	.a(n25294),
	.b(FE_OFN491_n24022),
	.c(n17787),
	.d(n24021));
   na02f02 U27563 (.o(n24025),
	.a(n24024),
	.b(n24023));
   na02f01 U27564 (.o(n24034),
	.a(n24033),
	.b(n24032));
   in01s01 U27565 (.o(n24035),
	.a(n24034));
   ao22f01 U27566 (.o(n24041),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__3_),
	.c(FE_OFN188_n24453),
	.d(proc_input_NIB_storage_data_f_2__3_));
   ao22f01 U27567 (.o(n24040),
	.a(n18077),
	.b(proc_input_NIB_storage_data_f_5__3_),
	.c(FE_OCPN25834_n),
	.d(proc_input_NIB_storage_data_f_0__3_));
   ao22f01 U27568 (.o(n24039),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__3_),
	.c(FE_OFN25645_n21748),
	.d(proc_input_NIB_storage_data_f_8__3_));
   ao22f01 U27569 (.o(n24038),
	.a(n20056),
	.b(proc_input_NIB_storage_data_f_9__3_),
	.c(n17742),
	.d(proc_input_NIB_storage_data_f_4__3_));
   ao22f01 U27570 (.o(n24045),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__3_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__3_));
   ao22f01 U27571 (.o(n24044),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__3_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__3_));
   ao22f01 U27572 (.o(n24043),
	.a(FE_OFN25635_n19595),
	.b(proc_input_NIB_storage_data_f_15__3_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__3_));
   ao22f01 U27573 (.o(n24049),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__3_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__3_));
   ao22f01 U27574 (.o(n24048),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__3_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__3_));
   na02f04 U27575 (.o(n24685),
	.a(n24049),
	.b(n24048));
   ao22f01 U27576 (.o(n24051),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__3_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__3_));
   ao22f01 U27577 (.o(n24050),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__3_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__3_));
   ao22f01 U27578 (.o(n24057),
	.a(n19019),
	.b(n24685),
	.c(n19017),
	.d(FE_OFN229_n24684));
   ao22f01 U27579 (.o(n24053),
	.a(FE_RN_13),
	.b(south_input_NIB_storage_data_f_3__3_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__3_));
   na02f02 U27580 (.o(n24687),
	.a(n24053),
	.b(n24052));
   ao22f01 U27581 (.o(n24055),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__3_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__3_));
   ao22f01 U27582 (.o(n24054),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__3_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__3_));
   na02f03 U27583 (.o(n24686),
	.a(n24055),
	.b(n24054));
   ao22f01 U27585 (.o(n24064),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__4_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__4_));
   ao22f01 U27586 (.o(n24063),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__4_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__4_));
   ao22f01 U27587 (.o(n24062),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__4_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__4_));
   ao22f01 U27588 (.o(n24061),
	.a(n24060),
	.b(proc_input_NIB_storage_data_f_9__4_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__4_));
   ao22f01 U27589 (.o(n24069),
	.a(FE_OCPN25814_FE_OFN186_n24453),
	.b(proc_input_NIB_storage_data_f_2__4_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__4_));
   ao22f01 U27590 (.o(n24068),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__4_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__4_));
   ao22f01 U27591 (.o(n24066),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__4_),
	.c(FE_OFN167_n24343),
	.d(proc_input_NIB_storage_data_f_8__4_));
   ao22f01 U27592 (.o(n24073),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__4_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__4_));
   ao22f01 U27593 (.o(n24072),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__4_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__4_));
   na02f02 U27594 (.o(n24702),
	.a(n24073),
	.b(n24072));
   ao22f01 U27595 (.o(n24075),
	.a(FE_RN_13),
	.b(south_input_NIB_storage_data_f_3__4_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__4_));
   ao22f01 U27596 (.o(n24074),
	.a(n21365),
	.b(south_input_NIB_storage_data_f_2__4_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__4_));
   ao22f01 U27597 (.o(n24077),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__4_),
	.c(FE_OFN24800_n20506),
	.d(east_input_NIB_storage_data_f_3__4_));
   ao22f01 U27598 (.o(n24076),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__4_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__4_));
   ao22f01 U27599 (.o(n24079),
	.a(FE_OFN28_n18974),
	.b(west_input_NIB_storage_data_f_0__4_),
	.c(n24466),
	.d(west_input_NIB_storage_data_f_2__4_));
   ao22f01 U27600 (.o(n24078),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__4_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__4_));
   na02f02 U27601 (.o(n24705),
	.a(n24079),
	.b(n24078));
   na02f02 U27602 (.o(n24082),
	.a(n24081),
	.b(n24080));
   in01s01 U27603 (.o(n24083),
	.a(n24082));
   ao22f01 U27604 (.o(n24087),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__1_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__1_));
   ao22f01 U27605 (.o(n24086),
	.a(FE_OCPN25814_FE_OFN186_n24453),
	.b(proc_input_NIB_storage_data_f_2__1_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__1_));
   ao22f01 U27606 (.o(n24085),
	.a(FE_OFN24731_n18131),
	.b(proc_input_NIB_storage_data_f_0__1_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__1_));
   ao22f01 U27607 (.o(n24084),
	.a(FE_OFN25680_n17814),
	.b(proc_input_NIB_storage_data_f_9__1_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__1_));
   ao22f01 U27608 (.o(n24092),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__1_),
	.c(FE_OFN168_n24343),
	.d(proc_input_NIB_storage_data_f_8__1_));
   ao22f01 U27609 (.o(n24091),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__1_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__1_));
   ao22f01 U27610 (.o(n24090),
	.a(n24454),
	.b(proc_input_NIB_storage_data_f_13__1_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__1_));
   ao22f01 U27611 (.o(n24089),
	.a(n19707),
	.b(proc_input_NIB_storage_data_f_3__1_),
	.c(FE_OCPN25954_n18039),
	.d(proc_input_NIB_storage_data_f_10__1_));
   ao22f01 U27612 (.o(n24096),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__1_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__1_));
   ao22f01 U27613 (.o(n24095),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__1_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__1_));
   na02f04 U27614 (.o(n24663),
	.a(n24096),
	.b(n24095));
   ao22f01 U27615 (.o(n24098),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__1_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__1_));
   ao22f01 U27616 (.o(n24097),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__1_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__1_));
   ao22f01 U27617 (.o(n24100),
	.a(FE_OFN24788_n24965),
	.b(south_input_NIB_storage_data_f_3__1_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__1_));
   ao22f01 U27618 (.o(n24099),
	.a(n17782),
	.b(south_input_NIB_storage_data_f_2__1_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__1_));
   ao22f01 U27619 (.o(n24102),
	.a(FE_OFN28_n18974),
	.b(west_input_NIB_storage_data_f_0__1_),
	.c(n24466),
	.d(west_input_NIB_storage_data_f_2__1_));
   ao22f01 U27620 (.o(n24101),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__1_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__1_));
   na02f04 U27621 (.o(n24665),
	.a(n24102),
	.b(n24101));
   na02f02 U27622 (.o(n24105),
	.a(n24104),
	.b(n24103));
   ao22f01 U27624 (.o(n24110),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__11_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__11_));
   ao22f01 U27625 (.o(n24107),
	.a(FE_OCPN25909_n19547),
	.b(proc_input_NIB_storage_data_f_11__11_),
	.c(FE_OFN168_n24343),
	.d(proc_input_NIB_storage_data_f_8__11_));
   ao22f01 U27626 (.o(n24113),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__11_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__11_));
   ao22f01 U27627 (.o(n24112),
	.a(n19707),
	.b(proc_input_NIB_storage_data_f_3__11_),
	.c(FE_OCPN25837_n24342),
	.d(proc_input_NIB_storage_data_f_0__11_));
   ao22f01 U27628 (.o(n24111),
	.a(FE_OFN25680_n17814),
	.b(proc_input_NIB_storage_data_f_9__11_),
	.c(FE_OCPN25954_n18039),
	.d(proc_input_NIB_storage_data_f_10__11_));
   ao22f01 U27629 (.o(n24118),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__11_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__11_));
   na02f02 U27631 (.o(n24577),
	.a(n24118),
	.b(n24117));
   ao22f01 U27632 (.o(n24120),
	.a(FE_OCPN25935_n24965),
	.b(south_input_NIB_storage_data_f_3__11_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__11_));
   ao22f01 U27633 (.o(n24119),
	.a(n17782),
	.b(south_input_NIB_storage_data_f_2__11_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__11_));
   na02f02 U27634 (.o(n24576),
	.a(n24120),
	.b(n24119));
   ao22f01 U27635 (.o(n24122),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__11_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__11_));
   ao22f01 U27636 (.o(n24121),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__11_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__11_));
   ao22f01 U27637 (.o(n24124),
	.a(FE_OFN28_n18974),
	.b(west_input_NIB_storage_data_f_0__11_),
	.c(FE_RN_27),
	.d(west_input_NIB_storage_data_f_1__11_));
   ao22f01 U27638 (.o(n24123),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__11_),
	.c(n24466),
	.d(west_input_NIB_storage_data_f_2__11_));
   na02f02 U27639 (.o(n24579),
	.a(n24124),
	.b(n24123));
   na02f02 U27640 (.o(n24127),
	.a(n24126),
	.b(n24125));
   in01s01 U27641 (.o(n24128),
	.a(n24127));
   ao22f01 U27642 (.o(n24133),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__2_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__2_));
   ao22f01 U27643 (.o(n24131),
	.a(FE_OCPN25834_n),
	.b(proc_input_NIB_storage_data_f_0__2_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__2_));
   ao22f01 U27644 (.o(n24130),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__2_),
	.c(FE_RN_51),
	.d(proc_input_NIB_storage_data_f_1__2_));
   ao22f01 U27645 (.o(n24137),
	.a(n18077),
	.b(proc_input_NIB_storage_data_f_5__2_),
	.c(FE_OFN25645_n21748),
	.d(proc_input_NIB_storage_data_f_8__2_));
   ao22f01 U27646 (.o(n24136),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__2_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__2_));
   ao22f01 U27647 (.o(n24135),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__2_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__2_));
   ao22f01 U27648 (.o(n24134),
	.a(n24060),
	.b(proc_input_NIB_storage_data_f_9__2_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__2_));
   no02f04 U27649 (.o(n24701),
	.a(n24139),
	.b(n24138));
   ao22f01 U27650 (.o(n24141),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__2_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__2_));
   ao22f01 U27651 (.o(n24140),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__2_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__2_));
   ao22f01 U27652 (.o(n24143),
	.a(n21365),
	.b(south_input_NIB_storage_data_f_2__2_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__2_));
   na02f02 U27653 (.o(n24694),
	.a(n24144),
	.b(n24143));
   ao22f01 U27654 (.o(n24146),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__2_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__2_));
   ao22f01 U27655 (.o(n24145),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__2_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__2_));
   na02f02 U27656 (.o(n24695),
	.a(n24146),
	.b(n24145));
   ao22f01 U27657 (.o(n24148),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__2_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__2_));
   ao22f01 U27658 (.o(n24147),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__2_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__2_));
   na02f02 U27659 (.o(n24696),
	.a(n24148),
	.b(n24147));
   na02f02 U27660 (.o(n24151),
	.a(n24150),
	.b(n24149));
   in01s01 U27661 (.o(n24152),
	.a(n24151));
   ao22f01 U27662 (.o(n24156),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__17_),
	.c(FE_OFN188_n24453),
	.d(proc_input_NIB_storage_data_f_2__17_));
   ao22f01 U27663 (.o(n24155),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__17_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__17_));
   ao22f01 U27664 (.o(n24153),
	.a(n20056),
	.b(proc_input_NIB_storage_data_f_9__17_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__17_));
   ao22f01 U27665 (.o(n24160),
	.a(n24454),
	.b(proc_input_NIB_storage_data_f_13__17_),
	.c(FE_OFN25645_n21748),
	.d(proc_input_NIB_storage_data_f_8__17_));
   ao22f01 U27666 (.o(n24159),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__17_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__17_));
   ao22f01 U27667 (.o(n24157),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__17_),
	.c(FE_OFN165_n24129),
	.d(proc_input_NIB_storage_data_f_1__17_));
   ao22f01 U27668 (.o(n24164),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__17_),
	.c(FE_OFN24800_n20506),
	.d(east_input_NIB_storage_data_f_3__17_));
   ao22f01 U27669 (.o(n24163),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__17_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__17_));
   ao22f01 U27670 (.o(n24167),
	.a(FE_OCPN25938_n24965),
	.b(south_input_NIB_storage_data_f_3__17_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__17_));
   ao22f01 U27671 (.o(n24166),
	.a(n24165),
	.b(south_input_NIB_storage_data_f_2__17_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__17_));
   na02f02 U27672 (.o(n24638),
	.a(n24167),
	.b(n24166));
   ao22f01 U27673 (.o(n24173),
	.a(FE_OFN44_n19054),
	.b(FE_OFN217_n24637),
	.c(FE_OFN366_n17753),
	.d(n24638));
   ao22f01 U27674 (.o(n24169),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__17_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__17_));
   ao22f01 U27675 (.o(n24168),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__17_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__17_));
   na02f04 U27676 (.o(n24639),
	.a(n24169),
	.b(n24168));
   ao22f01 U27677 (.o(n24171),
	.a(FE_OFN28_n18974),
	.b(west_input_NIB_storage_data_f_0__17_),
	.c(n24466),
	.d(west_input_NIB_storage_data_f_2__17_));
   ao22f01 U27678 (.o(n24170),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__17_),
	.c(FE_RN_27),
	.d(west_input_NIB_storage_data_f_1__17_));
   na02f02 U27679 (.o(n24640),
	.a(n24171),
	.b(n24170));
   na02f02 U27680 (.o(n24174),
	.a(n24173),
	.b(n24172));
   ao22f01 U27682 (.o(n24179),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__20_),
	.c(FE_OCPN25828_n21745),
	.d(proc_input_NIB_storage_data_f_2__20_));
   ao22f01 U27683 (.o(n24178),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__20_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__20_));
   ao22f02 U27684 (.o(n24176),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__20_),
	.c(FE_OCPN25819_n24342),
	.d(proc_input_NIB_storage_data_f_0__20_));
   ao22f01 U27685 (.o(n24182),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__20_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__20_));
   ao22f01 U27686 (.o(n24181),
	.a(FE_OCPN25909_n19547),
	.b(proc_input_NIB_storage_data_f_11__20_),
	.c(n17743),
	.d(proc_input_NIB_storage_data_f_4__20_));
   ao22f01 U27687 (.o(n24180),
	.a(n24060),
	.b(proc_input_NIB_storage_data_f_9__20_),
	.c(FE_OFN167_n24343),
	.d(proc_input_NIB_storage_data_f_8__20_));
   ao22f01 U27688 (.o(n24187),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__20_),
	.c(FE_OFN24800_n20506),
	.d(east_input_NIB_storage_data_f_3__20_));
   ao22f01 U27689 (.o(n24186),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__20_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__20_));
   ao22f01 U27690 (.o(n24189),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__20_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__20_));
   ao22f01 U27691 (.o(n24188),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__20_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__20_));
   na02f04 U27692 (.o(n24721),
	.a(n24189),
	.b(n24188));
   ao22f01 U27693 (.o(n24191),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__20_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__20_));
   ao22f01 U27694 (.o(n24190),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__20_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__20_));
   na02f02 U27695 (.o(n24723),
	.a(n24191),
	.b(n24190));
   ao22f01 U27696 (.o(n24193),
	.a(FE_OCPN25938_n24965),
	.b(south_input_NIB_storage_data_f_3__20_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__20_));
   ao22f01 U27697 (.o(n24192),
	.a(n21365),
	.b(south_input_NIB_storage_data_f_2__20_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__20_));
   na02f02 U27698 (.o(n24722),
	.a(n24193),
	.b(n24192));
   na02f02 U27699 (.o(n24196),
	.a(n24195),
	.b(n24194));
   ao22f01 U27701 (.o(n24201),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__19_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__19_));
   ao22f01 U27702 (.o(n24200),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__19_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__19_));
   ao22f01 U27703 (.o(n24199),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__19_),
	.c(FE_OFN25645_n21748),
	.d(proc_input_NIB_storage_data_f_8__19_));
   ao22f01 U27704 (.o(n24198),
	.a(n17754),
	.b(proc_input_NIB_storage_data_f_3__19_),
	.c(n24060),
	.d(proc_input_NIB_storage_data_f_9__19_));
   ao22f01 U27705 (.o(n24203),
	.a(FE_OCPN25834_n),
	.b(proc_input_NIB_storage_data_f_0__19_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__19_));
   ao22f01 U27706 (.o(n24210),
	.a(FE_OCPN25937_n24965),
	.b(south_input_NIB_storage_data_f_3__19_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__19_));
   ao22f01 U27707 (.o(n24209),
	.a(n24142),
	.b(south_input_NIB_storage_data_f_2__19_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__19_));
   na02f02 U27708 (.o(n24740),
	.a(n24210),
	.b(n24209));
   ao22f01 U27709 (.o(n24212),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__19_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__19_));
   ao22f01 U27710 (.o(n24211),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__19_),
	.c(FE_RN_27),
	.d(west_input_NIB_storage_data_f_1__19_));
   ao22f01 U27711 (.o(n24214),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__19_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__19_));
   ao22f01 U27712 (.o(n24213),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__19_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__19_));
   na02f03 U27713 (.o(n24742),
	.a(n24214),
	.b(n24213));
   ao22f01 U27714 (.o(n24216),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__19_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__19_));
   ao22f01 U27715 (.o(n24215),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__19_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__19_));
   na02f02 U27716 (.o(n24219),
	.a(n24218),
	.b(n24217));
   in01s01 U27717 (.o(n24220),
	.a(n24219));
   ao22f01 U27718 (.o(n24225),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__15_),
	.c(FE_OFN25689_n19503),
	.d(proc_input_NIB_storage_data_f_6__15_));
   ao22m02 U27719 (.o(n24224),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__15_),
	.c(FE_OCPN25834_n),
	.d(proc_input_NIB_storage_data_f_0__15_));
   ao22f01 U27720 (.o(n24223),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__15_),
	.c(n17743),
	.d(proc_input_NIB_storage_data_f_4__15_));
   ao22f01 U27721 (.o(n24222),
	.a(n21768),
	.b(proc_input_NIB_storage_data_f_3__15_),
	.c(n24060),
	.d(proc_input_NIB_storage_data_f_9__15_));
   ao22f01 U27722 (.o(n24229),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__15_),
	.c(FE_OCPN25954_n18039),
	.d(proc_input_NIB_storage_data_f_10__15_));
   ao22f01 U27723 (.o(n24226),
	.a(FE_RN_51),
	.b(proc_input_NIB_storage_data_f_1__15_),
	.c(n24343),
	.d(proc_input_NIB_storage_data_f_8__15_));
   ao22f01 U27724 (.o(n24233),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__15_),
	.c(FE_OFN24800_n20506),
	.d(east_input_NIB_storage_data_f_3__15_));
   ao22f01 U27725 (.o(n24232),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__15_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__15_));
   ao22f01 U27726 (.o(n24235),
	.a(n24472),
	.b(south_input_NIB_storage_data_f_0__15_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__15_));
   ao22f01 U27727 (.o(n24234),
	.a(FE_OCPN25940_n24965),
	.b(south_input_NIB_storage_data_f_3__15_),
	.c(FE_OFN25648_n18762),
	.d(south_input_NIB_storage_data_f_2__15_));
   na02f02 U27728 (.o(n24620),
	.a(n24235),
	.b(n24234));
   ao22f01 U27729 (.o(n24241),
	.a(n19054),
	.b(FE_OFN207_n24619),
	.c(FE_OFN366_n17753),
	.d(n24620));
   ao22f01 U27730 (.o(n24237),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__15_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__15_));
   ao22f01 U27731 (.o(n24236),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__15_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__15_));
   na02f03 U27732 (.o(n24621),
	.a(n24237),
	.b(n24236));
   ao22f01 U27733 (.o(n24239),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__15_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__15_));
   ao22f01 U27734 (.o(n24238),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__15_),
	.c(FE_RN_27),
	.d(west_input_NIB_storage_data_f_1__15_));
   na02f04 U27735 (.o(n24622),
	.a(n24239),
	.b(n24238));
   na02f02 U27736 (.o(n24242),
	.a(n24241),
	.b(n24240));
   in01s01 U27737 (.o(n24243),
	.a(n24242));
   ao22f01 U27738 (.o(n24248),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__14_),
	.c(FE_OFN20_n17779),
	.d(proc_input_NIB_storage_data_f_7__14_));
   ao22f01 U27739 (.o(n24246),
	.a(n24454),
	.b(proc_input_NIB_storage_data_f_13__14_),
	.c(n17743),
	.d(proc_input_NIB_storage_data_f_4__14_));
   ao22f01 U27740 (.o(n24245),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__14_),
	.c(n19705),
	.d(proc_input_NIB_storage_data_f_9__14_));
   ao22f01 U27741 (.o(n24252),
	.a(FE_OCPN25827_n21745),
	.b(proc_input_NIB_storage_data_f_2__14_),
	.c(FE_OCPN25954_n18039),
	.d(proc_input_NIB_storage_data_f_10__14_));
   ao22f01 U27743 (.o(n24250),
	.a(n21768),
	.b(proc_input_NIB_storage_data_f_3__14_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__14_));
   ao22f01 U27744 (.o(n24249),
	.a(FE_OFN161_n24129),
	.b(proc_input_NIB_storage_data_f_1__14_),
	.c(FE_OFN167_n24343),
	.d(proc_input_NIB_storage_data_f_8__14_));
   ao22f01 U27745 (.o(n24256),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__14_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__14_));
   ao22f01 U27746 (.o(n24255),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__14_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__14_));
   na02f02 U27747 (.o(n24676),
	.a(n24256),
	.b(n24255));
   ao22f01 U27748 (.o(n24258),
	.a(FE_OCPN25937_n24965),
	.b(south_input_NIB_storage_data_f_3__14_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__14_));
   ao22f01 U27749 (.o(n24257),
	.a(n17782),
	.b(south_input_NIB_storage_data_f_2__14_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__14_));
   na02f02 U27750 (.o(n24675),
	.a(n24258),
	.b(n24257));
   ao22f01 U27751 (.o(n24259),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__14_),
	.c(FE_OFN24800_n20506),
	.d(east_input_NIB_storage_data_f_3__14_));
   ao22f01 U27752 (.o(n24262),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__14_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__14_));
   ao22f01 U27753 (.o(n24261),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__14_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__14_));
   na02f04 U27754 (.o(n24678),
	.a(n24262),
	.b(n24261));
   na02f02 U27755 (.o(n24265),
	.a(n24264),
	.b(n24263));
   ao22f01 U27757 (.o(n24270),
	.a(n18077),
	.b(proc_input_NIB_storage_data_f_5__13_),
	.c(FE_OFN20_n17779),
	.d(proc_input_NIB_storage_data_f_7__13_));
   ao22f01 U27758 (.o(n24267),
	.a(n19709),
	.b(proc_input_NIB_storage_data_f_3__13_),
	.c(n24060),
	.d(proc_input_NIB_storage_data_f_9__13_));
   ao22f01 U27759 (.o(n24274),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__13_),
	.c(FE_OFN25604_n19530),
	.d(proc_input_NIB_storage_data_f_13__13_));
   ao22f01 U27760 (.o(n24273),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__13_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__13_));
   ao22f01 U27761 (.o(n24272),
	.a(FE_OFN25635_n19595),
	.b(proc_input_NIB_storage_data_f_15__13_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__13_));
   ao22f01 U27762 (.o(n24271),
	.a(FE_OFN25645_n21748),
	.b(proc_input_NIB_storage_data_f_8__13_),
	.c(n17743),
	.d(proc_input_NIB_storage_data_f_4__13_));
   ao22f01 U27763 (.o(n24278),
	.a(FE_RN_13),
	.b(south_input_NIB_storage_data_f_3__13_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__13_));
   ao22f01 U27764 (.o(n24277),
	.a(n17782),
	.b(south_input_NIB_storage_data_f_2__13_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__13_));
   na02f02 U27765 (.o(n24598),
	.a(n24278),
	.b(n24277));
   ao22f01 U27766 (.o(n24280),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__13_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__13_));
   ao22f01 U27767 (.o(n24279),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__13_),
	.c(FE_RN_27),
	.d(west_input_NIB_storage_data_f_1__13_));
   na02f02 U27768 (.o(n24599),
	.a(n24280),
	.b(n24279));
   ao22f01 U27769 (.o(n24282),
	.a(FE_OFN24771_n19075),
	.b(north_input_NIB_storage_data_f_0__13_),
	.c(n19220),
	.d(north_input_NIB_storage_data_f_2__13_));
   ao22f01 U27770 (.o(n24281),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__13_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__13_));
   ao22f01 U27771 (.o(n24284),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__13_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__13_));
   ao22f01 U27772 (.o(n24283),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__13_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__13_));
   na02f02 U27773 (.o(n24287),
	.a(n24286),
	.b(n24285));
   in01s01 U27774 (.o(n24288),
	.a(n24287));
   ao22f01 U27775 (.o(n24292),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__12_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__12_));
   ao22f01 U27776 (.o(n24291),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__12_),
	.c(n21768),
	.d(proc_input_NIB_storage_data_f_3__12_));
   ao22f01 U27777 (.o(n24290),
	.a(FE_OCPN25837_n24342),
	.b(proc_input_NIB_storage_data_f_0__12_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__12_));
   ao22f01 U27778 (.o(n24289),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__12_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__12_));
   ao22f01 U27779 (.o(n24296),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__12_),
	.c(FE_OFN168_n24343),
	.d(proc_input_NIB_storage_data_f_8__12_));
   ao22f01 U27780 (.o(n24295),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__12_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__12_));
   ao22f01 U27781 (.o(n24294),
	.a(FE_OCPN25814_FE_OFN186_n24453),
	.b(proc_input_NIB_storage_data_f_2__12_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__12_));
   ao22f01 U27782 (.o(n24293),
	.a(FE_OFN25680_n17814),
	.b(proc_input_NIB_storage_data_f_9__12_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__12_));
   ao22f01 U27783 (.o(n24300),
	.a(n19193),
	.b(north_input_NIB_storage_data_f_3__12_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__12_));
   ao22f01 U27784 (.o(n24299),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__12_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__12_));
   na02f02 U27785 (.o(n24586),
	.a(n24300),
	.b(n24299));
   ao22f01 U27786 (.o(n24302),
	.a(FE_OCPN25939_n24965),
	.b(south_input_NIB_storage_data_f_3__12_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__12_));
   ao22f01 U27787 (.o(n24301),
	.a(n24142),
	.b(south_input_NIB_storage_data_f_2__12_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__12_));
   na02m02 U27788 (.o(n24585),
	.a(n24302),
	.b(n24301));
   ao22f01 U27789 (.o(n24304),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__12_),
	.c(FE_OFN24800_n20506),
	.d(east_input_NIB_storage_data_f_3__12_));
   ao22f01 U27790 (.o(n24303),
	.a(FE_OFN24778_n19932),
	.b(east_input_NIB_storage_data_f_0__12_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__12_));
   ao22f01 U27791 (.o(n24306),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__12_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__12_));
   ao22f01 U27792 (.o(n24305),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__12_),
	.c(FE_RN_27),
	.d(west_input_NIB_storage_data_f_1__12_));
   na02f02 U27793 (.o(n24588),
	.a(n24306),
	.b(n24305));
   na02f02 U27794 (.o(n24309),
	.a(n24308),
	.b(n24307));
   ao22f01 U27796 (.o(n24314),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__21_),
	.c(FE_OCPN25814_FE_OFN186_n24453),
	.d(proc_input_NIB_storage_data_f_2__21_));
   ao22f01 U27797 (.o(n24313),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__21_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__21_));
   ao22f01 U27798 (.o(n24311),
	.a(n20056),
	.b(proc_input_NIB_storage_data_f_9__21_),
	.c(FE_OCPN25834_n),
	.d(proc_input_NIB_storage_data_f_0__21_));
   ao22f01 U27799 (.o(n24318),
	.a(n24454),
	.b(proc_input_NIB_storage_data_f_13__21_),
	.c(FE_OFN168_n24343),
	.d(proc_input_NIB_storage_data_f_8__21_));
   ao22f01 U27800 (.o(n24316),
	.a(n17754),
	.b(proc_input_NIB_storage_data_f_3__21_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__21_));
   ao22f01 U27801 (.o(n24315),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__21_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__21_));
   ao22f01 U27802 (.o(n24323),
	.a(FE_OFN24788_n24965),
	.b(south_input_NIB_storage_data_f_3__21_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__21_));
   ao22f01 U27803 (.o(n24322),
	.a(n24321),
	.b(south_input_NIB_storage_data_f_2__21_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__21_));
   na02m02 U27804 (.o(n24711),
	.a(n24323),
	.b(n24322));
   ao22f01 U27805 (.o(n24325),
	.a(FE_OFN24771_n19075),
	.b(north_input_NIB_storage_data_f_0__21_),
	.c(n19220),
	.d(north_input_NIB_storage_data_f_2__21_));
   ao22f01 U27806 (.o(n24324),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__21_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__21_));
   na02f02 U27807 (.o(n24712),
	.a(n24325),
	.b(n24324));
   ao22m02 U27808 (.o(n24327),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__21_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__21_));
   ao22m02 U27809 (.o(n24326),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__21_),
	.c(FE_RN_31),
	.d(west_input_NIB_storage_data_f_1__21_));
   na02f03 U27810 (.o(n24714),
	.a(n24327),
	.b(n24326));
   ao22f01 U27811 (.o(n24329),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__21_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__21_));
   ao22f01 U27812 (.o(n24328),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__21_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__21_));
   ao22f01 U27813 (.o(n24330),
	.a(n19019),
	.b(n24714),
	.c(n19017),
	.d(n24713));
   in01s01 U27814 (.o(n24333),
	.a(n24332));
   in01s01 U27816 (.o(n24341),
	.a(n24340));
   ao22f01 U27817 (.o(n24348),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__0_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__0_));
   ao22f02 U27818 (.o(n24347),
	.a(FE_OCPN25834_n),
	.b(proc_input_NIB_storage_data_f_0__0_),
	.c(FE_RN_51),
	.d(proc_input_NIB_storage_data_f_1__0_));
   ao22f01 U27819 (.o(n24346),
	.a(n17754),
	.b(proc_input_NIB_storage_data_f_3__0_),
	.c(FE_OFN25645_n21748),
	.d(proc_input_NIB_storage_data_f_8__0_));
   ao22m02 U27820 (.o(n24345),
	.a(n24060),
	.b(proc_input_NIB_storage_data_f_9__0_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__0_));
   ao22f01 U27821 (.o(n24354),
	.a(FE_RN_49),
	.b(proc_input_NIB_storage_data_f_5__0_),
	.c(FE_OCPN25954_n18039),
	.d(proc_input_NIB_storage_data_f_10__0_));
   ao22f01 U27822 (.o(n24353),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__0_),
	.c(n24454),
	.d(proc_input_NIB_storage_data_f_13__0_));
   ao22f01 U27823 (.o(n24352),
	.a(FE_OFN188_n24453),
	.b(proc_input_NIB_storage_data_f_2__0_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__0_));
   ao22f01 U27824 (.o(n24351),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__0_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__0_));
   ao22m02 U27825 (.o(n24358),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__0_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__0_));
   ao22f01 U27826 (.o(n24357),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__0_),
	.c(FE_RN_27),
	.d(west_input_NIB_storage_data_f_1__0_));
   na02f02 U27827 (.o(n24732),
	.a(n24358),
	.b(n24357));
   ao22f01 U27828 (.o(n24361),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__0_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__0_));
   ao22f01 U27829 (.o(n24360),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__0_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__0_));
   ao22f01 U27830 (.o(n24363),
	.a(FE_RN_13),
	.b(south_input_NIB_storage_data_f_3__0_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__0_));
   ao22f01 U27831 (.o(n24362),
	.a(n17782),
	.b(south_input_NIB_storage_data_f_2__0_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__0_));
   na02f02 U27832 (.o(n24734),
	.a(n24363),
	.b(n24362));
   ao22f01 U27833 (.o(n24367),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__0_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__0_));
   ao22f01 U27834 (.o(n24366),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__0_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__0_));
   na02f02 U27835 (.o(n24733),
	.a(n24367),
	.b(n24366));
   ao22f01 U27836 (.o(n24373),
	.a(n19019),
	.b(n24721),
	.c(n19017),
	.d(n24720));
   na02f02 U27837 (.o(n24374),
	.a(n24373),
	.b(n24372));
   ao22f01 U27839 (.o(n24376),
	.a(n19017),
	.b(FE_OFN242_n24744),
	.c(n19020),
	.d(n24742));
   na02f02 U27840 (.o(n24378),
	.a(n24377),
	.b(n24376));
   ao22f01 U27842 (.o(n24382),
	.a(FE_OFN25688_n19500),
	.b(proc_input_NIB_storage_data_f_12__18_),
	.c(FE_OFN25644_n19504),
	.d(proc_input_NIB_storage_data_f_14__18_));
   ao22f02 U27843 (.o(n24380),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__18_),
	.c(n21740),
	.d(proc_input_NIB_storage_data_f_0__18_));
   ao22f01 U27844 (.o(n24387),
	.a(n19503),
	.b(proc_input_NIB_storage_data_f_6__18_),
	.c(FE_OFN168_n24343),
	.d(proc_input_NIB_storage_data_f_8__18_));
   ao22f01 U27845 (.o(n24386),
	.a(n24454),
	.b(proc_input_NIB_storage_data_f_13__18_),
	.c(FE_OFN25635_n19595),
	.d(proc_input_NIB_storage_data_f_15__18_));
   ao22f01 U27846 (.o(n24384),
	.a(FE_OFN25680_n17814),
	.b(proc_input_NIB_storage_data_f_9__18_),
	.c(n21749),
	.d(proc_input_NIB_storage_data_f_4__18_));
   ao22m02 U27847 (.o(n24392),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__18_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__18_));
   ao22f01 U27848 (.o(n24391),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__18_),
	.c(FE_RN_27),
	.d(west_input_NIB_storage_data_f_1__18_));
   na02f02 U27849 (.o(n24751),
	.a(n24392),
	.b(n24391));
   ao22f01 U27850 (.o(n24394),
	.a(FE_OCPN25935_n24965),
	.b(south_input_NIB_storage_data_f_3__18_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__18_));
   ao22f01 U27851 (.o(n24393),
	.a(n17782),
	.b(south_input_NIB_storage_data_f_2__18_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__18_));
   na02f02 U27852 (.o(n24750),
	.a(n24394),
	.b(n24393));
   ao22f01 U27853 (.o(n24401),
	.a(n19019),
	.b(FE_OFN546_n24751),
	.c(FE_OFN42_n19022),
	.d(n24750));
   ao22f01 U27854 (.o(n24396),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__18_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__18_));
   ao22f01 U27855 (.o(n24395),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__18_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__18_));
   ao22f01 U27856 (.o(n24399),
	.a(FE_OFN24771_n19075),
	.b(north_input_NIB_storage_data_f_0__18_),
	.c(n19220),
	.d(north_input_NIB_storage_data_f_2__18_));
   ao22f01 U27857 (.o(n24398),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__18_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__18_));
   na02f03 U27858 (.o(n24754),
	.a(n24399),
	.b(n24398));
   ao22f01 U27859 (.o(n24400),
	.a(n19017),
	.b(n24752),
	.c(n19020),
	.d(n24754));
   na02f02 U27860 (.o(n24402),
	.a(n24401),
	.b(n24400));
   na02f02 U27862 (.o(n24406),
	.a(n24405),
	.b(n24404));
   ao22f01 U27863 (.o(n24409),
	.a(n19017),
	.b(FE_OFN217_n24637),
	.c(n19022),
	.d(n24638));
   ao22f01 U27864 (.o(n24408),
	.a(n19019),
	.b(n24640),
	.c(n19020),
	.d(n24639));
   na02f02 U27865 (.o(n24410),
	.a(n24409),
	.b(n24408));
   ao22f01 U27867 (.o(n24413),
	.a(n19017),
	.b(FE_OFN207_n24619),
	.c(n19022),
	.d(n24620));
   na02f02 U27868 (.o(n24418),
	.a(n24417),
	.b(n24416));
   ao22f01 U27870 (.o(n24420),
	.a(n19019),
	.b(n24678),
	.c(n19017),
	.d(FE_OFN227_n24677));
   in01s01 U27871 (.o(n24423),
	.a(n24422));
   ao22f01 U27872 (.o(n24425),
	.a(n19019),
	.b(n24599),
	.c(n19022),
	.d(n24598));
   in01s01 U27873 (.o(n24427),
	.a(n24426));
   na02f02 U27876 (.o(n24438),
	.a(n24437),
	.b(n24436));
   in01s01 U27877 (.o(n24443),
	.a(n24442));
   na02f02 U27878 (.o(n24446),
	.a(n24445),
	.b(n24444));
   in01s01 U27879 (.o(n24447),
	.a(n24446));
   ao22f01 U27880 (.o(n24452),
	.a(FE_OFN20_n17779),
	.b(proc_input_NIB_storage_data_f_7__16_),
	.c(n19503),
	.d(proc_input_NIB_storage_data_f_6__16_));
   ao22f01 U27881 (.o(n24450),
	.a(FE_OFN25644_n19504),
	.b(proc_input_NIB_storage_data_f_14__16_),
	.c(n17742),
	.d(proc_input_NIB_storage_data_f_4__16_));
   ao22f01 U27882 (.o(n24449),
	.a(FE_OCPN25954_n18039),
	.b(proc_input_NIB_storage_data_f_10__16_),
	.c(FE_OFN161_n24129),
	.d(proc_input_NIB_storage_data_f_1__16_));
   ao22f01 U27883 (.o(n24459),
	.a(FE_OCPN25814_FE_OFN186_n24453),
	.b(proc_input_NIB_storage_data_f_2__16_),
	.c(FE_OFN168_n24343),
	.d(proc_input_NIB_storage_data_f_8__16_));
   ao22f01 U27884 (.o(n24457),
	.a(FE_OFN25635_n19595),
	.b(proc_input_NIB_storage_data_f_15__16_),
	.c(FE_OCPN25909_n19547),
	.d(proc_input_NIB_storage_data_f_11__16_));
   no02f02 U27885 (.o(n24636),
	.a(n24461),
	.b(n24460));
   ao22f01 U27886 (.o(n24464),
	.a(n25428),
	.b(north_input_NIB_storage_data_f_3__16_),
	.c(FE_OFN24771_n19075),
	.d(north_input_NIB_storage_data_f_0__16_));
   ao22f01 U27887 (.o(n24463),
	.a(n19220),
	.b(north_input_NIB_storage_data_f_2__16_),
	.c(FE_OFN178_n24364),
	.d(north_input_NIB_storage_data_f_1__16_));
   na02f04 U27888 (.o(n24628),
	.a(n24464),
	.b(n24463));
   ao22f01 U27889 (.o(n24468),
	.a(FE_OCPN25811_n18959),
	.b(west_input_NIB_storage_data_f_3__16_),
	.c(FE_OFN28_n18974),
	.d(west_input_NIB_storage_data_f_0__16_));
   ao22f01 U27890 (.o(n24467),
	.a(n24466),
	.b(west_input_NIB_storage_data_f_2__16_),
	.c(FE_RN_27),
	.d(west_input_NIB_storage_data_f_1__16_));
   na02f04 U27891 (.o(n24629),
	.a(n24468),
	.b(n24467));
   ao22f01 U27892 (.o(n24471),
	.a(FE_OFN25659_n19914),
	.b(east_input_NIB_storage_data_f_2__16_),
	.c(FE_OFN24799_n20506),
	.d(east_input_NIB_storage_data_f_3__16_));
   ao22f01 U27893 (.o(n24470),
	.a(FE_OFN24779_n19932),
	.b(east_input_NIB_storage_data_f_0__16_),
	.c(FE_OCPN25905_n19306),
	.d(east_input_NIB_storage_data_f_1__16_));
   ao22f01 U27894 (.o(n24475),
	.a(FE_OCPN25936_n24965),
	.b(south_input_NIB_storage_data_f_3__16_),
	.c(n24472),
	.d(south_input_NIB_storage_data_f_0__16_));
   ao22f01 U27895 (.o(n24474),
	.a(n17782),
	.b(south_input_NIB_storage_data_f_2__16_),
	.c(FE_OFN24741_n18683),
	.d(south_input_NIB_storage_data_f_1__16_));
   ao22f01 U27896 (.o(n24476),
	.a(FE_OFN44_n19054),
	.b(FE_OFN211_n24630),
	.c(FE_OFN366_n17753),
	.d(n24631));
   na02f02 U27897 (.o(n24478),
	.a(n24477),
	.b(n24476));
   ao22f01 U27899 (.o(n24481),
	.a(n19019),
	.b(n24629),
	.c(n19020),
	.d(n24628));
   ao22f01 U27900 (.o(n24480),
	.a(n19017),
	.b(FE_OFN211_n24630),
	.c(FE_OFN42_n19022),
	.d(n24631));
   na02f01 U27901 (.o(n24482),
	.a(n24481),
	.b(n24480));
   ao22f01 U27903 (.o(n24485),
	.a(n19493),
	.b(FE_OFN528_n24732),
	.c(FE_OFN577_n25498),
	.d(FE_OFN237_n24730));
   ao22f01 U27904 (.o(n24484),
	.a(FE_OFN105_n22517),
	.b(n24734),
	.c(FE_OFN93_n21667),
	.d(FE_OFN530_n24733));
   na02f02 U27905 (.o(n24486),
	.a(n24485),
	.b(n24484));
   in01f02 U27906 (.o(n24487),
	.a(n24486));
   ao22f01 U27907 (.o(n24489),
	.a(n19493),
	.b(n24629),
	.c(FE_OFN93_n21667),
	.d(n24628));
   ao22f01 U27908 (.o(n24488),
	.a(FE_OFN105_n22517),
	.b(n24631),
	.c(n25498),
	.d(FE_OFN211_n24630));
   na02f02 U27909 (.o(n24490),
	.a(n24489),
	.b(n24488));
   ao22f01 U27911 (.o(n24493),
	.a(FE_OFN105_n22517),
	.b(n24585),
	.c(FE_OFN93_n21667),
	.d(FE_OFN497_n24586));
   ao22f01 U27912 (.o(n24492),
	.a(n19493),
	.b(n24588),
	.c(n25498),
	.d(n24587));
   na02f02 U27913 (.o(n24494),
	.a(n24493),
	.b(n24492));
   in01s01 U27914 (.o(n24495),
	.a(n24494));
   ao22f01 U27915 (.o(n24497),
	.a(FE_OFN105_n22517),
	.b(n24576),
	.c(FE_OFN93_n21667),
	.d(FE_OFN493_n24577));
   ao22f01 U27916 (.o(n24496),
	.a(n19493),
	.b(FE_OFN495_n24579),
	.c(FE_OFN577_n25498),
	.d(n24578));
   na02f02 U27917 (.o(n24498),
	.a(n24497),
	.b(n24496));
   ao22f01 U27919 (.o(n24501),
	.a(FE_OFN105_n22517),
	.b(n24675),
	.c(FE_OFN93_n21667),
	.d(n24676));
   ao22f01 U27920 (.o(n24500),
	.a(n19493),
	.b(n24678),
	.c(n25498),
	.d(FE_OFN227_n24677));
   na02f02 U27921 (.o(n24502),
	.a(n24501),
	.b(n24500));
   in01s01 U27922 (.o(n24503),
	.a(n24502));
   ao22f01 U27923 (.o(n24505),
	.a(n25498),
	.b(FE_OFN221_n24662),
	.c(FE_OFN93_n21667),
	.d(n24663));
   ao22f01 U27924 (.o(n24504),
	.a(n19493),
	.b(n24665),
	.c(FE_OFN105_n22517),
	.d(FE_OFN223_n24664));
   na02f02 U27925 (.o(n24506),
	.a(n24505),
	.b(n24504));
   in01s01 U27926 (.o(n24507),
	.a(n24506));
   ao22f01 U27927 (.o(n24509),
	.a(n19493),
	.b(n24599),
	.c(FE_OFN105_n22517),
	.d(n24598));
   ao22f01 U27928 (.o(n24508),
	.a(n25498),
	.b(FE_OFN203_n24600),
	.c(FE_OFN93_n21667),
	.d(FE_OFN499_n24601));
   na02f02 U27929 (.o(n24510),
	.a(n24509),
	.b(n24508));
   ao22f01 U27931 (.o(n24513),
	.a(FE_OFN105_n22517),
	.b(n24620),
	.c(n25498),
	.d(FE_OFN207_n24619));
   ao22f01 U27932 (.o(n24512),
	.a(n19493),
	.b(n24622),
	.c(FE_OFN93_n21667),
	.d(n24621));
   na02f02 U27933 (.o(n24514),
	.a(n24513),
	.b(n24512));
   in01s01 U27934 (.o(n24515),
	.a(n24514));
   ao22f01 U27935 (.o(n24517),
	.a(n19493),
	.b(n24685),
	.c(FE_OFN577_n25498),
	.d(FE_OFN229_n24684));
   ao22f01 U27936 (.o(n24516),
	.a(FE_OFN105_n22517),
	.b(n24687),
	.c(FE_OFN93_n21667),
	.d(n24686));
   na02f02 U27937 (.o(n24518),
	.a(n24517),
	.b(n24516));
   ao22f01 U27939 (.o(n24520),
	.a(n19493),
	.b(n24705),
	.c(n25498),
	.d(FE_OFN231_n24704));
   na02f02 U27940 (.o(n24522),
	.a(n24521),
	.b(n24520));
   in01f01 U27941 (.o(n24523),
	.a(n24522));
   ao22f01 U27942 (.o(n24525),
	.a(FE_OFN105_n22517),
	.b(n24638),
	.c(n25498),
	.d(FE_OFN217_n24637));
   ao22f01 U27943 (.o(n24524),
	.a(n19493),
	.b(n24640),
	.c(FE_OFN93_n21667),
	.d(n24639));
   na02f02 U27944 (.o(n24526),
	.a(n24525),
	.b(n24524));
   ao22f01 U27946 (.o(n24529),
	.a(FE_OFN105_n22517),
	.b(n24711),
	.c(FE_OFN93_n21667),
	.d(FE_OFN517_n24712));
   ao22f01 U27947 (.o(n24528),
	.a(n19493),
	.b(n24714),
	.c(FE_OFN577_n25498),
	.d(n24713));
   na02f02 U27948 (.o(n24530),
	.a(n24529),
	.b(n24528));
   ao22f01 U27950 (.o(n24533),
	.a(n19493),
	.b(n24721),
	.c(n25498),
	.d(n24720));
   ao22f01 U27951 (.o(n24532),
	.a(FE_OFN105_n22517),
	.b(n24722),
	.c(FE_OFN93_n21667),
	.d(FE_OFN521_n24723));
   in01s01 U27952 (.o(n24535),
	.a(n24534));
   na02f02 U27953 (.o(n24538),
	.a(n24537),
	.b(n24536));
   in01f01 U27954 (.o(n24539),
	.a(n24538));
   na02f02 U27955 (.o(n24542),
	.a(n24541),
	.b(n24540));
   na02f02 U27957 (.o(n24546),
	.a(n24545),
	.b(n24544));
   na02f02 U27958 (.o(n24550),
	.a(n24549),
	.b(n24548));
   ao22f01 U27960 (.o(n24553),
	.a(FE_OFN105_n22517),
	.b(n24694),
	.c(FE_OFN577_n25498),
	.d(n24693));
   ao22f01 U27961 (.o(n24552),
	.a(n19493),
	.b(n24696),
	.c(FE_OFN93_n21667),
	.d(FE_OFN513_n24695));
   na02f02 U27962 (.o(n24554),
	.a(n24553),
	.b(n24552));
   ao22f01 U27964 (.o(n24556),
	.a(FE_OFN389_n17786),
	.b(FE_OFN495_n24579),
	.c(FE_OFN111_n22773),
	.d(n24578));
   na02f02 U27965 (.o(n24558),
	.a(n24557),
	.b(n24556));
   ao22f01 U27967 (.o(n24561),
	.a(n17786),
	.b(n24721),
	.c(FE_OFN111_n22773),
	.d(n24720));
   na02f01 U27968 (.o(n24562),
	.a(n24561),
	.b(n24560));
   ao22f01 U27970 (.o(n24564),
	.a(n17786),
	.b(n24678),
	.c(FE_OFN111_n22773),
	.d(FE_OFN227_n24677));
   na02f02 U27971 (.o(n24566),
	.a(n24565),
	.b(n24564));
   ao22f01 U27973 (.o(n24568),
	.a(FE_OFN389_n17786),
	.b(n24714),
	.c(FE_OFN111_n22773),
	.d(n24713));
   na02f01 U27974 (.o(n24570),
	.a(n24569),
	.b(n24568));
   ao22f01 U27976 (.o(n24572),
	.a(n17786),
	.b(n24588),
	.c(FE_OFN111_n22773),
	.d(n24587));
   na02f02 U27977 (.o(n24574),
	.a(n24573),
	.b(n24572));
   ao22f01 U27979 (.o(n24581),
	.a(FE_OFN257_n25294),
	.b(FE_OFN493_n24577),
	.c(n17787),
	.d(n24576));
   ao22f01 U27981 (.o(n24590),
	.a(n25294),
	.b(FE_OFN497_n24586),
	.c(n17787),
	.d(n24585));
   in01s01 U27982 (.o(n24592),
	.a(n24591));
   ao22f01 U27983 (.o(n24595),
	.a(n25295),
	.b(n24741),
	.c(n17787),
	.d(n24740));
   in01f01 U27984 (.o(n24597),
	.a(n24596));
   ao22f01 U27985 (.o(n24603),
	.a(n25295),
	.b(n24599),
	.c(n17787),
	.d(n24598));
   in01s01 U27986 (.o(n24605),
	.a(n24604));
   ao22f01 U27987 (.o(n24608),
	.a(n25295),
	.b(n24629),
	.c(n25294),
	.d(n24628));
   ao22f01 U27989 (.o(n24611),
	.a(n25295),
	.b(n24622),
	.c(n25294),
	.d(n24621));
   in01f01 U27990 (.o(n24614),
	.a(n24613));
   ao22f01 U27991 (.o(n24615),
	.a(n25295),
	.b(n24640),
	.c(n25294),
	.d(n24639));
   ao22f01 U27993 (.o(n24623),
	.a(n17786),
	.b(n24622),
	.c(n17755),
	.d(n24621));
   na02f02 U27994 (.o(n24625),
	.a(n24624),
	.b(n24623));
   ao22f01 U27996 (.o(n24633),
	.a(FE_OFN389_n17786),
	.b(n24629),
	.c(n17755),
	.d(n24628));
   na02f02 U27997 (.o(n24634),
	.a(n24633),
	.b(n24632));
   ao22f01 U27999 (.o(n24641),
	.a(FE_OFN389_n17786),
	.b(n24640),
	.c(n17755),
	.d(n24639));
   na02f02 U28000 (.o(n24643),
	.a(n24642),
	.b(n24641));
   ao22f01 U28002 (.o(n24646),
	.a(n25295),
	.b(n24696),
	.c(n25294),
	.d(FE_OFN513_n24695));
   ao22f01 U28004 (.o(n24650),
	.a(FE_OFN257_n25294),
	.b(n24686),
	.c(n17787),
	.d(n24687));
   ao22f01 U28006 (.o(n24655),
	.a(n25294),
	.b(FE_OFN515_n24702),
	.c(n17787),
	.d(n24703));
   in01f01 U28007 (.o(n24657),
	.a(n24656));
   ao22f01 U28008 (.o(n24658),
	.a(FE_OFN257_n25294),
	.b(FE_OFN530_n24733),
	.c(n17787),
	.d(n24734));
   in01f01 U28009 (.o(n24661),
	.a(n24660));
   ao22m02 U28010 (.o(n24666),
	.a(n25295),
	.b(n24665),
	.c(n17787),
	.d(FE_OFN223_n24664));
   in01s01 U28011 (.o(n24669),
	.a(n24668));
   ao22f01 U28012 (.o(n24672),
	.a(n19493),
	.b(FE_OFN546_n24751),
	.c(FE_OFN105_n22517),
	.d(n24750));
   ao22f01 U28013 (.o(n24671),
	.a(FE_OFN577_n25498),
	.b(n24752),
	.c(FE_OFN93_n21667),
	.d(n24754));
   na02f02 U28014 (.o(n24673),
	.a(n24672),
	.b(n24671));
   ao22f01 U28016 (.o(n24680),
	.a(n25294),
	.b(n24676),
	.c(n17787),
	.d(n24675));
   ao22f01 U28017 (.o(n24689),
	.a(FE_OFN389_n17786),
	.b(n24685),
	.c(FE_OFN111_n22773),
	.d(FE_OFN229_n24684));
   na02f02 U28018 (.o(n24690),
	.a(n24689),
	.b(n24688));
   ao22f01 U28020 (.o(n24697),
	.a(FE_OFN389_n17786),
	.b(n24696),
	.c(n17755),
	.d(FE_OFN513_n24695));
   na02f02 U28021 (.o(n24699),
	.a(n24698),
	.b(n24697));
   ao22f01 U28023 (.o(n24706),
	.a(FE_OFN389_n17786),
	.b(n24705),
	.c(FE_OFN111_n22773),
	.d(FE_OFN231_n24704));
   na02f02 U28024 (.o(n24708),
	.a(n24707),
	.b(n24706));
   ao22f01 U28025 (.o(n24716),
	.a(FE_OFN257_n25294),
	.b(FE_OFN517_n24712),
	.c(n17787),
	.d(n24711));
   ao22f01 U28027 (.o(n24724),
	.a(n25294),
	.b(FE_OFN521_n24723),
	.c(n17787),
	.d(n24722));
   ao22f01 U28029 (.o(n24736),
	.a(FE_OFN389_n17786),
	.b(FE_OFN528_n24732),
	.c(FE_OFN111_n22773),
	.d(FE_OFN237_n24730));
   na02f02 U28030 (.o(n24737),
	.a(n24736),
	.b(n24735));
   in01f02 U28031 (.o(n24738),
	.a(n24737));
   ao22f01 U28032 (.o(n24746),
	.a(n19493),
	.b(n24741),
	.c(FE_OFN105_n22517),
	.d(n24740));
   ao22f01 U28033 (.o(n24745),
	.a(FE_OFN577_n25498),
	.b(FE_OFN242_n24744),
	.c(FE_OFN93_n21667),
	.d(n24742));
   na02f02 U28034 (.o(n24747),
	.a(n24746),
	.b(n24745));
   ao22f01 U28036 (.o(n24756),
	.a(n25295),
	.b(FE_OFN546_n24751),
	.c(n17787),
	.d(n24750));
   in01s01 U28039 (.o(n24763),
	.a(east_input_NIB_storage_data_f_1__61_));
   na02s01 U28040 (.o(n24762),
	.a(dataIn_E_61_),
	.b(FE_OFN555_n24761));
   oa12s01 U28041 (.o(n11143),
	.a(n24762),
	.b(FE_OFN555_n24761),
	.c(n24763));
   na02s01 U28042 (.o(n24764),
	.a(dataIn_E_62_),
	.b(FE_OFN555_n24761));
   na02s01 U28043 (.o(n24766),
	.a(dataIn_E_60_),
	.b(FE_OFN555_n24761));
   oa12s01 U28044 (.o(n11148),
	.a(n24766),
	.b(FE_OFN555_n24761),
	.c(n24767));
   in01s01 U28045 (.o(n24769),
	.a(east_input_NIB_storage_data_f_1__56_));
   na02s01 U28046 (.o(n24768),
	.a(dataIn_E_56_),
	.b(FE_OFN555_n24761));
   oa12s01 U28047 (.o(n11168),
	.a(n24768),
	.b(FE_OFN555_n24761),
	.c(n24769));
   na02s01 U28048 (.o(n24770),
	.a(dataIn_E_58_),
	.b(FE_OFN555_n24761));
   oa12s01 U28049 (.o(n11158),
	.a(n24770),
	.b(FE_OFN555_n24761),
	.c(n24771));
   in01s01 U28050 (.o(n24773),
	.a(east_input_NIB_storage_data_f_1__52_));
   na02s01 U28051 (.o(n24772),
	.a(dataIn_E_52_),
	.b(FE_OFN555_n24761));
   oa12s01 U28052 (.o(n11188),
	.a(n24772),
	.b(FE_OFN555_n24761),
	.c(n24773));
   in01s01 U28053 (.o(n24775),
	.a(east_input_NIB_storage_data_f_1__63_));
   na02s01 U28054 (.o(n24774),
	.a(dataIn_E_63_),
	.b(FE_OFN555_n24761));
   oa12s01 U28055 (.o(n11133),
	.a(n24774),
	.b(FE_OFN555_n24761),
	.c(n24775));
   na02s01 U28056 (.o(n24776),
	.a(dataIn_E_41_),
	.b(n24761));
   oa12s01 U28057 (.o(n11243),
	.a(n24776),
	.b(n24761),
	.c(n24777));
   in01s01 U28058 (.o(n24779),
	.a(east_input_NIB_storage_data_f_1__51_));
   na02s01 U28059 (.o(n24778),
	.a(dataIn_E_51_),
	.b(FE_OFN555_n24761));
   oa12s01 U28060 (.o(n11193),
	.a(n24778),
	.b(FE_OFN555_n24761),
	.c(n24779));
   in01s01 U28061 (.o(n24781),
	.a(east_input_NIB_storage_data_f_1__59_));
   na02s01 U28062 (.o(n24780),
	.a(dataIn_E_59_),
	.b(FE_OFN555_n24761));
   oa12s01 U28063 (.o(n11153),
	.a(n24780),
	.b(FE_OFN555_n24761),
	.c(n24781));
   na02s01 U28064 (.o(n24782),
	.a(dataIn_E_54_),
	.b(FE_OFN555_n24761));
   na02s01 U28065 (.o(n24784),
	.a(dataIn_E_57_),
	.b(FE_OFN555_n24761));
   oa12s01 U28066 (.o(n11163),
	.a(n24784),
	.b(FE_OFN555_n24761),
	.c(n24785));
   na02s01 U28067 (.o(n24786),
	.a(dataIn_E_30_),
	.b(n24761));
   oa12s01 U28068 (.o(n11298),
	.a(n24786),
	.b(n24761),
	.c(n24787));
   in01s01 U28069 (.o(n24789),
	.a(east_input_NIB_storage_data_f_1__55_));
   na02s01 U28070 (.o(n24788),
	.a(dataIn_E_55_),
	.b(FE_OFN555_n24761));
   oa12s01 U28071 (.o(n11173),
	.a(n24788),
	.b(FE_OFN555_n24761),
	.c(n24789));
   in01s01 U28072 (.o(n24791),
	.a(east_input_NIB_storage_data_f_1__50_));
   oa12s01 U28073 (.o(n11198),
	.a(n24790),
	.b(FE_OFN555_n24761),
	.c(n24791));
   na02s01 U28074 (.o(n24792),
	.a(dataIn_E_53_),
	.b(FE_OFN555_n24761));
   oa12s01 U28075 (.o(n11183),
	.a(n24792),
	.b(FE_OFN555_n24761),
	.c(n24793));
   oa22s01 U28076 (.o(n24794),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_17_),
	.c(south_input_NIB_storage_data_f_0__17_),
	.d(FE_OFN83_n20814));
   in01s01 U28077 (.o(n9753),
	.a(n24794));
   oa22s01 U28078 (.o(n24795),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_21_),
	.c(south_input_NIB_storage_data_f_0__21_),
	.d(FE_OFN83_n20814));
   in01s01 U28079 (.o(n9733),
	.a(n24795));
   oa22s01 U28080 (.o(n24796),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_18_),
	.c(south_input_NIB_storage_data_f_0__18_),
	.d(FE_OFN83_n20814));
   in01s01 U28081 (.o(n9748),
	.a(n24796));
   oa22s01 U28082 (.o(n24797),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_13_),
	.c(south_input_NIB_storage_data_f_0__13_),
	.d(FE_OFN83_n20814));
   in01s01 U28083 (.o(n9773),
	.a(n24797));
   oa22s01 U28084 (.o(n24798),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_19_),
	.c(south_input_NIB_storage_data_f_0__19_),
	.d(FE_OFN83_n20814));
   in01s01 U28085 (.o(n9743),
	.a(n24798));
   oa22s01 U28086 (.o(n24799),
	.a(FE_OFN952_n25916),
	.b(dataIn_S_16_),
	.c(south_input_NIB_storage_data_f_0__16_),
	.d(FE_OFN83_n20814));
   in01s01 U28087 (.o(n9758),
	.a(n24799));
   in01s01 U28088 (.o(n9768),
	.a(n24800));
   oa22m01 U28089 (.o(n24801),
	.a(FE_OFN25749_FE_OFN24796_n20854),
	.b(dataIn_W_14_),
	.c(west_input_NIB_storage_data_f_0__14_),
	.d(n20855));
   in01s01 U28090 (.o(n8478),
	.a(n24801));
   oa22m01 U28091 (.o(n24802),
	.a(FE_OFN25750_FE_OFN24796_n20854),
	.b(dataIn_W_18_),
	.c(west_input_NIB_storage_data_f_0__18_),
	.d(n20855));
   in01s01 U28092 (.o(n8458),
	.a(n24802));
   oa22m01 U28093 (.o(n24803),
	.a(FE_OFN25749_FE_OFN24796_n20854),
	.b(dataIn_W_12_),
	.c(west_input_NIB_storage_data_f_0__12_),
	.d(n20855));
   in01s01 U28094 (.o(n8488),
	.a(n24803));
   oa22m01 U28095 (.o(n24804),
	.a(FE_OFN25749_FE_OFN24796_n20854),
	.b(dataIn_W_15_),
	.c(west_input_NIB_storage_data_f_0__15_),
	.d(n20855));
   in01s01 U28096 (.o(n8473),
	.a(n24804));
   oa22m01 U28097 (.o(n24805),
	.a(FE_OFN25750_FE_OFN24796_n20854),
	.b(dataIn_W_16_),
	.c(west_input_NIB_storage_data_f_0__16_),
	.d(n20855));
   in01s01 U28098 (.o(n8468),
	.a(n24805));
   oa22m01 U28099 (.o(n24806),
	.a(FE_OFN25749_FE_OFN24796_n20854),
	.b(dataIn_W_20_),
	.c(west_input_NIB_storage_data_f_0__20_),
	.d(n20855));
   in01s01 U28100 (.o(n8448),
	.a(n24806));
   oa22s01 U28101 (.o(n24807),
	.a(FE_OFN1102_n25965),
	.b(dataIn_W_19_),
	.c(west_input_NIB_storage_data_f_0__19_),
	.d(n20855));
   in01s01 U28102 (.o(n8453),
	.a(n24807));
   oa22s01 U28103 (.o(n24808),
	.a(FE_OFN24794_n20854),
	.b(dataIn_W_33_),
	.c(west_input_NIB_storage_data_f_0__33_),
	.d(n20855));
   in01s01 U28104 (.o(n8383),
	.a(n24808));
   oa22m01 U28105 (.o(n24809),
	.a(FE_OFN25749_FE_OFN24796_n20854),
	.b(dataIn_W_21_),
	.c(west_input_NIB_storage_data_f_0__21_),
	.d(n20855));
   oa22s01 U28106 (.o(n24810),
	.a(FE_OFN1090_n20855),
	.b(dataIn_W_13_),
	.c(west_input_NIB_storage_data_f_0__13_),
	.d(n20855));
   in01s01 U28107 (.o(n8483),
	.a(n24810));
   oa22s01 U28108 (.o(n24811),
	.a(FE_OFN25785_n17770),
	.b(dataIn_S_19_),
	.c(south_input_NIB_storage_data_f_1__19_),
	.d(n20797));
   in01s01 U28109 (.o(n10063),
	.a(n24811));
   oa22s01 U28110 (.o(n24812),
	.a(n17770),
	.b(dataIn_S_16_),
	.c(south_input_NIB_storage_data_f_1__16_),
	.d(n20797));
   in01s01 U28111 (.o(n10078),
	.a(n24812));
   oa22f01 U28112 (.o(n24813),
	.a(FE_OFN25787_n17770),
	.b(dataIn_S_13_),
	.c(south_input_NIB_storage_data_f_1__13_),
	.d(n20797));
   oa22s01 U28113 (.o(n24814),
	.a(n17770),
	.b(dataIn_S_18_),
	.c(south_input_NIB_storage_data_f_1__18_),
	.d(n20797));
   in01s01 U28114 (.o(n10068),
	.a(n24814));
   in01s01 U28115 (.o(n10053),
	.a(n24815));
   oa22s01 U28116 (.o(n24816),
	.a(FE_OFN25785_n17770),
	.b(dataIn_S_17_),
	.c(south_input_NIB_storage_data_f_1__17_),
	.d(n20797));
   in01s01 U28117 (.o(n10073),
	.a(n24816));
   oa22s01 U28118 (.o(n24817),
	.a(n17770),
	.b(dataIn_S_11_),
	.c(south_input_NIB_storage_data_f_1__11_),
	.d(n20797));
   in01s01 U28119 (.o(n10103),
	.a(n24817));
   oa22s01 U28120 (.o(n24818),
	.a(FE_OFN25785_n17770),
	.b(dataIn_S_14_),
	.c(south_input_NIB_storage_data_f_1__14_),
	.d(n20797));
   in01s01 U28121 (.o(n10088),
	.a(n24818));
   oa22m01 U28122 (.o(n24819),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_33_),
	.c(west_input_NIB_storage_data_f_1__33_),
	.d(FE_OFN380_n17772));
   in01s01 U28123 (.o(n8703),
	.a(n24819));
   oa22m01 U28124 (.o(n24820),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_13_),
	.c(west_input_NIB_storage_data_f_1__13_),
	.d(FE_OFN380_n17772));
   in01s01 U28125 (.o(n8803),
	.a(n24820));
   oa22m01 U28126 (.o(n24821),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_21_),
	.c(west_input_NIB_storage_data_f_1__21_),
	.d(FE_OFN380_n17772));
   in01s01 U28127 (.o(n8763),
	.a(n24821));
   oa22m01 U28128 (.o(n24822),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_18_),
	.c(west_input_NIB_storage_data_f_1__18_),
	.d(FE_OFN380_n17772));
   in01s01 U28129 (.o(n8778),
	.a(n24822));
   oa22m01 U28130 (.o(n24823),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_15_),
	.c(west_input_NIB_storage_data_f_1__15_),
	.d(FE_OFN380_n17772));
   in01s01 U28131 (.o(n8793),
	.a(n24823));
   oa22m01 U28132 (.o(n24824),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_12_),
	.c(west_input_NIB_storage_data_f_1__12_),
	.d(FE_OFN380_n17772));
   in01s01 U28133 (.o(n8808),
	.a(n24824));
   oa22m01 U28134 (.o(n24825),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_20_),
	.c(west_input_NIB_storage_data_f_1__20_),
	.d(FE_OFN380_n17772));
   in01s01 U28135 (.o(n8768),
	.a(n24825));
   oa22m01 U28136 (.o(n24826),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_19_),
	.c(west_input_NIB_storage_data_f_1__19_),
	.d(FE_OFN380_n17772));
   in01s01 U28137 (.o(n8773),
	.a(n24826));
   oa22m01 U28138 (.o(n24827),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_16_),
	.c(west_input_NIB_storage_data_f_1__16_),
	.d(FE_OFN380_n17772));
   in01s01 U28139 (.o(n8788),
	.a(n24827));
   oa22m01 U28140 (.o(n24828),
	.a(FE_OFN382_n17772),
	.b(dataIn_W_14_),
	.c(west_input_NIB_storage_data_f_1__14_),
	.d(FE_OFN380_n17772));
   in01s01 U28141 (.o(n8798),
	.a(n24828));
   in01s01 U28142 (.o(n12358),
	.a(n24829));
   in01s01 U28143 (.o(n12338),
	.a(n24830));
   in01s01 U28144 (.o(n12348),
	.a(n24831));
   in01s01 U28145 (.o(n12253),
	.a(n24833));
   in01s01 U28146 (.o(n12333),
	.a(n24834));
   in01s01 U28147 (.o(n12318),
	.a(n24835));
   oa22f01 U28148 (.o(n24836),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_17_),
	.c(south_input_NIB_storage_data_f_2__17_),
	.d(n20972));
   in01s01 U28149 (.o(n10718),
	.a(n24837));
   in01s01 U28150 (.o(n10703),
	.a(n24838));
   oa22f01 U28151 (.o(n24839),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_14_),
	.c(south_input_NIB_storage_data_f_2__14_),
	.d(n20972));
   in01s01 U28152 (.o(n10408),
	.a(n24839));
   oa22f01 U28153 (.o(n24840),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_19_),
	.c(south_input_NIB_storage_data_f_2__19_),
	.d(n20972));
   in01s01 U28154 (.o(n10383),
	.a(n24840));
   in01s01 U28155 (.o(n10733),
	.a(n24841));
   in01s01 U28156 (.o(n10713),
	.a(n24842));
   oa22f01 U28157 (.o(n24843),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_16_),
	.c(south_input_NIB_storage_data_f_2__16_),
	.d(n20972));
   in01s01 U28158 (.o(n10398),
	.a(n24843));
   in01s01 U28159 (.o(n10728),
	.a(n24844));
   oa22f01 U28160 (.o(n24845),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_18_),
	.c(south_input_NIB_storage_data_f_2__18_),
	.d(n20972));
   in01s01 U28161 (.o(n10388),
	.a(n24845));
   in01s01 U28162 (.o(n10373),
	.a(n24846));
   in01s01 U28163 (.o(n10708),
	.a(n24848));
   oa22f01 U28164 (.o(n24849),
	.a(FE_OFN84_n20972),
	.b(dataIn_S_13_),
	.c(south_input_NIB_storage_data_f_2__13_),
	.d(n20972));
   in01s01 U28165 (.o(n10413),
	.a(n24849));
   in01s01 U28166 (.o(n9443),
	.a(n24850));
   in01s01 U28167 (.o(n9088),
	.a(n24851));
   oa22f01 U28168 (.o(n24852),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_33_),
	.c(west_input_NIB_storage_data_f_2__33_),
	.d(n25945));
   in01s01 U28169 (.o(n9023),
	.a(n24852));
   oa22f01 U28170 (.o(n24853),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_14_),
	.c(west_input_NIB_storage_data_f_2__14_),
	.d(n25945));
   oa22f01 U28171 (.o(n24854),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_18_),
	.c(west_input_NIB_storage_data_f_2__18_),
	.d(n25945));
   in01s01 U28172 (.o(n9098),
	.a(n24854));
   oa22f01 U28173 (.o(n24855),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_12_),
	.c(west_input_NIB_storage_data_f_2__12_),
	.d(n25945));
   in01s01 U28174 (.o(n9128),
	.a(n24855));
   oa22f01 U28175 (.o(n24856),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_14_),
	.c(west_input_NIB_storage_data_f_3__14_),
	.d(n21070));
   in01s01 U28176 (.o(n9438),
	.a(n24856));
   oa22f01 U28177 (.o(n24857),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_19_),
	.c(west_input_NIB_storage_data_f_3__19_),
	.d(n21070));
   in01s01 U28178 (.o(n9413),
	.a(n24857));
   oa22f01 U28179 (.o(n24858),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_16_),
	.c(west_input_NIB_storage_data_f_2__16_),
	.d(n25945));
   in01s01 U28180 (.o(n9108),
	.a(n24858));
   oa22f01 U28181 (.o(n24859),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_20_),
	.c(west_input_NIB_storage_data_f_3__20_),
	.d(n21070));
   in01s01 U28182 (.o(n9408),
	.a(n24859));
   in01s01 U28183 (.o(n9403),
	.a(n24860));
   oa22f01 U28184 (.o(n24861),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_12_),
	.c(west_input_NIB_storage_data_f_3__12_),
	.d(n21070));
   in01s01 U28185 (.o(n9448),
	.a(n24861));
   oa22f01 U28186 (.o(n24862),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_15_),
	.c(west_input_NIB_storage_data_f_3__15_),
	.d(n21070));
   in01s01 U28187 (.o(n9433),
	.a(n24862));
   oa22f01 U28188 (.o(n24863),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_16_),
	.c(west_input_NIB_storage_data_f_3__16_),
	.d(n21070));
   in01s01 U28189 (.o(n9428),
	.a(n24863));
   oa22f01 U28190 (.o(n24864),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_21_),
	.c(west_input_NIB_storage_data_f_2__21_),
	.d(n25945));
   in01s01 U28191 (.o(n9083),
	.a(n24864));
   oa22f01 U28192 (.o(n24865),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_15_),
	.c(west_input_NIB_storage_data_f_2__15_),
	.d(n25945));
   in01s01 U28193 (.o(n9113),
	.a(n24865));
   oa22f01 U28194 (.o(n24866),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_19_),
	.c(west_input_NIB_storage_data_f_2__19_),
	.d(n25945));
   in01s01 U28195 (.o(n9093),
	.a(n24866));
   oa22f01 U28196 (.o(n24867),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_18_),
	.c(west_input_NIB_storage_data_f_3__18_),
	.d(n21070));
   oa22f01 U28197 (.o(n24868),
	.a(FE_OFN24767_n21069),
	.b(dataIn_W_33_),
	.c(west_input_NIB_storage_data_f_3__33_),
	.d(n21070));
   oa22f01 U28198 (.o(n24869),
	.a(FE_OFN25791_n21053),
	.b(dataIn_W_13_),
	.c(west_input_NIB_storage_data_f_2__13_),
	.d(n25945));
   in01s01 U28199 (.o(n9123),
	.a(n24869));
   in01s01 U28200 (.o(n24871),
	.a(east_input_NIB_storage_data_f_1__28_));
   na02s01 U28201 (.o(n24870),
	.a(dataIn_E_28_),
	.b(n24761));
   in01s01 U28202 (.o(n24873),
	.a(east_input_NIB_storage_data_f_1__22_));
   na02s01 U28203 (.o(n24872),
	.a(dataIn_E_22_),
	.b(n24761));
   in01s01 U28204 (.o(n24875),
	.a(east_input_NIB_storage_data_f_1__23_));
   na02s01 U28205 (.o(n24874),
	.a(dataIn_E_23_),
	.b(n24761));
   in01s01 U28206 (.o(n24877),
	.a(east_input_NIB_storage_data_f_1__24_));
   na02s01 U28207 (.o(n24876),
	.a(dataIn_E_24_),
	.b(n24761));
   in01s01 U28208 (.o(n24879),
	.a(east_input_NIB_storage_data_f_1__25_));
   na02s01 U28209 (.o(n24878),
	.a(dataIn_E_25_),
	.b(FE_OFN555_n24761));
   in01s01 U28210 (.o(n24881),
	.a(east_input_NIB_storage_data_f_1__26_));
   na02s01 U28211 (.o(n24880),
	.a(dataIn_E_26_),
	.b(n24761));
   in01s01 U28212 (.o(n24883),
	.a(east_input_NIB_storage_data_f_1__27_));
   oa12s01 U28213 (.o(n11313),
	.a(n24882),
	.b(FE_OFN555_n24761),
	.c(n24883));
   in01s01 U28214 (.o(n24885),
	.a(east_input_NIB_storage_data_f_1__29_));
   na02s01 U28215 (.o(n24884),
	.a(dataIn_E_29_),
	.b(n24761));
   na02s01 U28216 (.o(n24886),
	.a(dataIn_E_32_),
	.b(n24761));
   in01s01 U28217 (.o(n24889),
	.a(east_input_NIB_storage_data_f_1__31_));
   na02s01 U28218 (.o(n24888),
	.a(dataIn_E_31_),
	.b(n24761));
   oa12s01 U28219 (.o(n11293),
	.a(n24888),
	.b(n24761),
	.c(n24889));
   na02s01 U28220 (.o(n24890),
	.a(dataIn_E_40_),
	.b(n24761));
   oa12s01 U28221 (.o(n11248),
	.a(n24890),
	.b(n24761),
	.c(n24891));
   na02s01 U28222 (.o(n24892),
	.a(dataIn_E_34_),
	.b(n24761));
   oa12s01 U28223 (.o(n11278),
	.a(n24892),
	.b(n24761),
	.c(n24893));
   na02s01 U28224 (.o(n24894),
	.a(dataIn_E_43_),
	.b(n24761));
   oa12s01 U28225 (.o(n11233),
	.a(n24894),
	.b(n24761),
	.c(n24895));
   in01s01 U28226 (.o(n24897),
	.a(east_input_NIB_storage_data_f_1__44_));
   na02s01 U28227 (.o(n24896),
	.a(dataIn_E_44_),
	.b(n24761));
   oa12s01 U28228 (.o(n11228),
	.a(n24896),
	.b(n24761),
	.c(n24897));
   in01s01 U28229 (.o(n24899),
	.a(east_input_NIB_storage_data_f_1__35_));
   oa12s01 U28230 (.o(n11273),
	.a(n24898),
	.b(n24761),
	.c(n24899));
   in01s01 U28231 (.o(n24901),
	.a(east_input_NIB_storage_data_f_1__36_));
   na02s01 U28232 (.o(n24900),
	.a(dataIn_E_36_),
	.b(n24761));
   oa12s01 U28233 (.o(n11268),
	.a(n24900),
	.b(n24761),
	.c(n24901));
   in01s01 U28234 (.o(n24903),
	.a(east_input_NIB_storage_data_f_1__37_));
   na02s01 U28235 (.o(n24902),
	.a(dataIn_E_37_),
	.b(n24761));
   oa12s01 U28236 (.o(n11263),
	.a(n24902),
	.b(n24761),
	.c(n24903));
   na02s01 U28237 (.o(n24904),
	.a(dataIn_E_38_),
	.b(n24761));
   oa12s01 U28238 (.o(n11258),
	.a(n24904),
	.b(n24761),
	.c(n24905));
   na02s01 U28239 (.o(n24906),
	.a(dataIn_E_39_),
	.b(n24761));
   oa12s01 U28240 (.o(n11253),
	.a(n24906),
	.b(n24761),
	.c(n24907));
   na02s01 U28241 (.o(n24908),
	.a(dataIn_E_48_),
	.b(n24761));
   oa12s01 U28242 (.o(n11208),
	.a(n24908),
	.b(n24761),
	.c(n24909));
   na02s01 U28243 (.o(n24910),
	.a(dataIn_E_42_),
	.b(n24761));
   oa12s01 U28244 (.o(n11238),
	.a(n24910),
	.b(n24761),
	.c(n24911));
   in01s01 U28245 (.o(n24913),
	.a(east_input_NIB_storage_data_f_1__47_));
   na02s01 U28246 (.o(n24912),
	.a(dataIn_E_47_),
	.b(n24761));
   oa12s01 U28247 (.o(n11213),
	.a(n24912),
	.b(n24761),
	.c(n24913));
   in01s01 U28248 (.o(n24915),
	.a(east_input_NIB_storage_data_f_1__45_));
   na02s01 U28249 (.o(n24914),
	.a(dataIn_E_45_),
	.b(n24761));
   oa12s01 U28250 (.o(n11223),
	.a(n24914),
	.b(n24761),
	.c(n24915));
   in01s01 U28251 (.o(n24917),
	.a(east_input_NIB_storage_data_f_1__46_));
   na02s01 U28252 (.o(n24916),
	.a(dataIn_E_46_),
	.b(n24761));
   oa12s01 U28253 (.o(n11218),
	.a(n24916),
	.b(n24761),
	.c(n24917));
   na02s01 U28254 (.o(n24918),
	.a(dataIn_E_49_),
	.b(n24761));
   oa12s01 U28255 (.o(n11203),
	.a(n24918),
	.b(n24761),
	.c(n24919));
   na02f01 U28256 (.o(n24922),
	.a(east_input_NIB_storage_data_f_3__43_),
	.b(n24921));
   na02s01 U28257 (.o(n24924),
	.a(east_input_NIB_storage_data_f_3__34_),
	.b(n24921));
   na02s01 U28258 (.o(n24926),
	.a(east_input_NIB_storage_data_f_3__48_),
	.b(n24921));
   na02s01 U28259 (.o(n24928),
	.a(east_input_NIB_storage_data_f_3__38_),
	.b(n24921));
   na02s01 U28260 (.o(n24930),
	.a(east_input_NIB_storage_data_f_3__40_),
	.b(n24921));
   na02s01 U28261 (.o(n24932),
	.a(east_input_NIB_storage_data_f_3__39_),
	.b(n24921));
   na02s01 U28262 (.o(n24934),
	.a(east_input_NIB_storage_data_f_3__49_),
	.b(n24921));
   na02s01 U28263 (.o(n24936),
	.a(east_input_NIB_storage_data_f_3__42_),
	.b(n24921));
   na02s01 U28264 (.o(n24938),
	.a(east_input_NIB_storage_data_f_3__35_),
	.b(n24921));
   na02s01 U28265 (.o(n24940),
	.a(east_input_NIB_storage_data_f_3__37_),
	.b(n24921));
   na02s01 U28266 (.o(n24942),
	.a(east_input_NIB_storage_data_f_3__36_),
	.b(n24921));
   na02s01 U28267 (.o(n24944),
	.a(east_input_NIB_storage_data_f_3__45_),
	.b(n24921));
   na02s01 U28268 (.o(n24946),
	.a(east_input_NIB_storage_data_f_3__44_),
	.b(n24921));
   na02s01 U28269 (.o(n24948),
	.a(east_input_NIB_storage_data_f_3__47_),
	.b(n24921));
   na02s01 U28270 (.o(n24950),
	.a(east_input_NIB_storage_data_f_3__46_),
	.b(n24921));
   in01m01 U28271 (.o(n24961),
	.a(south_output_current_route_connection_2_));
   oa22f02 U28272 (.o(south_output_control_N469),
	.a(n24963),
	.b(n24962),
	.c(n24961),
	.d(n24988));
   na02f01 U28273 (.o(n24967),
	.a(south_input_NIB_head_ptr_f_1_),
	.b(n25433));
   no02f04 U28274 (.o(n24985),
	.a(n24982),
	.b(n24981));
   oa22f02 U28275 (.o(south_output_control_N468),
	.a(n24991),
	.b(n24990),
	.c(n24989),
	.d(n24988));
   in01s01 U28276 (.o(n24994),
	.a(n25005));
   no04f04 U28277 (.o(n25016),
	.a(n25408),
	.b(n17757),
	.c(n20501),
	.d(n25055));
   na03m02 U28278 (.o(n25004),
	.a(n25003),
	.b(n25002),
	.c(n25001));
   oa22f02 U28279 (.o(n25015),
	.a(n25014),
	.b(n25013),
	.c(n25409),
	.d(n25012));
   ao12f02 U28280 (.o(n25039),
	.a(n25015),
	.b(n25016),
	.c(n25049));
   oa22f02 U28281 (.o(proc_output_control_N468),
	.a(n25039),
	.b(n25423),
	.c(n25038),
	.d(n25421));
   na02f01 U28282 (.o(n25472),
	.a(proc_input_NIB_elements_in_array_f_0_),
	.b(proc_input_NIB_elements_in_array_f_1_));
   no02s01 U28283 (.o(n25040),
	.a(n25974),
	.b(n25472));
   no04f01 U28284 (.o(n25042),
	.a(reset),
	.b(proc_input_NIB_elements_in_array_f_2_),
	.c(n18408),
	.d(n25041));
   na02s01 U28285 (.o(n25464),
	.a(n25979),
	.b(n25472));
   na02f01 U28286 (.o(n25043),
	.a(n25974),
	.b(proc_input_NIB_elements_in_array_f_1_));
   na03s01 U28287 (.o(n25045),
	.a(n25044),
	.b(n25464),
	.c(n25043));
   na02f01 U28288 (.o(n25047),
	.a(proc_input_NIB_elements_in_array_f_2_),
	.b(n25045));
   in01f02 U28289 (.o(n25059),
	.a(n25049));
   in01m01 U28290 (.o(n25407),
	.a(n25050));
   ao12f02 U28291 (.o(n25056),
	.a(proc_output_current_route_connection_2_),
	.b(n25054),
	.c(n25053));
   na02f02 U28292 (.o(n25057),
	.a(n25056),
	.b(n25055));
   ao22f02 U28293 (.o(n25058),
	.a(n25414),
	.b(n20501),
	.c(n25407),
	.d(n25057));
   oa22f02 U28294 (.o(proc_output_control_N469),
	.a(n25061),
	.b(n25421),
	.c(n25423),
	.d(n25060));
   no03f02 U28295 (.o(n25067),
	.a(east_output_current_route_connection_2_),
	.b(n25063),
	.c(n25387));
   in01s01 U28296 (.o(n25064),
	.a(east_output_current_route_connection_1_));
   na02f01 U28297 (.o(n25076),
	.a(west_input_NIB_head_ptr_f_1_),
	.b(n25463));
   in01s01 U28298 (.o(n25089),
	.a(north_output_control_planned_f));
   na03f04 U28299 (.o(n25100),
	.a(n25101),
	.b(n25102),
	.c(n25093));
   ao12f02 U28300 (.o(n25108),
	.a(n25099),
	.b(n25105),
	.c(n25100));
   in01f02 U28302 (.o(n25103),
	.a(n25102));
   no03f02 U28304 (.o(north_output_control_N470),
	.a(FE_OFN5_reset),
	.b(n25108),
	.c(n25107));
   no02f03 U28305 (.o(n25122),
	.a(n25119),
	.b(n25118));
   no02f01 U28306 (.o(n25121),
	.a(FE_OFN255_n25247),
	.b(FE_OFN563_n25120));
   no04f04 U28307 (.o(n25125),
	.a(n25123),
	.b(n19057),
	.c(n25122),
	.d(n25121));
   no02f02 U28308 (.o(n25136),
	.a(n25125),
	.b(n25124));
   na02f02 U28309 (.o(n2868),
	.a(n25144),
	.b(n25143));
   na02f01 U28310 (.o(n25148),
	.a(east_input_NIB_head_ptr_f_0_),
	.b(FE_OFN25596_reset));
   no02f01 U28311 (.o(n25145),
	.a(FE_OFN25600_reset),
	.b(east_input_NIB_head_ptr_f_0_));
   na02f02 U28312 (.o(n2858),
	.a(n25151),
	.b(n25150));
   na02s01 U28313 (.o(n25167),
	.a(west_output_current_route_connection_2_),
	.b(FE_OFN575_n25463));
   in01s01 U28314 (.o(n25157),
	.a(n25156));
   na02s01 U28315 (.o(n25164),
	.a(n25163),
	.b(n25162));
   no02f02 U28316 (.o(n25166),
	.a(n25184),
	.b(n25165));
   in01s01 U28318 (.o(n25171),
	.a(n25168));
   in01f02 U28319 (.o(n25185),
	.a(n25184));
   in01s01 U28320 (.o(n12363),
	.a(n25188));
   na02s01 U28321 (.o(n25189),
	.a(east_input_NIB_storage_data_f_3__41_),
	.b(n24921));
   na02s01 U28322 (.o(n25191),
	.a(east_input_NIB_storage_data_f_3__59_),
	.b(FE_OFN943_n24921));
   na02s01 U28323 (.o(n25193),
	.a(east_input_NIB_storage_data_f_3__58_),
	.b(FE_OFN943_n24921));
   na02s01 U28324 (.o(n25197),
	.a(east_input_NIB_storage_data_f_3__63_),
	.b(FE_OFN943_n24921));
   na02s01 U28325 (.o(n25199),
	.a(east_input_NIB_storage_data_f_3__52_),
	.b(FE_OFN943_n24921));
   na02s01 U28326 (.o(n25207),
	.a(east_input_NIB_storage_data_f_3__61_),
	.b(FE_OFN943_n24921));
   na02s01 U28327 (.o(n25211),
	.a(east_input_NIB_storage_data_f_3__50_),
	.b(FE_OFN943_n24921));
   na02s01 U28328 (.o(n25213),
	.a(east_input_NIB_storage_data_f_3__51_),
	.b(FE_OFN943_n24921));
   na02s01 U28329 (.o(n25215),
	.a(east_input_NIB_storage_data_f_3__56_),
	.b(FE_OFN943_n24921));
   na02s01 U28330 (.o(n25219),
	.a(east_input_NIB_storage_data_f_3__30_),
	.b(n24921));
   na02s01 U28331 (.o(n25223),
	.a(east_input_NIB_storage_data_f_3__31_),
	.b(n24921));
   na02f01 U28332 (.o(n25228),
	.a(n25227),
	.b(n25225));
   no02s01 U28333 (.o(n25226),
	.a(west_input_control_count_f_6_),
	.b(west_input_control_count_f_7_));
   ao22s01 U28334 (.o(n25235),
	.a(west_input_NIB_elements_in_array_f_0_),
	.b(n25929),
	.c(validIn_W),
	.d(n25234));
   in01s01 U28335 (.o(n25251),
	.a(n26026));
   in01s01 U28336 (.o(n25249),
	.a(n25239));
   no03s01 U28337 (.o(n25243),
	.a(south_input_control_count_f_6_),
	.b(south_input_control_count_f_1_),
	.c(n25242));
   in01s01 U28338 (.o(n25244),
	.a(n25243));
   no02f01 U28340 (.o(south_input_control_N52),
	.a(n25251),
	.b(n25462));
   na02s01 U28341 (.o(n25252),
	.a(east_input_NIB_storage_data_f_3__22_),
	.b(n24921));
   na02s01 U28342 (.o(n25256),
	.a(east_input_NIB_storage_data_f_3__26_),
	.b(n24921));
   na02s01 U28343 (.o(n25262),
	.a(east_input_NIB_storage_data_f_3__25_),
	.b(n24921));
   na02s01 U28344 (.o(n25264),
	.a(east_input_NIB_storage_data_f_3__27_),
	.b(n24921));
   ao22s01 U28345 (.o(n25270),
	.a(south_input_NIB_elements_in_array_f_0_),
	.b(n25897),
	.c(validIn_S),
	.d(n25268));
   in01s01 U28346 (.o(n25269),
	.a(n25270));
   in01f01 U28347 (.o(south_output_space_N46),
	.a(n25273));
   na02s01 U28348 (.o(n25281),
	.a(validIn_N),
	.b(north_input_NIB_elements_in_array_f_0_));
   no02s01 U28349 (.o(n25279),
	.a(north_input_NIB_elements_in_array_f_0_),
	.b(validIn_N));
   ao22s01 U28350 (.o(n25274),
	.a(north_input_NIB_elements_in_array_f_0_),
	.b(validIn_N),
	.c(n25830),
	.d(n25289));
   na02s01 U28351 (.o(n25283),
	.a(north_input_NIB_elements_in_array_f_2_),
	.b(n17888));
   in01s01 U28352 (.o(n25284),
	.a(n25281));
   na02s01 U28353 (.o(n25282),
	.a(north_input_NIB_elements_in_array_f_2_),
	.b(n25288));
   oa22s01 U28354 (.o(n25285),
	.a(n25284),
	.b(n25283),
	.c(n25282),
	.d(n25287));
   na02s01 U28355 (.o(n25297),
	.a(n25294),
	.b(proc_output_control_planned_f));
   na02s01 U28356 (.o(n25296),
	.a(FE_OFN259_n25295),
	.b(proc_output_control_planned_f));
   ao22f02 U28357 (.o(n25298),
	.a(n25412),
	.b(n25297),
	.c(n17757),
	.d(n25296));
   na02s01 U28358 (.o(n25299),
	.a(FE_OFN79_n20501),
	.b(proc_output_control_planned_f));
   na02f04 U28359 (.o(n25304),
	.a(n25303),
	.b(n25302));
   na02f04 U28360 (.o(n25306),
	.a(n25305),
	.b(n25304));
   no02f04 U28361 (.o(n25314),
	.a(n25307),
	.b(n25306));
   no02m02 U28362 (.o(n25308),
	.a(proc_output_control_planned_f),
	.b(n25408));
   no02m02 U28363 (.o(n25310),
	.a(n25309),
	.b(n25308));
   in01f01 U28364 (.o(n25318),
	.a(n26008));
   no02f02 U28365 (.o(n25324),
	.a(n25998),
	.b(n25984));
   in01s01 U28366 (.o(n25320),
	.a(n25319));
   na02s01 U28367 (.o(n25323),
	.a(FE_OFN25596_reset),
	.b(n25320));
   na02s01 U28368 (.o(n25334),
	.a(validIn_E),
	.b(east_input_NIB_elements_in_array_f_0_));
   in01s01 U28369 (.o(n25326),
	.a(n25334));
   no02s01 U28370 (.o(n25327),
	.a(east_input_NIB_elements_in_array_f_2_),
	.b(n25326));
   in01s01 U28371 (.o(n25331),
	.a(east_input_NIB_elements_in_array_f_2_));
   no02s01 U28372 (.o(n25340),
	.a(n25328),
	.b(n25331));
   in01s01 U28373 (.o(n25332),
	.a(east_input_NIB_elements_in_array_f_1_));
   oa22s01 U28374 (.o(n25333),
	.a(east_input_NIB_elements_in_array_f_2_),
	.b(n25332),
	.c(east_input_NIB_elements_in_array_f_1_),
	.d(n25331));
   in01f01 U28375 (.o(n25335),
	.a(n25998));
   ao22s01 U28376 (.o(n25344),
	.a(south_input_NIB_elements_in_array_f_1_),
	.b(n25343),
	.c(n18616),
	.d(n25345));
   in01s01 U28377 (.o(n25346),
	.a(n25347));
   ao22s01 U28378 (.o(n25348),
	.a(south_input_NIB_elements_in_array_f_1_),
	.b(n25347),
	.c(n25346),
	.d(n25345));
   in01s01 U28379 (.o(n25351),
	.a(north_output_space_yummy_f));
   in01s01 U28380 (.o(n25369),
	.a(north_output_space_count_f_0_));
   in01s01 U28381 (.o(n25358),
	.a(n25352));
   na02s01 U28382 (.o(n25367),
	.a(n25372),
	.b(north_output_space_count_f_2_));
   na02s01 U28383 (.o(n25357),
	.a(n25370),
	.b(n25367));
   in01s01 U28384 (.o(n25353),
	.a(north_output_space_count_f_1_));
   no02s01 U28385 (.o(n25354),
	.a(north_output_space_count_f_0_),
	.b(n25353));
   in01s01 U28386 (.o(n25356),
	.a(n25355));
   in01s01 U28387 (.o(n25371),
	.a(north_output_space_count_f_2_));
   in01s01 U28388 (.o(n25361),
	.a(n25374));
   na02s01 U28389 (.o(n25360),
	.a(north_output_space_count_f_0_),
	.b(north_output_space_count_f_1_));
   in01s01 U28390 (.o(n25362),
	.a(n25363));
   na02s01 U28391 (.o(n25366),
	.a(n25371),
	.b(n25362));
   na02s01 U28392 (.o(n25365),
	.a(north_output_space_count_f_2_),
	.b(n25363));
   na02s01 U28393 (.o(n25364),
	.a(n25370),
	.b(n25372));
   no02s01 U28394 (.o(n25376),
	.a(north_output_space_count_f_0_),
	.b(n25368));
   na02s01 U28395 (.o(n25373),
	.a(n25372),
	.b(n25371));
   ao22s01 U28396 (.o(n25378),
	.a(west_input_NIB_elements_in_array_f_1_),
	.b(n25377),
	.c(n18641),
	.d(n25379));
   in01s01 U28397 (.o(n25380),
	.a(n25381));
   na02s01 U28398 (.o(n25402),
	.a(east_output_current_route_connection_1_),
	.b(FE_OFN25598_reset));
   in01s01 U28399 (.o(n25410),
	.a(n25409));
   in01s01 U28401 (.o(n25439),
	.a(west_output_space_count_f_0_));
   no02s01 U28402 (.o(n25435),
	.a(n25459),
	.b(west_output_space_count_f_1_));
   in01s01 U28403 (.o(n25443),
	.a(n25435));
   na02s01 U28404 (.o(n25453),
	.a(n25457),
	.b(west_output_space_count_f_2_));
   in01s01 U28405 (.o(n25437),
	.a(n25453));
   no02s01 U28406 (.o(n25438),
	.a(n25437),
	.b(n25491));
   in01s01 U28407 (.o(n25442),
	.a(n25438));
   na02s01 U28408 (.o(n25440),
	.a(west_output_space_count_f_1_),
	.b(n25439));
   na02s01 U28409 (.o(n25441),
	.a(n25491),
	.b(n25440));
   in01s01 U28410 (.o(n25456),
	.a(west_output_space_count_f_2_));
   in01s01 U28411 (.o(n25446),
	.a(n25459));
   na02s01 U28412 (.o(n25445),
	.a(west_output_space_count_f_0_),
	.b(west_output_space_count_f_1_));
   in01s01 U28413 (.o(n25447),
	.a(n25448));
   na02s01 U28414 (.o(n25452),
	.a(n25456),
	.b(n25447));
   na02s01 U28415 (.o(n25451),
	.a(west_output_space_count_f_2_),
	.b(n25448));
   in01s01 U28416 (.o(n25449),
	.a(n25491));
   na02s01 U28417 (.o(n25450),
	.a(n25449),
	.b(n25457));
   na02s01 U28418 (.o(n25454),
	.a(n25459),
	.b(n25453));
   na02s01 U28419 (.o(n25455),
	.a(west_output_space_count_f_0_),
	.b(n25491));
   na02s01 U28420 (.o(n25458),
	.a(n25457),
	.b(n25456));
   no02s01 U28421 (.o(west_output_space_N47),
	.a(n25821),
	.b(west_output_space_N48));
   ao12f02 U28422 (.o(south_input_control_N51),
	.a(n26026),
	.b(FE_OFN575_n25463),
	.c(n25462));
   no02s01 U28423 (.o(n25468),
	.a(n25464),
	.b(n25482));
   in01f01 U28424 (.o(n25471),
	.a(proc_input_NIB_elements_in_array_f_2_));
   na03f01 U28425 (.o(n25466),
	.a(n25979),
	.b(proc_input_NIB_elements_in_array_f_3_),
	.c(n25471));
   na03f01 U28426 (.o(n25465),
	.a(n25974),
	.b(proc_input_NIB_elements_in_array_f_2_),
	.c(proc_input_NIB_elements_in_array_f_3_));
   no02s01 U28427 (.o(n25480),
	.a(n25468),
	.b(n25467));
   no02s01 U28428 (.o(n25473),
	.a(n25472),
	.b(n25471));
   in01f02 U28429 (.o(n25488),
	.a(n25485));
   na02f01 U28430 (.o(n25487),
	.a(proc_input_NIB_elements_in_array_f_3_),
	.b(n25486));
   in01s01 U28431 (.o(n25493),
	.a(west_output_space_is_two_or_more_f));
   ao22s01 U28432 (.o(n25501),
	.a(FE_OFN396_n19493),
	.b(n25516),
	.c(FE_OFN93_n21667),
	.d(n25518));
   na03f01 U28433 (.o(dataOut_S_59_),
	.a(n25502),
	.b(n25501),
	.c(n25500));
   ao22f01 U28434 (.o(n25504),
	.a(FE_OFN35_n19017),
	.b(n25512),
	.c(n19020),
	.d(FE_OFN579_n25511));
   na03m02 U28435 (.o(dataOut_E_51_),
	.a(n25505),
	.b(n25504),
	.c(n25503));
   ao22f01 U28436 (.o(n25508),
	.a(FE_OFN35_n19017),
	.b(n25497),
	.c(n19020),
	.d(n25518));
   na03m02 U28437 (.o(dataOut_E_59_),
	.a(n25509),
	.b(n25508),
	.c(n25507));
   ao22f01 U28438 (.o(n25514),
	.a(FE_OFN44_n19054),
	.b(n25512),
	.c(FE_OFN47_n19056),
	.d(FE_OFN579_n25511));
   ao22f01 U28440 (.o(n25523),
	.a(FE_OFN44_n19054),
	.b(n25497),
	.c(FE_OFN47_n19056),
	.d(n25518));
   na03f02 U28441 (.o(dataOut_N_59_),
	.a(n25524),
	.b(n25523),
	.c(n25522));
   in01s01 U28442 (.o(n3243),
	.a(n25525));
   in01s01 U28443 (.o(n3303),
	.a(n25526));
   in01s01 U28444 (.o(n3308),
	.a(n25527));
   in01s01 U28445 (.o(n3313),
	.a(n25528));
   in01s01 U28446 (.o(n3318),
	.a(n25529));
   in01s01 U28447 (.o(n3323),
	.a(n25530));
   in01s01 U28448 (.o(n3328),
	.a(n25531));
   in01s01 U28449 (.o(n3333),
	.a(n25532));
   in01s01 U28450 (.o(n3338),
	.a(n25533));
   in01s01 U28451 (.o(n3348),
	.a(n25535));
   in01s01 U28452 (.o(n3353),
	.a(n25536));
   in01s01 U28453 (.o(n3358),
	.a(n25537));
   in01s01 U28454 (.o(n3363),
	.a(n25538));
   in01s01 U28455 (.o(n3368),
	.a(n25539));
   in01s01 U28456 (.o(n3373),
	.a(n25540));
   in01s01 U28457 (.o(n3378),
	.a(n25541));
   in01s01 U28458 (.o(n3383),
	.a(n25542));
   in01s01 U28459 (.o(n3388),
	.a(n25543));
   in01s01 U28460 (.o(n3393),
	.a(n25544));
   in01s01 U28461 (.o(n3398),
	.a(n25545));
   in01s01 U28462 (.o(n3403),
	.a(n25546));
   in01s01 U28463 (.o(n3408),
	.a(n25548));
   oa22m01 U28464 (.o(n25549),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_1__33_),
	.d(n25571));
   in01s01 U28465 (.o(n3563),
	.a(n25549));
   oa22m01 U28466 (.o(n25550),
	.a(FE_OFN374_n17762),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_1__21_),
	.d(n25571));
   in01s01 U28467 (.o(n3623),
	.a(n25550));
   oa22m01 U28468 (.o(n25551),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_1__20_),
	.d(n25571));
   in01s01 U28469 (.o(n3628),
	.a(n25551));
   oa22m01 U28470 (.o(n25552),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_1__19_),
	.d(n25571));
   in01s01 U28471 (.o(n3633),
	.a(n25552));
   oa22m01 U28472 (.o(n25553),
	.a(FE_OFN374_n17762),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_1__18_),
	.d(n25571));
   in01s01 U28473 (.o(n3638),
	.a(n25553));
   oa22m01 U28474 (.o(n25554),
	.a(FE_OFN374_n17762),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_1__17_),
	.d(n25571));
   oa22m01 U28475 (.o(n25555),
	.a(FE_OFN374_n17762),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_1__16_),
	.d(n25571));
   in01s01 U28476 (.o(n3648),
	.a(n25555));
   oa22m01 U28477 (.o(n25556),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_1__15_),
	.d(n25571));
   in01s01 U28478 (.o(n3653),
	.a(n25556));
   oa22m01 U28479 (.o(n25557),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_1__14_),
	.d(n25571));
   in01s01 U28480 (.o(n3658),
	.a(n25557));
   oa22m01 U28481 (.o(n25558),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_1__13_),
	.d(n25571));
   in01s01 U28482 (.o(n3663),
	.a(n25558));
   oa22m01 U28483 (.o(n25559),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_1__12_),
	.d(n25571));
   in01s01 U28484 (.o(n3668),
	.a(n25559));
   oa22m01 U28485 (.o(n25560),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_1__11_),
	.d(n25571));
   in01s01 U28486 (.o(n3673),
	.a(n25560));
   oa22m01 U28487 (.o(n25561),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_1__10_),
	.d(n25571));
   in01s01 U28488 (.o(n3678),
	.a(n25561));
   in01s01 U28489 (.o(n3683),
	.a(n25562));
   oa22m01 U28490 (.o(n25563),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_1__8_),
	.d(n25571));
   in01s01 U28491 (.o(n3688),
	.a(n25563));
   oa22m01 U28492 (.o(n25564),
	.a(FE_OFN374_n17762),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_1__7_),
	.d(n25571));
   in01s01 U28493 (.o(n3693),
	.a(n25564));
   oa22m01 U28494 (.o(n25565),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_1__6_),
	.d(n25571));
   in01s01 U28495 (.o(n3698),
	.a(n25565));
   oa22m01 U28496 (.o(n25566),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_1__5_),
	.d(n25571));
   in01s01 U28497 (.o(n3703),
	.a(n25566));
   oa22m01 U28498 (.o(n25567),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_1__4_),
	.d(n25571));
   in01s01 U28499 (.o(n3708),
	.a(n25567));
   oa22m01 U28500 (.o(n25568),
	.a(FE_OFN374_n17762),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_1__3_),
	.d(n25571));
   in01s01 U28501 (.o(n3713),
	.a(n25568));
   oa22m01 U28502 (.o(n25569),
	.a(FE_OFN373_n17762),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_1__2_),
	.d(n25571));
   oa22m01 U28503 (.o(n25570),
	.a(FE_OFN374_n17762),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_1__1_),
	.d(n25571));
   in01s01 U28504 (.o(n3723),
	.a(n25570));
   in01s01 U28505 (.o(n3728),
	.a(n25572));
   oa22m01 U28506 (.o(n25573),
	.a(n17764),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_2__33_),
	.d(n25595));
   in01s01 U28507 (.o(n3883),
	.a(n25573));
   oa22m01 U28508 (.o(n25574),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_2__21_),
	.d(n25595));
   oa22m01 U28509 (.o(n25575),
	.a(n17764),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_2__20_),
	.d(n25595));
   in01s01 U28510 (.o(n3948),
	.a(n25575));
   oa22m01 U28511 (.o(n25576),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_2__19_),
	.d(n25595));
   in01s01 U28512 (.o(n3953),
	.a(n25576));
   oa22m01 U28513 (.o(n25577),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_2__18_),
	.d(n25595));
   in01s01 U28514 (.o(n3958),
	.a(n25577));
   oa22m01 U28515 (.o(n25578),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_2__17_),
	.d(n25595));
   in01s01 U28516 (.o(n3963),
	.a(n25578));
   oa22m01 U28517 (.o(n25579),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_2__16_),
	.d(n25595));
   in01s01 U28518 (.o(n3968),
	.a(n25579));
   in01s01 U28519 (.o(n3973),
	.a(n25580));
   oa22m01 U28520 (.o(n25581),
	.a(n17764),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_2__14_),
	.d(n25595));
   in01s01 U28521 (.o(n3978),
	.a(n25581));
   oa22m01 U28522 (.o(n25582),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_2__13_),
	.d(n25595));
   in01s01 U28523 (.o(n3983),
	.a(n25582));
   oa22m01 U28524 (.o(n25583),
	.a(n17764),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_2__12_),
	.d(n25595));
   in01s01 U28525 (.o(n3988),
	.a(n25583));
   oa22m01 U28526 (.o(n25584),
	.a(FE_OFN272_n25595),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_2__11_),
	.d(n25595));
   in01s01 U28527 (.o(n3993),
	.a(n25584));
   in01s01 U28528 (.o(n3998),
	.a(n25585));
   in01s01 U28529 (.o(n4003),
	.a(n25586));
   in01s01 U28530 (.o(n4008),
	.a(n25587));
   in01s01 U28531 (.o(n4013),
	.a(n25588));
   in01s01 U28532 (.o(n4023),
	.a(n25590));
   in01s01 U28533 (.o(n4028),
	.a(n25591));
   in01s01 U28534 (.o(n4033),
	.a(n25592));
   in01s01 U28535 (.o(n4038),
	.a(n25593));
   in01s01 U28536 (.o(n4043),
	.a(n25594));
   in01s01 U28537 (.o(n4048),
	.a(n25596));
   oa22m01 U28538 (.o(n25597),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_3__33_),
	.d(n25619));
   in01s01 U28539 (.o(n4203),
	.a(n25597));
   in01s01 U28540 (.o(n4263),
	.a(n25598));
   oa22m01 U28541 (.o(n25599),
	.a(FE_OFN25777_FE_OFN582_n25619),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_3__20_),
	.d(n17763));
   in01s01 U28542 (.o(n4268),
	.a(n25599));
   oa22m01 U28543 (.o(n25600),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_19_),
	.c(proc_input_NIB_storage_data_f_3__19_),
	.d(n25619));
   in01s01 U28544 (.o(n4273),
	.a(n25600));
   oa22m01 U28545 (.o(n25601),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_18_),
	.c(proc_input_NIB_storage_data_f_3__18_),
	.d(n25619));
   in01s01 U28546 (.o(n4278),
	.a(n25601));
   oa22m01 U28547 (.o(n25602),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_17_),
	.c(proc_input_NIB_storage_data_f_3__17_),
	.d(n25619));
   in01s01 U28548 (.o(n4283),
	.a(n25602));
   oa22m01 U28549 (.o(n25603),
	.a(FE_OFN25777_FE_OFN582_n25619),
	.b(dataIn_P_16_),
	.c(proc_input_NIB_storage_data_f_3__16_),
	.d(n17763));
   in01s01 U28550 (.o(n4288),
	.a(n25603));
   oa22m01 U28551 (.o(n25604),
	.a(FE_OFN582_n25619),
	.b(dataIn_P_15_),
	.c(proc_input_NIB_storage_data_f_3__15_),
	.d(n25619));
   in01s01 U28552 (.o(n4293),
	.a(n25604));
   oa22m01 U28553 (.o(n25605),
	.a(FE_OFN25777_FE_OFN582_n25619),
	.b(dataIn_P_14_),
	.c(proc_input_NIB_storage_data_f_3__14_),
	.d(n17763));
   in01s01 U28554 (.o(n4298),
	.a(n25605));
   oa22m01 U28555 (.o(n25606),
	.a(FE_OFN25776_FE_OFN582_n25619),
	.b(dataIn_P_13_),
	.c(proc_input_NIB_storage_data_f_3__13_),
	.d(n25619));
   in01s01 U28556 (.o(n4303),
	.a(n25606));
   oa22m01 U28557 (.o(n25607),
	.a(FE_OFN25777_FE_OFN582_n25619),
	.b(dataIn_P_12_),
	.c(proc_input_NIB_storage_data_f_3__12_),
	.d(n17763));
   in01s01 U28558 (.o(n4308),
	.a(n25607));
   oa22m01 U28559 (.o(n25608),
	.a(FE_OFN25777_FE_OFN582_n25619),
	.b(dataIn_P_11_),
	.c(proc_input_NIB_storage_data_f_3__11_),
	.d(n17763));
   in01s01 U28560 (.o(n4313),
	.a(n25608));
   in01s01 U28561 (.o(n4323),
	.a(n25610));
   in01s01 U28562 (.o(n4328),
	.a(n25611));
   in01s01 U28563 (.o(n4333),
	.a(n25612));
   in01s01 U28564 (.o(n4338),
	.a(n25613));
   in01s01 U28566 (.o(n4348),
	.a(n25615));
   in01s01 U28567 (.o(n4353),
	.a(n25616));
   in01s01 U28568 (.o(n4358),
	.a(n25617));
   in01s01 U28569 (.o(n4363),
	.a(n25618));
   in01s01 U28570 (.o(n4368),
	.a(n25620));
   oa22s01 U28571 (.o(n25621),
	.a(n22273),
	.b(dataIn_P_33_),
	.c(proc_input_NIB_storage_data_f_15__33_),
	.d(n25643));
   in01s01 U28572 (.o(n8043),
	.a(n25621));
   oa22s01 U28573 (.o(n25622),
	.a(FE_OFN584_n25643),
	.b(dataIn_P_21_),
	.c(proc_input_NIB_storage_data_f_15__21_),
	.d(n25643));
   in01s01 U28574 (.o(n8103),
	.a(n25622));
   oa22s01 U28575 (.o(n25623),
	.a(n22273),
	.b(dataIn_P_20_),
	.c(proc_input_NIB_storage_data_f_15__20_),
	.d(n25643));
   in01s01 U28576 (.o(n8108),
	.a(n25623));
   in01s01 U28577 (.o(n8113),
	.a(n25624));
   in01s01 U28578 (.o(n8118),
	.a(n25625));
   in01s01 U28579 (.o(n8123),
	.a(n25626));
   in01s01 U28580 (.o(n8128),
	.a(n25627));
   in01s01 U28581 (.o(n8133),
	.a(n25628));
   in01s01 U28582 (.o(n8138),
	.a(n25629));
   in01s01 U28583 (.o(n8148),
	.a(n25631));
   in01s01 U28584 (.o(n8153),
	.a(n25632));
   oa22s01 U28585 (.o(n25633),
	.a(FE_OFN584_n25643),
	.b(dataIn_P_10_),
	.c(proc_input_NIB_storage_data_f_15__10_),
	.d(n25643));
   in01s01 U28586 (.o(n8158),
	.a(n25633));
   oa22s01 U28587 (.o(n25634),
	.a(FE_OFN584_n25643),
	.b(dataIn_P_9_),
	.c(proc_input_NIB_storage_data_f_15__9_),
	.d(n25643));
   in01s01 U28588 (.o(n8163),
	.a(n25634));
   oa22s01 U28589 (.o(n25635),
	.a(FE_OFN584_n25643),
	.b(dataIn_P_8_),
	.c(proc_input_NIB_storage_data_f_15__8_),
	.d(n25643));
   in01s01 U28590 (.o(n8168),
	.a(n25635));
   oa22s01 U28591 (.o(n25636),
	.a(FE_OFN584_n25643),
	.b(dataIn_P_7_),
	.c(proc_input_NIB_storage_data_f_15__7_),
	.d(n25643));
   in01s01 U28592 (.o(n8173),
	.a(n25636));
   oa22s01 U28593 (.o(n25637),
	.a(FE_OFN584_n25643),
	.b(dataIn_P_6_),
	.c(proc_input_NIB_storage_data_f_15__6_),
	.d(n25643));
   in01s01 U28594 (.o(n8178),
	.a(n25637));
   oa22s01 U28595 (.o(n25638),
	.a(FE_OFN584_n25643),
	.b(dataIn_P_5_),
	.c(proc_input_NIB_storage_data_f_15__5_),
	.d(n25643));
   in01s01 U28596 (.o(n8183),
	.a(n25638));
   oa22s01 U28597 (.o(n25639),
	.a(n22273),
	.b(dataIn_P_4_),
	.c(proc_input_NIB_storage_data_f_15__4_),
	.d(n25643));
   in01s01 U28598 (.o(n8188),
	.a(n25639));
   oa22s01 U28599 (.o(n25640),
	.a(FE_OFN584_n25643),
	.b(dataIn_P_3_),
	.c(proc_input_NIB_storage_data_f_15__3_),
	.d(n25643));
   in01s01 U28600 (.o(n8193),
	.a(n25640));
   oa22s01 U28601 (.o(n25641),
	.a(FE_OFN584_n25643),
	.b(dataIn_P_2_),
	.c(proc_input_NIB_storage_data_f_15__2_),
	.d(n25643));
   in01s01 U28602 (.o(n8198),
	.a(n25641));
   oa22s01 U28603 (.o(n25642),
	.a(FE_OFN584_n25643),
	.b(dataIn_P_1_),
	.c(proc_input_NIB_storage_data_f_15__1_),
	.d(n25643));
   in01s01 U28604 (.o(n8203),
	.a(n25642));
   oa22s01 U28605 (.o(n25644),
	.a(FE_OFN584_n25643),
	.b(dataIn_P_0_),
	.c(proc_input_NIB_storage_data_f_15__0_),
	.d(n25643));
   in01s01 U28606 (.o(n8208),
	.a(n25644));
   oa22f01 U28607 (.o(n25645),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_33_),
	.c(east_input_NIB_storage_data_f_0__33_),
	.d(FE_OFN24862_n22945));
   in01s01 U28608 (.o(n10963),
	.a(n25645));
   oa22f01 U28609 (.o(n25646),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_21_),
	.c(east_input_NIB_storage_data_f_0__21_),
	.d(FE_OFN24862_n22945));
   in01s01 U28610 (.o(n11023),
	.a(n25646));
   oa22f01 U28611 (.o(n25647),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_20_),
	.c(east_input_NIB_storage_data_f_0__20_),
	.d(FE_OFN24862_n22945));
   in01s01 U28612 (.o(n11028),
	.a(n25647));
   oa22f01 U28613 (.o(n25648),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_19_),
	.c(east_input_NIB_storage_data_f_0__19_),
	.d(FE_OFN24862_n22945));
   in01s01 U28614 (.o(n11033),
	.a(n25648));
   oa22f01 U28615 (.o(n25649),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_18_),
	.c(east_input_NIB_storage_data_f_0__18_),
	.d(FE_OFN24862_n22945));
   in01s01 U28616 (.o(n11038),
	.a(n25649));
   oa22f01 U28617 (.o(n25650),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_17_),
	.c(east_input_NIB_storage_data_f_0__17_),
	.d(FE_OFN24862_n22945));
   in01s01 U28618 (.o(n11043),
	.a(n25650));
   oa22f01 U28619 (.o(n25651),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_15_),
	.c(east_input_NIB_storage_data_f_0__15_),
	.d(FE_OFN24862_n22945));
   in01s01 U28620 (.o(n11053),
	.a(n25651));
   oa22f01 U28621 (.o(n25652),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_13_),
	.c(east_input_NIB_storage_data_f_0__13_),
	.d(FE_OFN24862_n22945));
   in01s01 U28622 (.o(n11063),
	.a(n25652));
   oa22f01 U28623 (.o(n25653),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_12_),
	.c(east_input_NIB_storage_data_f_0__12_),
	.d(FE_OFN24862_n22945));
   oa22f01 U28624 (.o(n25654),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_11_),
	.c(east_input_NIB_storage_data_f_0__11_),
	.d(FE_OFN24862_n22945));
   in01s01 U28625 (.o(n11073),
	.a(n25654));
   oa22f01 U28626 (.o(n25655),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_10_),
	.c(east_input_NIB_storage_data_f_0__10_),
	.d(FE_OFN24862_n22945));
   in01s01 U28627 (.o(n11078),
	.a(n25655));
   oa22f01 U28628 (.o(n25656),
	.a(FE_OFN24861_n22945),
	.b(dataIn_E_9_),
	.c(east_input_NIB_storage_data_f_0__9_),
	.d(FE_OFN24862_n22945));
   in01s01 U28629 (.o(n11083),
	.a(n25656));
   in01s01 U28630 (.o(n11088),
	.a(n25657));
   in01s01 U28631 (.o(n11093),
	.a(n25658));
   in01s01 U28632 (.o(n11098),
	.a(n25659));
   in01s01 U28633 (.o(n11108),
	.a(n25660));
   in01s01 U28634 (.o(n11123),
	.a(n25661));
   in01s01 U28635 (.o(n11283),
	.a(n25662));
   in01s01 U28636 (.o(n11343),
	.a(n25663));
   in01s01 U28637 (.o(n11348),
	.a(n25664));
   in01s01 U28638 (.o(n11353),
	.a(n25665));
   in01s01 U28639 (.o(n11358),
	.a(n25666));
   in01s01 U28640 (.o(n11363),
	.a(n25667));
   in01s01 U28641 (.o(n11373),
	.a(n25668));
   in01s01 U28642 (.o(n11383),
	.a(n25669));
   in01s01 U28643 (.o(n11388),
	.a(n25670));
   in01s01 U28644 (.o(n11393),
	.a(n25671));
   in01s01 U28645 (.o(n11398),
	.a(n25672));
   in01s01 U28646 (.o(n11403),
	.a(n25673));
   in01s01 U28647 (.o(n11408),
	.a(n25674));
   in01s01 U28648 (.o(n11413),
	.a(n25675));
   in01s01 U28649 (.o(n11418),
	.a(n25676));
   in01s01 U28650 (.o(n11428),
	.a(n25677));
   oa22f01 U28651 (.o(n25679),
	.a(FE_OFN24808_n22958),
	.b(dataIn_E_33_),
	.c(east_input_NIB_storage_data_f_2__33_),
	.d(FE_OFN435_n22958));
   in01s01 U28652 (.o(n11603),
	.a(n25679));
   oa22f01 U28653 (.o(n25680),
	.a(FE_OFN24815_n22958),
	.b(dataIn_E_21_),
	.c(east_input_NIB_storage_data_f_2__21_),
	.d(FE_OFN435_n22958));
   in01s01 U28654 (.o(n11663),
	.a(n25680));
   oa22f01 U28655 (.o(n25681),
	.a(FE_OFN24807_n22958),
	.b(dataIn_E_20_),
	.c(east_input_NIB_storage_data_f_2__20_),
	.d(FE_OFN435_n22958));
   oa22f01 U28656 (.o(n25682),
	.a(FE_OFN24815_n22958),
	.b(dataIn_E_19_),
	.c(east_input_NIB_storage_data_f_2__19_),
	.d(FE_OFN435_n22958));
   in01s01 U28657 (.o(n11673),
	.a(n25682));
   oa22f01 U28658 (.o(n25683),
	.a(FE_OFN24812_n22958),
	.b(dataIn_E_18_),
	.c(east_input_NIB_storage_data_f_2__18_),
	.d(FE_OFN435_n22958));
   in01s01 U28659 (.o(n11678),
	.a(n25683));
   oa22f01 U28660 (.o(n25684),
	.a(FE_OFN24809_n22958),
	.b(dataIn_E_17_),
	.c(east_input_NIB_storage_data_f_2__17_),
	.d(FE_OFN435_n22958));
   in01s01 U28661 (.o(n11683),
	.a(n25684));
   oa22f01 U28662 (.o(n25685),
	.a(n22959),
	.b(dataIn_E_15_),
	.c(east_input_NIB_storage_data_f_2__15_),
	.d(FE_OFN435_n22958));
   in01s01 U28663 (.o(n11693),
	.a(n25685));
   oa22f01 U28664 (.o(n25686),
	.a(FE_OFN24810_n22958),
	.b(dataIn_E_13_),
	.c(east_input_NIB_storage_data_f_2__13_),
	.d(FE_OFN435_n22958));
   in01s01 U28665 (.o(n11703),
	.a(n25686));
   oa22f01 U28666 (.o(n25687),
	.a(FE_OFN438_n22958),
	.b(dataIn_E_12_),
	.c(east_input_NIB_storage_data_f_2__12_),
	.d(FE_OFN435_n22958));
   in01s01 U28667 (.o(n11708),
	.a(n25687));
   in01s01 U28668 (.o(n11713),
	.a(n25688));
   in01s01 U28669 (.o(n11718),
	.a(n25689));
   oa22f01 U28670 (.o(n25690),
	.a(FE_OFN24815_n22958),
	.b(dataIn_E_9_),
	.c(east_input_NIB_storage_data_f_2__9_),
	.d(FE_OFN435_n22958));
   in01s01 U28671 (.o(n11723),
	.a(n25690));
   oa22f01 U28672 (.o(n25691),
	.a(FE_OFN24814_n22958),
	.b(dataIn_E_8_),
	.c(east_input_NIB_storage_data_f_2__8_),
	.d(FE_OFN435_n22958));
   in01s01 U28673 (.o(n11728),
	.a(n25691));
   oa22f01 U28674 (.o(n25692),
	.a(FE_OFN24815_n22958),
	.b(dataIn_E_7_),
	.c(east_input_NIB_storage_data_f_2__7_),
	.d(FE_OFN435_n22958));
   in01s01 U28675 (.o(n11733),
	.a(n25692));
   in01s01 U28676 (.o(n11738),
	.a(n25693));
   in01s01 U28677 (.o(n11748),
	.a(n25694));
   in01s01 U28678 (.o(n11763),
	.a(n25695));
   in01s01 U28679 (.o(n11923),
	.a(n25696));
   in01s01 U28680 (.o(n11983),
	.a(n25697));
   in01s01 U28681 (.o(n11988),
	.a(n25698));
   in01s01 U28682 (.o(n11993),
	.a(n25699));
   in01s01 U28683 (.o(n11998),
	.a(n25700));
   in01s01 U28684 (.o(n12003),
	.a(n25701));
   in01s01 U28685 (.o(n12013),
	.a(n25702));
   in01s01 U28686 (.o(n12023),
	.a(n25703));
   in01s01 U28687 (.o(n12028),
	.a(n25704));
   in01s01 U28688 (.o(n12033),
	.a(n25705));
   in01s01 U28689 (.o(n12038),
	.a(n25706));
   in01s01 U28690 (.o(n12048),
	.a(n25708));
   in01s01 U28691 (.o(n12053),
	.a(n25709));
   in01s01 U28692 (.o(n12058),
	.a(n25710));
   in01s01 U28693 (.o(n12068),
	.a(n25711));
   in01s01 U28694 (.o(n12083),
	.a(n25712));
   in01s01 U28695 (.o(n25722),
	.a(ec_cfg_0_));
   ao22s01 U28696 (.o(n25716),
	.a(n25722),
	.b(ec_wants_to_send_but_cannot_P),
	.c(ec_cfg_0_),
	.d(ec_thanks_p_to_p_reg));
   in01s01 U28697 (.o(n25718),
	.a(ec_cfg_1_));
   no02s01 U28698 (.o(n25713),
	.a(n25718),
	.b(n25722));
   in01s01 U28699 (.o(n25715),
	.a(n25713));
   oa22s01 U28700 (.o(n25717),
	.a(ec_cfg_1_),
	.b(n25716),
	.c(n25715),
	.d(n25714));
   in01s01 U28701 (.o(n25734),
	.a(n25717));
   no02s01 U28702 (.o(n25732),
	.a(ec_cfg_0_),
	.b(n25718));
   ao22s01 U28703 (.o(n25719),
	.a(ec_thanks_e_to_p_reg),
	.b(n25722),
	.c(ec_thanks_n_to_p_reg),
	.d(ec_cfg_0_));
   no02s01 U28704 (.o(n25728),
	.a(ec_cfg_1_),
	.b(n25719));
   na02s01 U28705 (.o(n25724),
	.a(n25723),
	.b(ec_proc_input_valid_reg));
   in01s01 U28706 (.o(n25745),
	.a(ec_cfg_3_));
   in01s01 U28707 (.o(n25735),
	.a(ec_west_input_valid_reg));
   no02s01 U28708 (.o(n25740),
	.a(n25745),
	.b(n25735));
   no02s01 U28709 (.o(n25737),
	.a(ec_thanks_n_to_w_reg),
	.b(ec_thanks_p_to_w_reg));
   no03s01 U28710 (.o(n25736),
	.a(ec_thanks_e_to_w_reg),
	.b(ec_thanks_s_to_w_reg),
	.c(ec_thanks_w_to_w_reg));
   na02s01 U28711 (.o(n25739),
	.a(n25737),
	.b(n25736));
   na02s01 U28712 (.o(n25738),
	.a(ec_cfg_3_),
	.b(n25739));
   oa12s01 U28713 (.o(n25742),
	.a(n25738),
	.b(n25740),
	.c(n25739));
   ao22s01 U28714 (.o(n25741),
	.a(ec_thanks_n_to_w_reg),
	.b(ec_cfg_3_),
	.c(ec_thanks_e_to_w_reg),
	.d(n25745));
   in01s01 U28715 (.o(n25746),
	.a(ec_cfg_4_));
   na02s01 U28716 (.o(n25744),
	.a(ec_thanks_w_to_w_reg),
	.b(ec_cfg_4_));
   ao12s01 U28717 (.o(n25743),
	.a(n25746),
	.b(ec_cfg_3_),
	.c(ec_thanks_s_to_w_reg));
   oa22s01 U28718 (.o(n25749),
	.a(ec_cfg_3_),
	.b(n25744),
	.c(ec_cfg_5_),
	.d(n25743));
   ao22s01 U28719 (.o(n25747),
	.a(ec_thanks_p_to_w_reg),
	.b(ec_cfg_3_),
	.c(n25745),
	.d(ec_wants_to_send_but_cannot_W));
   na02s01 U28720 (.o(n25748),
	.a(n25747),
	.b(n25746));
   in01s01 U28721 (.o(ec_out_1_),
	.a(n25751));
   in01s01 U28722 (.o(n25758),
	.a(ec_cfg_7_));
   na02s01 U28723 (.o(n25764),
	.a(ec_cfg_6_),
	.b(n25758));
   in01s01 U28724 (.o(n25752),
	.a(ec_thanks_s_to_s_reg));
   no02s01 U28725 (.o(n25755),
	.a(n25757),
	.b(n25752));
   no02s01 U28726 (.o(n25754),
	.a(ec_cfg_7_),
	.b(n25753));
   oa22s01 U28727 (.o(n25772),
	.a(ec_thanks_p_to_s_reg),
	.b(n25764),
	.c(n25755),
	.d(n25754));
   no02s01 U28728 (.o(n25770),
	.a(ec_cfg_6_),
	.b(n25758));
   in01s01 U28729 (.o(n25757),
	.a(ec_cfg_6_));
   no04s01 U28730 (.o(n25761),
	.a(ec_thanks_w_to_s_reg),
	.b(n25758),
	.c(n25757),
	.d(n25756));
   no02s01 U28731 (.o(n25760),
	.a(ec_thanks_e_to_s_reg),
	.b(ec_thanks_n_to_s_reg));
   no02s01 U28732 (.o(n25759),
	.a(ec_thanks_s_to_s_reg),
	.b(ec_thanks_p_to_s_reg));
   na02s01 U28733 (.o(n25762),
	.a(n25760),
	.b(n25759));
   no02s01 U28734 (.o(n25768),
	.a(n25761),
	.b(n25762));
   in01s01 U28735 (.o(n25763),
	.a(n25762));
   no02s01 U28736 (.o(n25767),
	.a(n25770),
	.b(n25763));
   in01s01 U28737 (.o(n25777),
	.a(ec_cfg_10_));
   in01s01 U28738 (.o(n25773),
	.a(ec_thanks_s_to_e_reg));
   no02s01 U28739 (.o(n25776),
	.a(n25777),
	.b(n25773));
   in01s01 U28740 (.o(n25778),
	.a(ec_cfg_9_));
   ao22s01 U28741 (.o(n25774),
	.a(n25778),
	.b(ec_wants_to_send_but_cannot_E),
	.c(ec_cfg_9_),
	.d(ec_thanks_p_to_e_reg));
   no02s01 U28742 (.o(n25775),
	.a(n25774),
	.b(ec_cfg_10_));
   oa22s01 U28743 (.o(n25795),
	.a(n25776),
	.b(n25775),
	.c(n25777),
	.d(ec_cfg_9_));
   no02s01 U28744 (.o(n25793),
	.a(ec_cfg_9_),
	.b(n25777));
   ao22s01 U28745 (.o(n25779),
	.a(ec_thanks_e_to_e_reg),
	.b(n25778),
	.c(ec_thanks_n_to_e_reg),
	.d(ec_cfg_9_));
   no02s01 U28746 (.o(n25789),
	.a(ec_cfg_10_),
	.b(n25779));
   no02s01 U28747 (.o(n25781),
	.a(ec_thanks_e_to_e_reg),
	.b(ec_thanks_p_to_e_reg));
   no03f01 U28748 (.o(n25780),
	.a(ec_thanks_n_to_e_reg),
	.b(ec_thanks_w_to_e_reg),
	.c(ec_thanks_s_to_e_reg));
   na02f02 U28749 (.o(n25785),
	.a(n25781),
	.b(n25780));
   na02s01 U28750 (.o(n25782),
	.a(ec_cfg_9_),
	.b(ec_east_input_valid_reg));
   in01s01 U28751 (.o(n25783),
	.a(n25782));
   ao12s01 U28752 (.o(n25786),
	.a(n25784),
	.b(n25785),
	.c(ec_cfg_9_));
   na02s01 U28753 (.o(n25787),
	.a(ec_cfg_10_),
	.b(n25786));
   in01s01 U28754 (.o(n25788),
	.a(n25787));
   in01s01 U28755 (.o(n25790),
	.a(ec_cfg_11_));
   in01s01 U28756 (.o(n25804),
	.a(ec_cfg_12_));
   in01s01 U28757 (.o(n25796),
	.a(ec_north_input_valid_reg));
   no02s01 U28758 (.o(n25801),
	.a(n25804),
	.b(n25796));
   no02s01 U28759 (.o(n25798),
	.a(ec_thanks_s_to_n_reg),
	.b(ec_thanks_e_to_n_reg));
   no03s01 U28760 (.o(n25797),
	.a(ec_thanks_p_to_n_reg),
	.b(ec_thanks_w_to_n_reg),
	.c(ec_thanks_n_to_n_reg));
   na02s01 U28761 (.o(n25800),
	.a(n25798),
	.b(n25797));
   na02s01 U28762 (.o(n25799),
	.a(ec_cfg_12_),
	.b(n25800));
   oa12s01 U28763 (.o(n25803),
	.a(n25799),
	.b(n25801),
	.c(n25800));
   ao22s01 U28764 (.o(n25802),
	.a(ec_cfg_12_),
	.b(ec_thanks_n_to_n_reg),
	.c(n25804),
	.d(ec_thanks_e_to_n_reg));
   in01s01 U28765 (.o(n25808),
	.a(ec_cfg_13_));
   ao22s01 U28766 (.o(n25807),
	.a(ec_thanks_p_to_n_reg),
	.b(ec_cfg_12_),
	.c(n25804),
	.d(ec_wants_to_send_but_cannot_N));
   in01s01 U28767 (.o(n25805),
	.a(ec_thanks_w_to_n_reg));
   ao22s01 U28768 (.o(n25811),
	.a(n25808),
	.b(n25807),
	.c(n25806),
	.d(n25805));
   no02s01 U28769 (.o(n25809),
	.a(n25808),
	.b(ec_thanks_s_to_n_reg));
   oa22s01 U28770 (.o(n25810),
	.a(ec_cfg_14_),
	.b(n25809),
	.c(ec_cfg_12_),
	.d(n25808));
   in01s01 U28771 (.o(ec_out_4_),
	.a(n25813));
   no02f01 U28772 (.o(north_output_space_N42),
	.a(FE_OFN25601_reset),
	.b(n25814));
   no02f01 U28773 (.o(north_output_space_N43),
	.a(FE_OFN25601_reset),
	.b(n25815));
   na02s01 U28774 (.o(north_output_space_N44),
	.a(FE_OFN25596_reset),
	.b(n25816));
   no02f01 U28775 (.o(east_output_space_N42),
	.a(FE_OFN25601_reset),
	.b(n25817));
   no02f01 U28776 (.o(east_output_space_N43),
	.a(FE_OFN25601_reset),
	.b(n25818));
   no02f01 U28777 (.o(south_output_space_N42),
	.a(reset),
	.b(n25819));
   no02f01 U28778 (.o(south_output_space_N43),
	.a(reset),
	.b(n25820));
   no02f01 U28779 (.o(west_output_space_N42),
	.a(FE_OFN25601_reset),
	.b(n25821));
   no02f01 U28780 (.o(west_output_space_N43),
	.a(FE_OFN25601_reset),
	.b(n25822));
   na02s01 U28781 (.o(west_output_space_N44),
	.a(FE_OFN25596_reset),
	.b(n25823));
   no02f01 U28782 (.o(proc_output_space_N42),
	.a(reset),
	.b(n25824));
   no02f01 U28783 (.o(proc_output_space_N43),
	.a(reset),
	.b(n25825));
   na02s01 U28785 (.o(n25828),
	.a(FE_OFN575_n25463),
	.b(n25830));
   in01s01 U28786 (.o(n25827),
	.a(n25826));
   oa12s01 U28787 (.o(n13388),
	.a(n25827),
	.b(n25829),
	.c(n25828));
   na03s01 U28788 (.o(n25831),
	.a(north_input_NIB_tail_ptr_f_1_),
	.b(FE_OFN575_n25463),
	.c(n25830));
   in01s01 U28789 (.o(n25832),
	.a(north_input_NIB_storage_data_f_3__6_));
   in01s01 U28790 (.o(n25853),
	.a(dataIn_N_13_));
   in01s01 U28791 (.o(n25833),
	.a(north_input_NIB_storage_data_f_3__13_));
   ao22f01 U28792 (.o(n13313),
	.a(n21175),
	.b(n25853),
	.c(n25833),
	.d(FE_OFN86_n21175));
   in01s01 U28793 (.o(n25834),
	.a(north_input_NIB_storage_data_f_3__18_));
   ao22f01 U28794 (.o(n13288),
	.a(n21175),
	.b(n25855),
	.c(n25834),
	.d(FE_OFN86_n21175));
   in01s01 U28795 (.o(n25857),
	.a(dataIn_N_19_));
   in01s01 U28796 (.o(n25835),
	.a(north_input_NIB_storage_data_f_3__19_));
   ao22f01 U28797 (.o(n13283),
	.a(n21175),
	.b(n25857),
	.c(n25835),
	.d(FE_OFN86_n21175));
   in01s01 U28798 (.o(n25859),
	.a(dataIn_N_21_));
   in01s01 U28799 (.o(n25837),
	.a(north_input_NIB_storage_data_f_3__21_));
   ao22f01 U28800 (.o(n13273),
	.a(n21175),
	.b(n25859),
	.c(n25837),
	.d(FE_OFN86_n21175));
   in01s01 U28801 (.o(n25838),
	.a(north_input_NIB_storage_data_f_2__6_));
   in01s01 U28802 (.o(n25839),
	.a(north_input_NIB_storage_data_f_2__13_));
   ao22f01 U28803 (.o(n12993),
	.a(n20656),
	.b(n25853),
	.c(n25839),
	.d(FE_OFN25876_n25842));
   in01s01 U28804 (.o(n25840),
	.a(north_input_NIB_storage_data_f_2__18_));
   ao22f01 U28805 (.o(n12968),
	.a(n20656),
	.b(n25855),
	.c(n25840),
	.d(FE_OFN25876_n25842));
   in01s01 U28806 (.o(n25841),
	.a(north_input_NIB_storage_data_f_2__19_));
   ao22f01 U28807 (.o(n12963),
	.a(n20656),
	.b(n25857),
	.c(n25841),
	.d(FE_OFN25876_n25842));
   in01s01 U28808 (.o(n25843),
	.a(north_input_NIB_storage_data_f_2__21_));
   ao22f01 U28809 (.o(n12953),
	.a(n20656),
	.b(n25859),
	.c(n25843),
	.d(FE_OFN25876_n25842));
   in01s01 U28810 (.o(n25844),
	.a(north_input_NIB_storage_data_f_1__6_));
   ao22f01 U28811 (.o(n12708),
	.a(n21220),
	.b(n25851),
	.c(n25844),
	.d(n25848));
   in01s01 U28812 (.o(n25845),
	.a(north_input_NIB_storage_data_f_1__13_));
   ao22f01 U28813 (.o(n12673),
	.a(n21220),
	.b(n25853),
	.c(n25845),
	.d(n25848));
   in01s01 U28814 (.o(n25846),
	.a(north_input_NIB_storage_data_f_1__18_));
   ao22f01 U28815 (.o(n12648),
	.a(n21220),
	.b(n25855),
	.c(n25846),
	.d(n25848));
   in01s01 U28816 (.o(n25847),
	.a(north_input_NIB_storage_data_f_1__19_));
   in01s01 U28817 (.o(n25849),
	.a(north_input_NIB_storage_data_f_1__21_));
   ao22f01 U28818 (.o(n12633),
	.a(n21220),
	.b(n25859),
	.c(n25849),
	.d(n25848));
   in01s01 U28819 (.o(n25850),
	.a(north_input_NIB_storage_data_f_0__6_));
   in01s01 U28820 (.o(n25852),
	.a(north_input_NIB_storage_data_f_0__13_));
   in01s01 U28821 (.o(n25854),
	.a(north_input_NIB_storage_data_f_0__18_));
   in01s01 U28822 (.o(n25856),
	.a(north_input_NIB_storage_data_f_0__19_));
   in01s01 U28823 (.o(n25858),
	.a(north_input_NIB_storage_data_f_0__21_));
   oa12s01 U28824 (.o(n25860),
	.a(FE_OFN25596_reset),
	.b(validIn_E),
	.c(east_input_NIB_tail_ptr_f_0_));
   ao12s01 U28825 (.o(n12098),
	.a(n25860),
	.b(validIn_E),
	.c(east_input_NIB_tail_ptr_f_0_));
   na02s01 U28826 (.o(n25861),
	.a(east_input_NIB_tail_ptr_f_1_),
	.b(FE_OFN25596_reset));
   oa12s01 U28827 (.o(n12093),
	.a(FE_OFN951_n25881),
	.b(n25862),
	.c(n25861));
   in01s01 U28828 (.o(n25884),
	.a(dataIn_E_0_));
   in01s01 U28829 (.o(n25863),
	.a(east_input_NIB_storage_data_f_3__0_));
   ao22s01 U28830 (.o(n12088),
	.a(FE_OFN940_n24921),
	.b(n25884),
	.c(n25863),
	.d(FE_OFN24823_n24921));
   in01s01 U28831 (.o(n25886),
	.a(dataIn_E_2_));
   in01s01 U28832 (.o(n25864),
	.a(east_input_NIB_storage_data_f_3__2_));
   ao22s01 U28833 (.o(n12078),
	.a(FE_OFN940_n24921),
	.b(n25886),
	.c(n25864),
	.d(FE_OFN24818_n24921));
   in01s01 U28834 (.o(n25888),
	.a(dataIn_E_3_));
   ao22s01 U28835 (.o(n12073),
	.a(FE_OFN940_n24921),
	.b(n25888),
	.c(n25865),
	.d(FE_OFN24824_n24921));
   in01s01 U28836 (.o(n25890),
	.a(dataIn_E_5_));
   in01s01 U28837 (.o(n25866),
	.a(east_input_NIB_storage_data_f_3__5_));
   ao22s01 U28838 (.o(n12063),
	.a(FE_OFN940_n24921),
	.b(n25890),
	.c(n25866),
	.d(FE_OFN24820_n24921));
   in01s01 U28839 (.o(n25892),
	.a(dataIn_E_14_));
   in01s01 U28840 (.o(n25867),
	.a(east_input_NIB_storage_data_f_3__14_));
   ao22s01 U28841 (.o(n12018),
	.a(FE_OFN940_n24921),
	.b(n25892),
	.c(n25867),
	.d(FE_OFN24817_n24921));
   in01s01 U28842 (.o(n25894),
	.a(dataIn_E_16_));
   in01s01 U28843 (.o(n25868),
	.a(east_input_NIB_storage_data_f_3__16_));
   ao22s01 U28844 (.o(n12008),
	.a(FE_OFN940_n24921),
	.b(n25894),
	.c(n25868),
	.d(FE_OFN24824_n24921));
   in01s01 U28845 (.o(n25870),
	.a(east_input_NIB_storage_data_f_2__0_));
   in01s01 U28846 (.o(n25871),
	.a(east_input_NIB_storage_data_f_2__2_));
   in01s01 U28847 (.o(n25872),
	.a(east_input_NIB_storage_data_f_2__3_));
   in01s01 U28848 (.o(n25873),
	.a(east_input_NIB_storage_data_f_2__5_));
   in01s01 U28849 (.o(n25874),
	.a(east_input_NIB_storage_data_f_2__14_));
   ao22f01 U28850 (.o(n11698),
	.a(FE_OFN435_n22958),
	.b(n25892),
	.c(n25874),
	.d(FE_OFN437_n22958));
   in01s01 U28851 (.o(n25875),
	.a(east_input_NIB_storage_data_f_2__16_));
   ao22f01 U28852 (.o(n11688),
	.a(FE_OFN435_n22958),
	.b(n25894),
	.c(n25875),
	.d(FE_OFN24814_n22958));
   in01s01 U28853 (.o(n25876),
	.a(east_input_NIB_storage_data_f_1__0_));
   ao22s01 U28854 (.o(n11448),
	.a(FE_OFN556_n24761),
	.b(n25884),
	.c(n25876),
	.d(n25881));
   in01s01 U28855 (.o(n25877),
	.a(east_input_NIB_storage_data_f_1__2_));
   ao22s01 U28856 (.o(n11438),
	.a(FE_OFN556_n24761),
	.b(n25886),
	.c(n25877),
	.d(n25881));
   in01s01 U28857 (.o(n25878),
	.a(east_input_NIB_storage_data_f_1__3_));
   ao22s01 U28858 (.o(n11433),
	.a(n24761),
	.b(n25888),
	.c(n25878),
	.d(n25881));
   ao22s01 U28859 (.o(n11423),
	.a(n24761),
	.b(n25890),
	.c(n25879),
	.d(n25881));
   in01s01 U28860 (.o(n25880),
	.a(east_input_NIB_storage_data_f_1__14_));
   ao22s01 U28861 (.o(n11378),
	.a(n24761),
	.b(n25892),
	.c(n25880),
	.d(n25881));
   in01s01 U28862 (.o(n25882),
	.a(east_input_NIB_storage_data_f_1__16_));
   ao22s01 U28863 (.o(n11368),
	.a(FE_OFN556_n24761),
	.b(n25894),
	.c(n25882),
	.d(n25881));
   in01s01 U28864 (.o(n25883),
	.a(east_input_NIB_storage_data_f_0__0_));
   in01s01 U28865 (.o(n25885),
	.a(east_input_NIB_storage_data_f_0__2_));
   in01s01 U28866 (.o(n25887),
	.a(east_input_NIB_storage_data_f_0__3_));
   in01s01 U28867 (.o(n25889),
	.a(east_input_NIB_storage_data_f_0__5_));
   in01s01 U28868 (.o(n25891),
	.a(east_input_NIB_storage_data_f_0__14_));
   ao22f01 U28869 (.o(n11058),
	.a(FE_OFN24862_n22945),
	.b(n25892),
	.c(n25891),
	.d(FE_OFN24861_n22945));
   ao22f01 U28870 (.o(n11048),
	.a(FE_OFN24862_n22945),
	.b(n25894),
	.c(n25893),
	.d(FE_OFN24861_n22945));
   ao22s01 U28871 (.o(n25895),
	.a(validIn_S),
	.b(n25896),
	.c(south_input_NIB_tail_ptr_f_0_),
	.d(n25897));
   no02f01 U28872 (.o(n10808),
	.a(FE_OFN5_reset),
	.b(n25895));
   no02s01 U28873 (.o(n25899),
	.a(n25897),
	.b(n25896));
   na02s01 U28874 (.o(n25898),
	.a(south_input_NIB_tail_ptr_f_1_),
	.b(FE_OFN575_n25463));
   oa12s01 U28875 (.o(n10803),
	.a(FE_OFN25785_n17770),
	.b(n25899),
	.c(n25898));
   in01s01 U28876 (.o(n25918),
	.a(dataIn_S_8_));
   in01s01 U28877 (.o(n25900),
	.a(south_input_NIB_storage_data_f_3__8_));
   ao22s01 U28878 (.o(n10758),
	.a(n20996),
	.b(n25918),
	.c(n25900),
	.d(FE_OFN896_n17769));
   in01s01 U28879 (.o(n25920),
	.a(dataIn_S_12_));
   in01s01 U28880 (.o(n25901),
	.a(south_input_NIB_storage_data_f_3__12_));
   ao22s01 U28881 (.o(n10738),
	.a(n20996),
	.b(n25920),
	.c(n25901),
	.d(n17769));
   in01s01 U28882 (.o(n25922),
	.a(dataIn_S_15_));
   in01s01 U28883 (.o(n25902),
	.a(south_input_NIB_storage_data_f_3__15_));
   ao22s01 U28884 (.o(n10723),
	.a(n20996),
	.b(n25922),
	.c(n25902),
	.d(n17769));
   in01s01 U28885 (.o(n25924),
	.a(dataIn_S_20_));
   in01s01 U28886 (.o(n25903),
	.a(south_input_NIB_storage_data_f_3__20_));
   ao22s01 U28887 (.o(n10698),
	.a(n20996),
	.b(n25924),
	.c(n25903),
	.d(n17769));
   in01s01 U28888 (.o(n25926),
	.a(dataIn_S_33_));
   in01s01 U28889 (.o(n25904),
	.a(south_input_NIB_storage_data_f_3__33_));
   ao22s01 U28890 (.o(n10633),
	.a(n20996),
	.b(n25926),
	.c(n25904),
	.d(n17769));
   in01s01 U28891 (.o(n25906),
	.a(south_input_NIB_storage_data_f_2__8_));
   in01s01 U28892 (.o(n25907),
	.a(south_input_NIB_storage_data_f_2__12_));
   ao22f01 U28893 (.o(n10418),
	.a(n20972),
	.b(n25920),
	.c(n25907),
	.d(FE_OFN84_n20972));
   in01s01 U28894 (.o(n25908),
	.a(south_input_NIB_storage_data_f_2__15_));
   in01s01 U28895 (.o(n25909),
	.a(south_input_NIB_storage_data_f_2__20_));
   ao22f01 U28896 (.o(n10378),
	.a(n20972),
	.b(n25924),
	.c(n25909),
	.d(FE_OFN84_n20972));
   in01s01 U28897 (.o(n25910),
	.a(south_input_NIB_storage_data_f_2__33_));
   ao22f01 U28898 (.o(n10313),
	.a(n20972),
	.b(n25926),
	.c(n25910),
	.d(FE_OFN84_n20972));
   in01s01 U28899 (.o(n25911),
	.a(south_input_NIB_storage_data_f_1__8_));
   ao22s01 U28900 (.o(n10118),
	.a(n20797),
	.b(n25918),
	.c(n25911),
	.d(FE_OFN25787_n17770));
   in01s01 U28901 (.o(n25912),
	.a(south_input_NIB_storage_data_f_1__12_));
   ao22s01 U28902 (.o(n10098),
	.a(n20797),
	.b(n25920),
	.c(n25912),
	.d(FE_OFN25785_n17770));
   in01s01 U28903 (.o(n25913),
	.a(south_input_NIB_storage_data_f_1__15_));
   ao22s01 U28904 (.o(n10083),
	.a(n20797),
	.b(n25922),
	.c(n25913),
	.d(FE_OFN25785_n17770));
   in01s01 U28905 (.o(n25914),
	.a(south_input_NIB_storage_data_f_1__20_));
   ao22s01 U28906 (.o(n10058),
	.a(n20797),
	.b(n25924),
	.c(n25914),
	.d(FE_OFN25787_n17770));
   in01s01 U28907 (.o(n25915),
	.a(south_input_NIB_storage_data_f_1__33_));
   ao22s01 U28908 (.o(n9993),
	.a(n20797),
	.b(n25926),
	.c(n25915),
	.d(FE_OFN25787_n17770));
   in01s01 U28909 (.o(n25917),
	.a(south_input_NIB_storage_data_f_0__8_));
   ao22s01 U28910 (.o(n9798),
	.a(FE_OFN83_n20814),
	.b(n25918),
	.c(n25917),
	.d(FE_OFN952_n25916));
   in01s01 U28911 (.o(n25919),
	.a(south_input_NIB_storage_data_f_0__12_));
   ao22s01 U28912 (.o(n9778),
	.a(FE_OFN83_n20814),
	.b(n25920),
	.c(n25919),
	.d(n25916));
   in01s01 U28913 (.o(n25921),
	.a(south_input_NIB_storage_data_f_0__15_));
   ao22s01 U28914 (.o(n9763),
	.a(FE_OFN83_n20814),
	.b(n25922),
	.c(n25921),
	.d(n25916));
   in01s01 U28915 (.o(n25923),
	.a(south_input_NIB_storage_data_f_0__20_));
   ao22s01 U28916 (.o(n9738),
	.a(FE_OFN83_n20814),
	.b(n25924),
	.c(n25923),
	.d(FE_OFN952_n25916));
   in01s01 U28917 (.o(n25925),
	.a(south_input_NIB_storage_data_f_0__33_));
   ao22s01 U28918 (.o(n9673),
	.a(FE_OFN83_n20814),
	.b(n25926),
	.c(n25925),
	.d(FE_OFN952_n25916));
   no02f01 U28919 (.o(n9518),
	.a(reset),
	.b(n25927));
   no02s01 U28920 (.o(n25931),
	.a(n25929),
	.b(n25928));
   na02s01 U28921 (.o(n25930),
	.a(west_input_NIB_tail_ptr_f_1_),
	.b(FE_OFN25598_reset));
   oa12s01 U28922 (.o(n9513),
	.a(FE_OFN381_n17772),
	.b(n25931),
	.c(n25930));
   in01s01 U28923 (.o(n25956),
	.a(dataIn_W_1_));
   in01s01 U28924 (.o(n25932),
	.a(west_input_NIB_storage_data_f_3__1_));
   in01s01 U28925 (.o(n25958),
	.a(dataIn_W_4_));
   in01s01 U28926 (.o(n25933),
	.a(west_input_NIB_storage_data_f_3__4_));
   in01s01 U28927 (.o(n25960),
	.a(dataIn_W_7_));
   in01s01 U28928 (.o(n25934),
	.a(west_input_NIB_storage_data_f_3__7_));
   in01s01 U28929 (.o(n25962),
	.a(dataIn_W_9_));
   in01s01 U28930 (.o(n25935),
	.a(west_input_NIB_storage_data_f_3__9_));
   in01s01 U28931 (.o(n25964),
	.a(dataIn_W_10_));
   in01s01 U28932 (.o(n25936),
	.a(west_input_NIB_storage_data_f_3__10_));
   in01s01 U28933 (.o(n25967),
	.a(dataIn_W_11_));
   in01s01 U28934 (.o(n25938),
	.a(west_input_NIB_storage_data_f_3__11_));
   ao22f01 U28935 (.o(n9453),
	.a(n21070),
	.b(n25967),
	.c(n25938),
	.d(FE_OFN24767_n21069));
   in01s01 U28936 (.o(n25969),
	.a(dataIn_W_17_));
   in01s01 U28937 (.o(n25939),
	.a(west_input_NIB_storage_data_f_3__17_));
   in01s01 U28938 (.o(n25940),
	.a(west_input_NIB_storage_data_f_2__1_));
   ao22f01 U28939 (.o(n9183),
	.a(n25945),
	.b(n25956),
	.c(n25940),
	.d(FE_OFN25791_n21053));
   in01s01 U28940 (.o(n25941),
	.a(west_input_NIB_storage_data_f_2__4_));
   ao22f01 U28941 (.o(n9168),
	.a(n25945),
	.b(n25958),
	.c(n25941),
	.d(FE_OFN25791_n21053));
   in01s01 U28942 (.o(n25942),
	.a(west_input_NIB_storage_data_f_2__7_));
   ao22f01 U28943 (.o(n9153),
	.a(n25945),
	.b(n25960),
	.c(n25942),
	.d(FE_OFN25791_n21053));
   ao22f01 U28944 (.o(n9143),
	.a(n25945),
	.b(n25962),
	.c(n25943),
	.d(FE_OFN25791_n21053));
   in01s01 U28945 (.o(n25944),
	.a(west_input_NIB_storage_data_f_2__10_));
   ao22f01 U28946 (.o(n9138),
	.a(n25945),
	.b(n25964),
	.c(n25944),
	.d(FE_OFN25791_n21053));
   in01s01 U28947 (.o(n25946),
	.a(west_input_NIB_storage_data_f_2__11_));
   in01s01 U28948 (.o(n25947),
	.a(west_input_NIB_storage_data_f_2__17_));
   ao22f01 U28949 (.o(n9103),
	.a(n25945),
	.b(n25969),
	.c(n25947),
	.d(FE_OFN25791_n21053));
   in01s01 U28950 (.o(n25948),
	.a(west_input_NIB_storage_data_f_1__1_));
   ao22s01 U28951 (.o(n8863),
	.a(FE_OFN380_n17772),
	.b(n25956),
	.c(n25948),
	.d(FE_OFN382_n17772));
   in01s01 U28952 (.o(n25949),
	.a(west_input_NIB_storage_data_f_1__4_));
   ao22s01 U28953 (.o(n8848),
	.a(FE_OFN380_n17772),
	.b(n25958),
	.c(n25949),
	.d(FE_OFN382_n17772));
   in01s01 U28954 (.o(n25950),
	.a(west_input_NIB_storage_data_f_1__7_));
   ao22s01 U28955 (.o(n8833),
	.a(FE_OFN380_n17772),
	.b(n25960),
	.c(n25950),
	.d(FE_OFN382_n17772));
   in01s01 U28956 (.o(n25951),
	.a(west_input_NIB_storage_data_f_1__9_));
   ao22s01 U28957 (.o(n8823),
	.a(FE_OFN380_n17772),
	.b(n25962),
	.c(n25951),
	.d(FE_OFN382_n17772));
   in01s01 U28958 (.o(n25952),
	.a(west_input_NIB_storage_data_f_1__10_));
   in01s01 U28959 (.o(n25953),
	.a(west_input_NIB_storage_data_f_1__11_));
   ao22s01 U28960 (.o(n8813),
	.a(FE_OFN380_n17772),
	.b(n25967),
	.c(n25953),
	.d(FE_OFN382_n17772));
   ao22s01 U28961 (.o(n8783),
	.a(FE_OFN380_n17772),
	.b(n25969),
	.c(n25954),
	.d(FE_OFN382_n17772));
   in01s01 U28962 (.o(n25955),
	.a(west_input_NIB_storage_data_f_0__1_));
   ao22s01 U28963 (.o(n8543),
	.a(n20855),
	.b(n25956),
	.c(n25955),
	.d(FE_OFN25750_FE_OFN24796_n20854));
   in01s01 U28964 (.o(n25957),
	.a(west_input_NIB_storage_data_f_0__4_));
   ao22s01 U28965 (.o(n8528),
	.a(n20855),
	.b(n25958),
	.c(n25957),
	.d(FE_OFN25749_FE_OFN24796_n20854));
   in01s01 U28966 (.o(n25959),
	.a(west_input_NIB_storage_data_f_0__7_));
   ao22s01 U28967 (.o(n8513),
	.a(n20855),
	.b(n25960),
	.c(n25959),
	.d(FE_OFN25750_FE_OFN24796_n20854));
   in01s01 U28968 (.o(n25961),
	.a(west_input_NIB_storage_data_f_0__9_));
   ao22s01 U28969 (.o(n8503),
	.a(n20855),
	.b(n25962),
	.c(n25961),
	.d(FE_OFN25750_FE_OFN24796_n20854));
   in01s01 U28970 (.o(n25963),
	.a(west_input_NIB_storage_data_f_0__10_));
   ao22s01 U28971 (.o(n8498),
	.a(n20855),
	.b(n25964),
	.c(n25963),
	.d(FE_OFN25749_FE_OFN24796_n20854));
   ao22s01 U28972 (.o(n8493),
	.a(n20855),
	.b(n25967),
	.c(n25966),
	.d(FE_OFN25750_FE_OFN24796_n20854));
   in01s01 U28973 (.o(n25968),
	.a(west_input_NIB_storage_data_f_0__17_));
   ao22s01 U28974 (.o(n8463),
	.a(n20855),
	.b(n25969),
	.c(n25968),
	.d(FE_OFN1101_n25965));
   ao22s01 U28975 (.o(n8228),
	.a(proc_input_NIB_tail_ptr_f_0_),
	.b(FE_OFN25843_n25972),
	.c(n25971),
	.d(n25970));
   ao22s01 U28976 (.o(n25975),
	.a(n25974),
	.b(proc_input_NIB_tail_ptr_f_1_),
	.c(n25979),
	.d(n25973));
   no02s01 U28977 (.o(n8223),
	.a(n25976),
	.b(n25975));
   in01s01 U28978 (.o(n25982),
	.a(proc_input_NIB_tail_ptr_f_3_));
   oa12s01 U28979 (.o(n8213),
	.a(n17767),
	.b(n25983),
	.c(n25982));
endmodule


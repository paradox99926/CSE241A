
module aes_sbox_4 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n48, n50, n51, n65, n68, n70, n72, n123, n142, n150, n151, n182, n187,
         n192, n226, n287, n288, n304, n305, n306, n313, n342, n398, n399,
         n400, n404, n405, n410, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842;

  AN2XD1 U28 ( .A1(n705), .A2(n704), .Z(n709) );
  OA21D1 U35 ( .A1(n691), .A2(n690), .B(n689), .Z(n696) );
  OR3D1 U88 ( .A1(n661), .A2(n793), .A3(n445), .Z(n623) );
  OA21D1 U101 ( .A1(n342), .A2(n442), .B(n604), .Z(n608) );
  OR4D1 U199 ( .A1(n646), .A2(n567), .A3(n516), .A4(n515), .Z(n518) );
  MAOI22D1 U209 ( .A1(n836), .A2(n447), .B1(n616), .B2(n757), .ZN(n509) );
  AN2XD1 U215 ( .A1(n517), .A2(n791), .Z(n516) );
  AN2XD1 U271 ( .A1(n529), .A2(n716), .Z(n466) );
  AOI21D2 U1 ( .A1(n51), .A2(a[1]), .B(n785), .ZN(n573) );
  OAI222D1 U2 ( .A1(n405), .A2(n529), .B1(n484), .B2(n735), .C1(n483), .C2(
        n739), .ZN(n488) );
  OA221D0 U3 ( .A1(n736), .A2(n48), .B1(n744), .B2(n757), .C(n50), .Z(n464) );
  INVD16 U4 ( .I(n837), .ZN(n48) );
  AOI21D1 U5 ( .A1(n70), .A2(n814), .B(n719), .ZN(n50) );
  INVD3 U6 ( .I(n736), .ZN(n782) );
  INVD0 U7 ( .I(n551), .ZN(n783) );
  OAI32D0 U8 ( .A1(n551), .A2(n741), .A3(n730), .B1(n511), .B2(n510), .ZN(n512) );
  INR4D1 U9 ( .A1(n659), .B1(n657), .B2(n658), .B3(n834), .ZN(n668) );
  OAI221D0 U10 ( .A1(n723), .A2(n716), .B1(n692), .B2(n728), .C(n583), .ZN(
        n591) );
  AOI221D1 U11 ( .A1(n814), .A2(n778), .B1(n582), .B2(n444), .C(n719), .ZN(
        n583) );
  OA222D2 U12 ( .A1(n556), .A2(n741), .B1(n555), .B2(n342), .C1(n735), .C2(
        n554), .Z(n151) );
  OAI222D1 U13 ( .A1(n765), .A2(n764), .B1(a[3]), .B2(n819), .C1(n763), .C2(
        n441), .ZN(n771) );
  AOI221D1 U14 ( .A1(n840), .A2(n444), .B1(n822), .B2(n704), .C(n522), .ZN(
        n524) );
  NR4D1 U15 ( .A1(n537), .A2(n536), .A3(n535), .A4(n534), .ZN(n538) );
  CKND2D2 U16 ( .A1(a[1]), .A2(n441), .ZN(n723) );
  OA221D1 U17 ( .A1(n730), .A2(n723), .B1(n739), .B2(n654), .C(n427), .Z(n667)
         );
  OAI221D1 U18 ( .A1(n723), .A2(n342), .B1(n730), .B2(n691), .C(n672), .ZN(
        n679) );
  OAI31D2 U19 ( .A1(n661), .A2(n65), .A3(n797), .B(n660), .ZN(n662) );
  CKAN2D4 U20 ( .A1(n439), .A2(n438), .Z(n65) );
  CKND0 U21 ( .I(n723), .ZN(n780) );
  CKND2D2 U22 ( .A1(n447), .A2(n798), .ZN(n739) );
  CKND0 U23 ( .I(a[3]), .ZN(n447) );
  ND2D3 U24 ( .A1(n437), .A2(n813), .ZN(n741) );
  OA31D0 U25 ( .A1(n692), .A2(n436), .A3(a[1]), .B(n627), .Z(n426) );
  AOI21D1 U26 ( .A1(n812), .A2(n821), .B(n830), .ZN(n655) );
  AOI221D1 U27 ( .A1(n815), .A2(n803), .B1(n801), .B2(n563), .C(n830), .ZN(
        n491) );
  OR2D0 U29 ( .A1(n708), .A2(n736), .Z(n306) );
  INVD1 U30 ( .I(n749), .ZN(n811) );
  NR2D1 U31 ( .A1(n798), .A2(n806), .ZN(n660) );
  INVD1 U32 ( .I(n733), .ZN(n801) );
  INVD2 U33 ( .I(n756), .ZN(n793) );
  INVD1 U34 ( .I(n666), .ZN(n797) );
  INVD2 U36 ( .I(a[1]), .ZN(n445) );
  ND2D0 U37 ( .A1(a[3]), .A2(n445), .ZN(n666) );
  INVD2 U38 ( .I(n692), .ZN(n827) );
  CKND3 U39 ( .I(a[0]), .ZN(n441) );
  OAI222D0 U40 ( .A1(n437), .A2(n755), .B1(n754), .B2(n753), .C1(n764), .C2(
        n752), .ZN(n762) );
  OAI222D0 U41 ( .A1(n730), .A2(n549), .B1(n404), .B2(n704), .C1(n731), .C2(
        n673), .ZN(n455) );
  AOI221D0 U42 ( .A1(n787), .A2(n532), .B1(n824), .B2(n531), .C(n530), .ZN(
        n533) );
  OAI222D0 U43 ( .A1(n729), .A2(n704), .B1(n753), .B2(n572), .C1(n734), .C2(
        n744), .ZN(n576) );
  INVD2 U44 ( .I(n437), .ZN(n818) );
  INVD2 U45 ( .I(n769), .ZN(n784) );
  NR2D1 U46 ( .A1(n65), .A2(n70), .ZN(n677) );
  ND2D2 U47 ( .A1(n437), .A2(a[6]), .ZN(n692) );
  ND2D2 U48 ( .A1(n813), .A2(n818), .ZN(n735) );
  ND2D1 U49 ( .A1(n798), .A2(n806), .ZN(n753) );
  ND2D1 U50 ( .A1(n670), .A2(n824), .ZN(n714) );
  ND2D1 U51 ( .A1(n809), .A2(n827), .ZN(n715) );
  ND2D2 U52 ( .A1(n821), .A2(n660), .ZN(n716) );
  ND2D1 U53 ( .A1(n821), .A2(n807), .ZN(n706) );
  ND2D1 U54 ( .A1(n806), .A2(n813), .ZN(n645) );
  OAI221D0 U55 ( .A1(n605), .A2(n749), .B1(n400), .B2(n744), .C(n490), .ZN(
        n493) );
  OAI222D0 U56 ( .A1(n736), .A2(n596), .B1(n595), .B2(n438), .C1(n594), .C2(
        n665), .ZN(n597) );
  INVD1 U57 ( .I(n715), .ZN(n831) );
  OAI222D0 U58 ( .A1(n742), .A2(n741), .B1(n740), .B2(n739), .C1(n439), .C2(
        n738), .ZN(n773) );
  ND2D1 U59 ( .A1(a[3]), .A2(n806), .ZN(n730) );
  INVD2 U60 ( .I(a[3]), .ZN(n446) );
  INVD1 U61 ( .I(n70), .ZN(n398) );
  CKAN2D1 U62 ( .A1(n438), .A2(n446), .Z(n51) );
  CKND1 U63 ( .I(n51), .ZN(n342) );
  INVD3 U64 ( .I(a[1]), .ZN(n444) );
  INVD2 U65 ( .I(a[0]), .ZN(n440) );
  AN2XD1 U66 ( .A1(a[3]), .A2(n434), .Z(n68) );
  AN2XD1 U67 ( .A1(n439), .A2(n444), .Z(n70) );
  ND2D1 U68 ( .A1(n435), .A2(n446), .ZN(n697) );
  ND2D1 U69 ( .A1(a[3]), .A2(n436), .ZN(n673) );
  AOI211D0 U70 ( .A1(n797), .A2(n439), .B(n68), .C(n791), .ZN(n594) );
  ND2D1 U71 ( .A1(n782), .A2(a[0]), .ZN(n551) );
  CKND2D2 U72 ( .A1(n434), .A2(n445), .ZN(n654) );
  CKND2D1 U73 ( .A1(n824), .A2(n811), .ZN(n767) );
  IIND4D2 U74 ( .A1(n72), .A2(n123), .B1(n571), .B2(n570), .ZN(d[4]) );
  OAI221D2 U75 ( .A1(n440), .A2(n142), .B1(n764), .B2(n150), .C(n151), .ZN(n72) );
  AO221D0 U76 ( .A1(n793), .A2(n823), .B1(n831), .B2(n796), .C(n541), .Z(n123)
         );
  OAI222D1 U77 ( .A1(n524), .A2(n759), .B1(n405), .B2(n615), .C1(n523), .C2(
        n704), .ZN(n536) );
  CKND2D0 U78 ( .A1(a[3]), .A2(n434), .ZN(n404) );
  OAI222D1 U79 ( .A1(n693), .A2(n716), .B1(a[0]), .B2(n533), .C1(n769), .C2(
        n758), .ZN(n534) );
  ND2D4 U80 ( .A1(n443), .A2(n438), .ZN(n769) );
  BUFFD8 U81 ( .I(n781), .Z(n438) );
  INVD2 U82 ( .I(n444), .ZN(n443) );
  ND2D1 U83 ( .A1(n789), .A2(n441), .ZN(n693) );
  OA211D1 U84 ( .A1(n690), .A2(n666), .B(n544), .C(n543), .Z(n142) );
  OA211D0 U85 ( .A1(n548), .A2(n704), .B(n547), .C(n546), .Z(n150) );
  CKND2D2 U86 ( .A1(n441), .A2(n444), .ZN(n728) );
  OAI22D1 U87 ( .A1(n728), .A2(n694), .B1(n629), .B2(n723), .ZN(n630) );
  OA222D1 U89 ( .A1(n464), .A2(n733), .B1(n673), .B2(n510), .C1(n463), .C2(
        n441), .Z(n429) );
  AOI222D1 U90 ( .A1(n789), .A2(n809), .B1(n787), .B2(n479), .C1(n783), .C2(
        n812), .ZN(n484) );
  OAI222D1 U91 ( .A1(n632), .A2(n404), .B1(n744), .B2(n746), .C1(n756), .C2(
        n631), .ZN(n633) );
  AOI221D1 U92 ( .A1(n794), .A2(n563), .B1(n562), .B2(n801), .C(n561), .ZN(
        n571) );
  ND2D1 U93 ( .A1(n443), .A2(a[0]), .ZN(n704) );
  AO31D1 U94 ( .A1(n784), .A2(n838), .A3(n670), .B(n703), .Z(n461) );
  AOI211XD0 U95 ( .A1(n842), .A2(n790), .B(n477), .C(n653), .ZN(n504) );
  OAI222D1 U96 ( .A1(n767), .A2(n572), .B1(n759), .B2(n627), .C1(n491), .C2(
        n747), .ZN(n492) );
  INVD1 U97 ( .I(n653), .ZN(n825) );
  CKND0 U98 ( .I(n728), .ZN(n779) );
  AOI221D1 U99 ( .A1(n839), .A2(n441), .B1(n831), .B2(n789), .C(n622), .ZN(
        n652) );
  AO221D1 U100 ( .A1(n835), .A2(n778), .B1(n838), .B2(n679), .C(n678), .Z(n431) );
  NR4D1 U102 ( .A1(n771), .A2(n772), .A3(n773), .A4(n770), .ZN(n774) );
  ND2D1 U103 ( .A1(n437), .A2(n806), .ZN(n712) );
  OAI222D1 U104 ( .A1(n715), .A2(n705), .B1(n685), .B2(n441), .C1(n684), .C2(
        n757), .ZN(n686) );
  AOI211XD0 U105 ( .A1(n785), .A2(n802), .B(n805), .C(n683), .ZN(n684) );
  INVD1 U106 ( .I(n753), .ZN(n807) );
  NR2D0 U107 ( .A1(n735), .A2(n753), .ZN(n680) );
  ND2D0 U108 ( .A1(n441), .A2(n438), .ZN(n747) );
  AOI22D1 U109 ( .A1(n809), .A2(n68), .B1(n787), .B2(n806), .ZN(n552) );
  AOI221D1 U110 ( .A1(n826), .A2(n441), .B1(n836), .B2(a[1]), .C(n630), .ZN(
        n631) );
  ND2D2 U111 ( .A1(n809), .A2(n821), .ZN(n708) );
  AOI221D1 U112 ( .A1(n821), .A2(n643), .B1(n824), .B2(n642), .C(n641), .ZN(
        n650) );
  INVD4 U113 ( .I(n764), .ZN(n821) );
  OA222D1 U114 ( .A1(a[0]), .A2(n668), .B1(n667), .B2(n735), .C1(n666), .C2(
        n665), .Z(n433) );
  CKND2D1 U115 ( .A1(n660), .A2(n838), .ZN(n758) );
  AN4D1 U116 ( .A1(n660), .A2(n796), .A3(n439), .A4(n824), .Z(n515) );
  ND2D2 U117 ( .A1(n784), .A2(n441), .ZN(n549) );
  AOI22D1 U118 ( .A1(n817), .A2(n787), .B1(n790), .B2(n816), .ZN(n467) );
  INVD2 U119 ( .I(n645), .ZN(n815) );
  OAI22D1 U120 ( .A1(n437), .A2(n645), .B1(n400), .B2(n712), .ZN(n450) );
  OA221D1 U121 ( .A1(n342), .A2(n664), .B1(n663), .B2(n769), .C(n662), .Z(n427) );
  AOI221D1 U122 ( .A1(n824), .A2(n459), .B1(n458), .B2(n441), .C(n457), .ZN(
        n476) );
  OAI222D1 U123 ( .A1(n792), .A2(n621), .B1(n549), .B2(n529), .C1(n528), .C2(
        n764), .ZN(n535) );
  OAI222D1 U124 ( .A1(n404), .A2(n625), .B1(n580), .B2(n579), .C1(n578), .C2(
        n741), .ZN(n581) );
  OA221D0 U125 ( .A1(n182), .A2(a[1]), .B1(n739), .B2(n187), .C(n192), .Z(n474) );
  OA21D0 U126 ( .A1(n404), .A2(n715), .B(n768), .Z(n182) );
  OA222D0 U127 ( .A1(n469), .A2(n694), .B1(n465), .B2(n692), .C1(n712), .C2(
        n713), .Z(n187) );
  OA22D1 U128 ( .A1(n467), .A2(n697), .B1(n466), .B2(n744), .Z(n192) );
  CKND1 U129 ( .I(n739), .ZN(n800) );
  IIND4D2 U130 ( .A1(n430), .A2(n431), .B1(n702), .B2(n701), .ZN(d[1]) );
  AOI221D1 U131 ( .A1(n688), .A2(n837), .B1(n68), .B2(n687), .C(n686), .ZN(
        n702) );
  OA221D1 U132 ( .A1(n733), .A2(n741), .B1(n756), .B2(n749), .C(n226), .Z(n523) );
  INVD4 U133 ( .I(n741), .ZN(n838) );
  OA221D1 U134 ( .A1(n444), .A2(n428), .B1(n588), .B2(n645), .C(n429), .Z(n475) );
  BUFFD6 U135 ( .I(a[7]), .Z(n437) );
  INVD4 U136 ( .I(n735), .ZN(n824) );
  OAI221D1 U137 ( .A1(n656), .A2(n666), .B1(n655), .B2(n654), .C(n825), .ZN(
        n658) );
  ND2D2 U138 ( .A1(n831), .A2(n441), .ZN(n627) );
  INVD2 U139 ( .I(n601), .ZN(n809) );
  OA221D0 U140 ( .A1(n600), .A2(n574), .B1(a[3]), .B2(n758), .C(n689), .Z(n226) );
  OAI222D1 U141 ( .A1(n736), .A2(n745), .B1(n677), .B2(n706), .C1(n676), .C2(
        n764), .ZN(n678) );
  AOI221D1 U142 ( .A1(n838), .A2(n634), .B1(n835), .B2(n784), .C(n633), .ZN(
        n651) );
  AOI211XD1 U143 ( .A1(n808), .A2(n577), .B(n575), .C(n576), .ZN(n578) );
  CKND1 U144 ( .I(n706), .ZN(n823) );
  OAI22D1 U145 ( .A1(n445), .A2(n706), .B1(a[1]), .B2(n626), .ZN(n628) );
  INVD4 U146 ( .I(n440), .ZN(n439) );
  CKND2D2 U147 ( .A1(n439), .A2(n434), .ZN(n744) );
  AOI221D1 U148 ( .A1(n824), .A2(n599), .B1(n598), .B2(n441), .C(n597), .ZN(
        n612) );
  AOI221D1 U149 ( .A1(n70), .A2(n671), .B1(n670), .B2(n787), .C(n669), .ZN(
        n672) );
  AOI22D1 U150 ( .A1(n793), .A2(n811), .B1(n51), .B2(n806), .ZN(n748) );
  AOI221D1 U151 ( .A1(n782), .A2(n803), .B1(n790), .B2(n810), .C(n750), .ZN(
        n765) );
  ND2D1 U152 ( .A1(n436), .A2(n446), .ZN(n752) );
  AOI221D1 U153 ( .A1(n821), .A2(n493), .B1(n783), .B2(n506), .C(n492), .ZN(
        n502) );
  CKND1 U154 ( .I(n767), .ZN(n826) );
  OR2D0 U155 ( .A1(n621), .A2(n744), .Z(n287) );
  OR2D0 U156 ( .A1(n432), .A2(n769), .Z(n288) );
  ND3D1 U157 ( .A1(n287), .A2(n288), .A3(n433), .ZN(n430) );
  CKND0 U158 ( .I(n680), .ZN(n432) );
  CKAN2D1 U159 ( .A1(n462), .A2(n789), .Z(n304) );
  AN2D1 U160 ( .A1(n831), .A2(n796), .Z(n305) );
  NR3D1 U161 ( .A1(n304), .A2(n305), .A3(n461), .ZN(n463) );
  OR2XD1 U162 ( .A1(n438), .A2(n714), .Z(n313) );
  CKND2D2 U163 ( .A1(n306), .A2(n313), .ZN(n653) );
  ND2D3 U164 ( .A1(n445), .A2(n438), .ZN(n736) );
  AOI221D1 U165 ( .A1(n780), .A2(n675), .B1(n812), .B2(n65), .C(n674), .ZN(
        n676) );
  INVD6 U166 ( .I(n436), .ZN(n806) );
  AOI221D1 U167 ( .A1(n801), .A2(n779), .B1(n810), .B2(n789), .C(n553), .ZN(
        n554) );
  INVD6 U168 ( .I(n435), .ZN(n798) );
  ND2D2 U169 ( .A1(a[6]), .A2(n818), .ZN(n764) );
  ND2D2 U170 ( .A1(a[6]), .A2(n806), .ZN(n757) );
  OAI211D0 U171 ( .A1(n806), .A2(n739), .B(n756), .C(n734), .ZN(n671) );
  AOI221D1 U172 ( .A1(n783), .A2(n829), .B1(n778), .B2(n842), .C(n581), .ZN(
        n614) );
  AOI21D0 U173 ( .A1(n673), .A2(n749), .B(n410), .ZN(n669) );
  OAI22D0 U174 ( .A1(n749), .A2(n759), .B1(a[1]), .B2(n748), .ZN(n750) );
  ND2D2 U175 ( .A1(n436), .A2(n798), .ZN(n749) );
  ND2D2 U176 ( .A1(a[3]), .A2(n438), .ZN(n756) );
  AOI221D1 U177 ( .A1(n795), .A2(n591), .B1(n821), .B2(n590), .C(n589), .ZN(
        n613) );
  CKND2D0 U178 ( .A1(n435), .A2(a[3]), .ZN(n399) );
  CKND2D0 U179 ( .A1(n435), .A2(a[3]), .ZN(n400) );
  CKND2D0 U180 ( .A1(n439), .A2(n438), .ZN(n410) );
  AOI211XD0 U181 ( .A1(n822), .A2(n439), .B(n628), .C(n832), .ZN(n632) );
  AOI211XD0 U182 ( .A1(n820), .A2(n790), .B(n482), .C(n481), .ZN(n483) );
  CKND2D0 U183 ( .A1(n439), .A2(n438), .ZN(n405) );
  ND2D0 U184 ( .A1(n780), .A2(n838), .ZN(n510) );
  CKND2D0 U185 ( .A1(n435), .A2(a[3]), .ZN(n734) );
  CKND2D0 U186 ( .A1(n434), .A2(n723), .ZN(n721) );
  ND2D0 U187 ( .A1(n439), .A2(n787), .ZN(n713) );
  NR2D0 U188 ( .A1(n615), .A2(n398), .ZN(n751) );
  NR2D0 U189 ( .A1(n789), .A2(n778), .ZN(n604) );
  CKND2D0 U190 ( .A1(n673), .A2(n733), .ZN(n675) );
  ND2D0 U191 ( .A1(n806), .A2(n818), .ZN(n600) );
  CKND2D0 U192 ( .A1(n810), .A2(n827), .ZN(n746) );
  CKND2D0 U193 ( .A1(n801), .A2(n827), .ZN(n596) );
  ND2D0 U194 ( .A1(n434), .A2(n446), .ZN(n759) );
  NR2XD0 U195 ( .A1(n839), .A2(n506), .ZN(n507) );
  CKND2D0 U196 ( .A1(n443), .A2(n434), .ZN(n731) );
  ND2D0 U197 ( .A1(n436), .A2(n818), .ZN(n694) );
  ND2D0 U198 ( .A1(n434), .A2(n798), .ZN(n616) );
  ND2D0 U200 ( .A1(n436), .A2(n813), .ZN(n505) );
  INR2D1 U201 ( .A1(n745), .B1(n495), .ZN(n496) );
  CKND2D0 U202 ( .A1(a[1]), .A2(a[6]), .ZN(n480) );
  OAI31D0 U203 ( .A1(n782), .A2(n70), .A3(n793), .B(n839), .ZN(n485) );
  AOI22D0 U204 ( .A1(n840), .A2(n784), .B1(n796), .B2(n826), .ZN(n543) );
  NR2D0 U205 ( .A1(n442), .A2(n743), .ZN(n726) );
  NR2D0 U206 ( .A1(n786), .A2(n782), .ZN(n469) );
  CKND2D0 U207 ( .A1(n713), .A2(n723), .ZN(n577) );
  AOI21D0 U208 ( .A1(n836), .A2(n796), .B(n682), .ZN(n685) );
  NR2D0 U210 ( .A1(n65), .A2(n779), .ZN(n605) );
  ND2D0 U211 ( .A1(n793), .A2(n833), .ZN(n557) );
  CKND0 U212 ( .I(n758), .ZN(n839) );
  NR2D0 U213 ( .A1(n793), .A2(n786), .ZN(n449) );
  CKND0 U214 ( .I(n572), .ZN(n794) );
  CKND2D0 U216 ( .A1(n443), .A2(a[3]), .ZN(n766) );
  ND3D0 U217 ( .A1(n68), .A2(n660), .A3(n824), .ZN(n743) );
  OAI22D0 U218 ( .A1(n739), .A2(n736), .B1(n644), .B2(n723), .ZN(n514) );
  CKND2D0 U219 ( .A1(n766), .A2(n342), .ZN(n519) );
  NR2D0 U220 ( .A1(n715), .A2(a[3]), .ZN(n682) );
  NR2D0 U221 ( .A1(n804), .A2(n809), .ZN(n592) );
  AOI22D0 U222 ( .A1(n441), .A2(n796), .B1(n447), .B2(n786), .ZN(n580) );
  AOI22D0 U223 ( .A1(n789), .A2(a[0]), .B1(a[1]), .B2(n68), .ZN(n478) );
  NR2D0 U224 ( .A1(n68), .A2(n802), .ZN(n644) );
  NR2D0 U225 ( .A1(n743), .A2(n439), .ZN(n699) );
  ND2D0 U226 ( .A1(n795), .A2(a[1]), .ZN(n705) );
  NR2D0 U227 ( .A1(n626), .A2(n707), .ZN(n725) );
  CKND2D0 U228 ( .A1(n841), .A2(n803), .ZN(n768) );
  ND2D0 U229 ( .A1(n809), .A2(n838), .ZN(n665) );
  CKND2D0 U230 ( .A1(n779), .A2(n446), .ZN(n707) );
  ND2D0 U231 ( .A1(n801), .A2(n841), .ZN(n745) );
  CKND2D0 U232 ( .A1(n800), .A2(n824), .ZN(n659) );
  CKND2D0 U233 ( .A1(n814), .A2(n803), .ZN(n529) );
  CKND2D0 U234 ( .A1(n766), .A2(n549), .ZN(n550) );
  NR2D0 U235 ( .A1(n836), .A2(n680), .ZN(n452) );
  NR2D0 U236 ( .A1(n703), .A2(n836), .ZN(n710) );
  OAI21D0 U237 ( .A1(a[0]), .A2(n673), .B(n733), .ZN(n479) );
  CKND2D1 U238 ( .A1(n486), .A2(n485), .ZN(n487) );
  AOI211XD0 U239 ( .A1(n838), .A2(n489), .B(n488), .C(n487), .ZN(n503) );
  OAI22D0 U240 ( .A1(n441), .A2(n706), .B1(n445), .B2(n716), .ZN(n522) );
  ND2D0 U241 ( .A1(n65), .A2(n811), .ZN(n635) );
  OAI21D0 U242 ( .A1(n735), .A2(n601), .B(n706), .ZN(n582) );
  AOI22D0 U243 ( .A1(n790), .A2(n837), .B1(n782), .B2(n816), .ZN(n560) );
  AOI21D0 U244 ( .A1(n840), .A2(n68), .B(n834), .ZN(n558) );
  NR2XD0 U245 ( .A1(n816), .A2(n827), .ZN(n629) );
  OAI33D0 U246 ( .A1(n739), .A2(n438), .A3(n712), .B1(n645), .B2(a[1]), .B3(
        n644), .ZN(n648) );
  NR2XD0 U247 ( .A1(n822), .A2(n833), .ZN(n656) );
  NR2D0 U248 ( .A1(n811), .A2(n793), .ZN(n511) );
  OAI22D0 U249 ( .A1(n769), .A2(n768), .B1(n767), .B2(n766), .ZN(n770) );
  AOI21D0 U250 ( .A1(n342), .A2(n574), .B(n398), .ZN(n453) );
  OAI22D0 U251 ( .A1(n749), .A2(n342), .B1(n677), .B2(n697), .ZN(n454) );
  OAI31D0 U252 ( .A1(n723), .A2(n802), .A3(n735), .B(n722), .ZN(n727) );
  AOI31D0 U253 ( .A1(n827), .A2(n721), .A3(n802), .B(n720), .ZN(n722) );
  AOI32D0 U254 ( .A1(n782), .A2(n441), .A3(n812), .B1(n780), .B2(n545), .ZN(
        n547) );
  CKND2D0 U255 ( .A1(n400), .A2(n729), .ZN(n545) );
  NR2D0 U256 ( .A1(n616), .A2(n704), .ZN(n688) );
  OAI21D0 U257 ( .A1(n399), .A2(n600), .B(n625), .ZN(n506) );
  AOI21D0 U258 ( .A1(n601), .A2(n645), .B(n342), .ZN(n495) );
  INR2D0 U259 ( .A1(n517), .B1(n654), .ZN(n698) );
  CKND2D0 U260 ( .A1(n807), .A2(n827), .ZN(n625) );
  AOI22D0 U261 ( .A1(n815), .A2(n732), .B1(n817), .B2(n787), .ZN(n740) );
  CKND2D0 U262 ( .A1(n747), .A2(n744), .ZN(n732) );
  ND2D0 U263 ( .A1(n438), .A2(n798), .ZN(n548) );
  NR2D0 U264 ( .A1(n505), .A2(n654), .ZN(n562) );
  CKND2D0 U265 ( .A1(n670), .A2(n827), .ZN(n621) );
  CKND0 U266 ( .I(n690), .ZN(n841) );
  CKND2D0 U267 ( .A1(n809), .A2(n444), .ZN(n664) );
  CKND2D0 U268 ( .A1(n811), .A2(n818), .ZN(n615) );
  CKND2D0 U269 ( .A1(n68), .A2(n798), .ZN(n593) );
  NR2D0 U270 ( .A1(n840), .A2(n826), .ZN(n460) );
  OAI22D0 U272 ( .A1(n456), .A2(n764), .B1(n731), .B2(n625), .ZN(n457) );
  AOI21D0 U273 ( .A1(n759), .A2(n729), .B(n764), .ZN(n617) );
  AOI21D0 U274 ( .A1(n835), .A2(a[1]), .B(n680), .ZN(n681) );
  ND4D0 U275 ( .A1(n70), .A2(n815), .A3(n435), .A4(n437), .ZN(n711) );
  AOI32D0 U276 ( .A1(n436), .A2(n441), .A3(n796), .B1(n807), .B2(n623), .ZN(
        n624) );
  AOI31D0 U277 ( .A1(n434), .A2(n806), .A3(n70), .B(n805), .ZN(n490) );
  CKND2D1 U278 ( .A1(n586), .A2(n585), .ZN(n590) );
  AOI21D0 U279 ( .A1(n788), .A2(n824), .B(n562), .ZN(n508) );
  NR2D0 U280 ( .A1(n791), .A2(a[3]), .ZN(n607) );
  CKND2D1 U281 ( .A1(n437), .A2(n494), .ZN(n497) );
  AOI21D0 U282 ( .A1(n801), .A2(n837), .B(n682), .ZN(n498) );
  NR2D0 U283 ( .A1(n791), .A2(n789), .ZN(n465) );
  AOI22D0 U284 ( .A1(n804), .A2(n779), .B1(n802), .B2(n434), .ZN(n564) );
  CKND2D0 U285 ( .A1(n704), .A2(n446), .ZN(n565) );
  CKND0 U286 ( .I(n751), .ZN(n819) );
  AOI22D0 U287 ( .A1(n784), .A2(n815), .B1(n793), .B2(n798), .ZN(n755) );
  OAI211D0 U288 ( .A1(n436), .A2(n766), .B(n616), .C(n733), .ZN(n531) );
  OAI33D0 U289 ( .A1(n404), .A2(n437), .A3(n753), .B1(n690), .B2(n438), .B3(
        n399), .ZN(n530) );
  OAI32D0 U290 ( .A1(n752), .A2(n469), .A3(n692), .B1(n468), .B2(n723), .ZN(
        n472) );
  AOI31D0 U291 ( .A1(n435), .A2(n813), .A3(n793), .B(n682), .ZN(n468) );
  AOI211D0 U292 ( .A1(n760), .A2(n645), .B(n574), .C(n398), .ZN(n470) );
  NR2D0 U293 ( .A1(a[3]), .A2(n436), .ZN(n670) );
  OAI31D0 U294 ( .A1(n731), .A2(n760), .A3(n733), .B(n603), .ZN(n610) );
  AOI33D0 U295 ( .A1(n602), .A2(n813), .A3(n784), .B1(n833), .B2(n446), .B3(
        n780), .ZN(n603) );
  OAI22D0 U296 ( .A1(a[3]), .A2(n601), .B1(n441), .B2(n600), .ZN(n602) );
  CKND0 U297 ( .I(n600), .ZN(n820) );
  OAI33D0 U298 ( .A1(n645), .A2(n439), .A3(n438), .B1(n480), .B2(n712), .B3(
        n744), .ZN(n481) );
  OAI22D0 U299 ( .A1(n813), .A2(n697), .B1(n798), .B2(n645), .ZN(n637) );
  AOI32D0 U300 ( .A1(n437), .A2(n798), .A3(n782), .B1(n787), .B2(n450), .ZN(
        n451) );
  CKND2D0 U301 ( .A1(n435), .A2(n438), .ZN(n574) );
  AOI21D0 U302 ( .A1(n715), .A2(n659), .B(n434), .ZN(n618) );
  AOI21D0 U303 ( .A1(n826), .A2(n68), .B(n737), .ZN(n738) );
  OAI33D0 U304 ( .A1(n736), .A2(n735), .A3(n399), .B1(n757), .B2(n438), .B3(
        n733), .ZN(n737) );
  NR2D0 U305 ( .A1(n779), .A2(n787), .ZN(n639) );
  AOI21D0 U306 ( .A1(n778), .A2(n637), .B(n636), .ZN(n640) );
  CKND2D1 U307 ( .A1(n757), .A2(n712), .ZN(n563) );
  OAI21D0 U308 ( .A1(n696), .A2(n723), .B(n695), .ZN(n700) );
  OA33D0 U309 ( .A1(n694), .A2(n399), .A3(n398), .B1(n693), .B2(n692), .B3(
        n752), .Z(n695) );
  CKND2D0 U310 ( .A1(n680), .A2(n728), .ZN(n424) );
  NR2D0 U311 ( .A1(n435), .A2(n813), .ZN(n462) );
  CKND2D0 U312 ( .A1(n436), .A2(a[6]), .ZN(n760) );
  AOI32D0 U313 ( .A1(n435), .A2(n818), .A3(n795), .B1(n68), .B2(n542), .ZN(
        n544) );
  OAI22D0 U314 ( .A1(a[6]), .A2(n435), .B1(n436), .B2(n741), .ZN(n542) );
  BUFFD4 U315 ( .I(a[5]), .Z(n436) );
  BUFFD4 U316 ( .I(a[4]), .Z(n435) );
  BUFFD4 U317 ( .I(a[2]), .Z(n434) );
  INVD1 U318 ( .I(n549), .ZN(n785) );
  INVD1 U319 ( .I(n557), .ZN(n834) );
  NR2D1 U320 ( .A1(n442), .A2(a[3]), .ZN(n661) );
  INVD1 U321 ( .I(n704), .ZN(n778) );
  INVD1 U322 ( .I(n766), .ZN(n796) );
  INVD1 U323 ( .I(n693), .ZN(n790) );
  INVD1 U324 ( .I(n665), .ZN(n840) );
  INVD1 U325 ( .I(n713), .ZN(n788) );
  INVD1 U326 ( .I(n768), .ZN(n842) );
  AOI222D0 U327 ( .A1(n789), .A2(n803), .B1(n801), .B2(n65), .C1(n810), .C2(
        n787), .ZN(n546) );
  INVD1 U328 ( .I(n579), .ZN(n836) );
  ND2D1 U329 ( .A1(n793), .A2(a[1]), .ZN(n572) );
  AO221D0 U330 ( .A1(n782), .A2(n812), .B1(n780), .B2(n795), .C(n688), .Z(n642) );
  INVD1 U331 ( .I(n747), .ZN(n786) );
  INVD1 U332 ( .I(n587), .ZN(n830) );
  INVD1 U333 ( .I(n625), .ZN(n835) );
  INVD1 U334 ( .I(n708), .ZN(n822) );
  INVD1 U335 ( .I(n626), .ZN(n833) );
  ND2D1 U336 ( .A1(n778), .A2(n804), .ZN(n588) );
  OAI22D1 U337 ( .A1(n398), .A2(n739), .B1(n592), .B2(n728), .ZN(n599) );
  ND2D1 U338 ( .A1(n799), .A2(n815), .ZN(n689) );
  INVD1 U339 ( .I(n730), .ZN(n808) );
  INVD1 U340 ( .I(n548), .ZN(n799) );
  INVD1 U341 ( .I(n596), .ZN(n828) );
  AOI221D0 U342 ( .A1(n785), .A2(n812), .B1(n807), .B2(n550), .C(n688), .ZN(
        n556) );
  INVD1 U343 ( .I(a[0]), .ZN(n442) );
  OAI222D0 U344 ( .A1(n626), .A2(n438), .B1(n600), .B2(n593), .C1(a[3]), .C2(
        n706), .ZN(n598) );
  OAI222D0 U345 ( .A1(n744), .A2(n752), .B1(n766), .B2(n635), .C1(n733), .C2(
        n693), .ZN(n643) );
  NR2D1 U346 ( .A1(n636), .A2(n751), .ZN(n595) );
  NR4D0 U347 ( .A1(n443), .A2(n818), .A3(n747), .A4(n739), .ZN(n683) );
  NR4D0 U348 ( .A1(n697), .A2(n747), .A3(n741), .A4(n806), .ZN(n720) );
  OAI222D0 U349 ( .A1(n404), .A2(n708), .B1(n580), .B2(n716), .C1(n626), .C2(
        n654), .ZN(n477) );
  OAI222D0 U350 ( .A1(n741), .A2(n616), .B1(a[3]), .B2(n615), .C1(n735), .C2(
        n752), .ZN(n619) );
  NR4D0 U351 ( .A1(n753), .A2(n741), .A3(n654), .A4(a[3]), .ZN(n724) );
  NR2D1 U352 ( .A1(n690), .A2(n728), .ZN(n719) );
  OAI32D1 U353 ( .A1(n574), .A2(n728), .A3(n673), .B1(n573), .B2(n749), .ZN(
        n575) );
  OAI222D0 U354 ( .A1(n654), .A2(n752), .B1(a[0]), .B2(n552), .C1(n734), .C2(
        n551), .ZN(n553) );
  ND2D1 U355 ( .A1(n827), .A2(n811), .ZN(n626) );
  OAI222D0 U356 ( .A1(n736), .A2(n673), .B1(n478), .B2(n749), .C1(a[1]), .C2(
        n400), .ZN(n489) );
  INVD1 U357 ( .I(n759), .ZN(n795) );
  NR4D0 U358 ( .A1(n527), .A2(n526), .A3(n525), .A4(n584), .ZN(n528) );
  NR3D0 U359 ( .A1(n723), .A2(a[3]), .A3(n749), .ZN(n526) );
  NR4D0 U360 ( .A1(n569), .A2(n568), .A3(n567), .A4(n724), .ZN(n570) );
  INVD1 U361 ( .I(n697), .ZN(n803) );
  OAI222D0 U362 ( .A1(n747), .A2(n746), .B1(n745), .B2(n744), .C1(a[1]), .C2(
        n743), .ZN(n772) );
  INVD1 U363 ( .I(n752), .ZN(n812) );
  INVD1 U364 ( .I(n654), .ZN(n787) );
  INVD1 U365 ( .I(n673), .ZN(n810) );
  INVD1 U366 ( .I(n712), .ZN(n837) );
  INVD1 U367 ( .I(n400), .ZN(n802) );
  NR3D0 U368 ( .A1(n505), .A2(n399), .A3(n769), .ZN(n471) );
  OAI222D0 U369 ( .A1(n560), .A2(n697), .B1(n559), .B2(n398), .C1(a[1]), .C2(
        n558), .ZN(n561) );
  AOI21D1 U370 ( .A1(n799), .A2(n841), .B(n828), .ZN(n559) );
  INVD1 U371 ( .I(n731), .ZN(n789) );
  ND2D1 U372 ( .A1(a[3]), .A2(n798), .ZN(n733) );
  NR2D1 U373 ( .A1(n694), .A2(n697), .ZN(n703) );
  INVD1 U374 ( .I(n505), .ZN(n814) );
  INVD1 U375 ( .I(n691), .ZN(n804) );
  AOI221D0 U376 ( .A1(n778), .A2(n51), .B1(n783), .B2(n808), .C(n584), .ZN(
        n585) );
  NR4D0 U377 ( .A1(n455), .A2(n454), .A3(n525), .A4(n453), .ZN(n456) );
  ND2D1 U378 ( .A1(n808), .A2(n827), .ZN(n587) );
  INVD1 U379 ( .I(n627), .ZN(n832) );
  INVD1 U380 ( .I(n721), .ZN(n792) );
  OAI222D0 U381 ( .A1(n434), .A2(n640), .B1(n639), .B2(n768), .C1(n638), .C2(
        n767), .ZN(n641) );
  NR3D0 U382 ( .A1(n661), .A2(n782), .A3(n795), .ZN(n638) );
  OAI221D0 U383 ( .A1(n399), .A2(n736), .B1(n697), .B2(n769), .C(n624), .ZN(
        n634) );
  AOI222D0 U384 ( .A1(n784), .A2(n800), .B1(n802), .B2(n786), .C1(n788), .C2(
        n436), .ZN(n586) );
  NR2XD0 U385 ( .A1(n762), .A2(n761), .ZN(n763) );
  OAI222D0 U386 ( .A1(n498), .A2(n728), .B1(n798), .B2(n497), .C1(n496), .C2(
        n704), .ZN(n500) );
  OAI222D0 U387 ( .A1(n566), .A2(n758), .B1(n767), .B2(n565), .C1(n564), .C2(
        n760), .ZN(n569) );
  NR4D0 U388 ( .A1(n673), .A2(n736), .A3(n764), .A4(n798), .ZN(n646) );
  OAI221D0 U389 ( .A1(n449), .A2(n601), .B1(n759), .B2(n704), .C(n448), .ZN(
        n459) );
  OAI221D0 U390 ( .A1(n452), .A2(n404), .B1(n756), .B2(n716), .C(n451), .ZN(
        n458) );
  OAI221D0 U391 ( .A1(n441), .A2(n716), .B1(n692), .B2(n704), .C(n681), .ZN(
        n687) );
  OAI221D0 U392 ( .A1(a[1]), .A2(n659), .B1(n707), .B2(n665), .C(n521), .ZN(
        n537) );
  AOI221D0 U393 ( .A1(n719), .A2(n795), .B1(n51), .B2(n718), .C(n717), .ZN(
        n776) );
  OAI221D0 U394 ( .A1(n723), .A2(n712), .B1(n443), .B2(n767), .C(n711), .ZN(
        n718) );
  NR3D0 U395 ( .A1(n723), .A2(n435), .A3(n600), .ZN(n636) );
  NR4D0 U396 ( .A1(n439), .A2(n813), .A3(n753), .A4(n759), .ZN(n568) );
  NR3D0 U397 ( .A1(n759), .A2(n437), .A3(n435), .ZN(n657) );
  NR3D0 U398 ( .A1(n442), .A2(n435), .A3(n673), .ZN(n584) );
  NR3D0 U399 ( .A1(n692), .A2(n806), .A3(n697), .ZN(n517) );
  ND2D1 U400 ( .A1(n436), .A2(n437), .ZN(n690) );
  OAI222D0 U401 ( .A1(a[1]), .A2(n760), .B1(n728), .B2(n741), .C1(n735), .C2(
        n731), .ZN(n482) );
  NR3D0 U402 ( .A1(n705), .A2(n435), .A3(n818), .ZN(n647) );
  AN3XD1 U403 ( .A1(n424), .A2(n425), .A3(n426), .Z(n555) );
  ND2D0 U404 ( .A1(a[1]), .A2(n833), .ZN(n425) );
  INVD1 U405 ( .I(n757), .ZN(n816) );
  ND2D1 U406 ( .A1(n434), .A2(n436), .ZN(n729) );
  ND2D1 U407 ( .A1(n435), .A2(n806), .ZN(n601) );
  INVD1 U408 ( .I(n434), .ZN(n781) );
  OAI222D0 U409 ( .A1(n608), .A2(n758), .B1(n607), .B2(n708), .C1(n606), .C2(
        n739), .ZN(n609) );
  OA22D0 U410 ( .A1(n760), .A2(n398), .B1(n712), .B2(n605), .Z(n606) );
  OAI222D0 U411 ( .A1(n509), .A2(n398), .B1(n508), .B2(n400), .C1(n507), .C2(
        n747), .ZN(n513) );
  INVD1 U412 ( .I(n760), .ZN(n817) );
  ND2D1 U413 ( .A1(n435), .A2(n434), .ZN(n691) );
  OAI22D1 U414 ( .A1(n445), .A2(n621), .B1(n620), .B2(n398), .ZN(n622) );
  NR4D0 U415 ( .A1(n619), .A2(n618), .A3(n828), .A4(n617), .ZN(n620) );
  NR4D0 U416 ( .A1(a[6]), .A2(n447), .A3(n712), .A4(n744), .ZN(n499) );
  ND4D1 U417 ( .A1(n614), .A2(n613), .A3(n612), .A4(n611), .ZN(d[3]) );
  NR2D1 U418 ( .A1(n610), .A2(n609), .ZN(n611) );
  ND4D1 U419 ( .A1(n502), .A2(n503), .A3(n504), .A4(n501), .ZN(d[6]) );
  NR4D0 U420 ( .A1(n500), .A2(n499), .A3(n515), .A4(n516), .ZN(n501) );
  ND4D1 U421 ( .A1(n476), .A2(n475), .A3(n474), .A4(n473), .ZN(d[7]) );
  NR4D0 U422 ( .A1(n472), .A2(n471), .A3(n699), .A4(n470), .ZN(n473) );
  ND4D1 U423 ( .A1(n652), .A2(n651), .A3(n650), .A4(n649), .ZN(d[2]) );
  NR4D0 U424 ( .A1(n648), .A2(n647), .A3(n646), .A4(n726), .ZN(n649) );
  NR4D0 U425 ( .A1(n727), .A2(n726), .A3(n725), .A4(n724), .ZN(n775) );
  ND3D1 U426 ( .A1(n540), .A2(n539), .A3(n538), .ZN(d[5]) );
  AOI211D1 U427 ( .A1(n841), .A2(n514), .B(n513), .C(n512), .ZN(n540) );
  INR4D0 U428 ( .A1(n743), .B1(n518), .B2(n725), .B3(n698), .ZN(n539) );
  NR4D0 U429 ( .A1(n700), .A2(n720), .A3(n699), .A4(n698), .ZN(n701) );
  INVD2 U430 ( .I(a[6]), .ZN(n813) );
  OAI222D0 U431 ( .A1(n710), .A2(n410), .B1(n709), .B2(n708), .C1(n707), .C2(
        n706), .ZN(n777) );
  OAI222D0 U432 ( .A1(n410), .A2(n587), .B1(n716), .B2(n666), .C1(n626), .C2(
        n744), .ZN(n541) );
  OAI222D0 U433 ( .A1(n712), .A2(n588), .B1(n405), .B2(n746), .C1(n604), .C2(
        n587), .ZN(n589) );
  ND2D1 U434 ( .A1(n410), .A2(n736), .ZN(n520) );
  OAI222D0 U435 ( .A1(n410), .A2(n733), .B1(n677), .B2(n673), .C1(n739), .C2(
        n549), .ZN(n527) );
  NR3D0 U436 ( .A1(n806), .A2(n443), .A3(n405), .ZN(n525) );
  OA221D0 U437 ( .A1(n460), .A2(n759), .B1(n706), .B2(n756), .C(n557), .Z(n428) );
  INVD1 U438 ( .I(n588), .ZN(n805) );
  NR3D0 U439 ( .A1(n704), .A2(n798), .A3(n714), .ZN(n567) );
  OAI21D0 U440 ( .A1(n645), .A2(n733), .B(n714), .ZN(n532) );
  AOI31D1 U441 ( .A1(n716), .A2(n715), .A3(n714), .B(n713), .ZN(n717) );
  IND4D1 U442 ( .A1(n777), .B1(n776), .B2(n775), .B3(n774), .ZN(d[0]) );
  NR2D1 U443 ( .A1(n785), .A2(n788), .ZN(n566) );
  OAI31D0 U444 ( .A1(n446), .A2(n785), .A3(n791), .B(n680), .ZN(n486) );
  OAI222D0 U445 ( .A1(n760), .A2(n769), .B1(n759), .B2(n758), .C1(n757), .C2(
        n756), .ZN(n761) );
  OAI22D0 U446 ( .A1(n404), .A2(n398), .B1(n728), .B2(n756), .ZN(n494) );
  NR2XD0 U447 ( .A1(n812), .A2(n808), .ZN(n663) );
  AOI22D0 U448 ( .A1(n831), .A2(n520), .B1(n680), .B2(n519), .ZN(n521) );
  OA222D0 U449 ( .A1(n731), .A2(n730), .B1(n729), .B2(n728), .C1(n733), .C2(
        n398), .Z(n742) );
  OAI22D0 U450 ( .A1(n730), .A2(n736), .B1(n749), .B2(n769), .ZN(n674) );
  AOI21D0 U451 ( .A1(a[3]), .A2(n838), .B(n797), .ZN(n754) );
  ND2D1 U452 ( .A1(n660), .A2(n827), .ZN(n579) );
  AOI22D0 U453 ( .A1(n808), .A2(n787), .B1(n784), .B2(n810), .ZN(n448) );
  INVD1 U454 ( .I(n621), .ZN(n829) );
  INVD1 U455 ( .I(n744), .ZN(n791) );
endmodule


module aes_sbox_3 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n48, n51, n53, n68, n70, n72, n187, n226, n310, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861;

  AN2XD1 U28 ( .A1(n721), .A2(n720), .Z(n725) );
  OA21D1 U35 ( .A1(n705), .A2(n704), .B(n703), .Z(n710) );
  OR3D1 U88 ( .A1(n673), .A2(n310), .A3(n445), .Z(n635) );
  OR4D1 U199 ( .A1(n658), .A2(n577), .A3(n522), .A4(n521), .Z(n524) );
  MAOI22D1 U209 ( .A1(n855), .A2(n447), .B1(n628), .B2(n775), .ZN(n515) );
  AN2XD1 U215 ( .A1(n523), .A2(n810), .Z(n522) );
  AN2XD1 U271 ( .A1(n536), .A2(n733), .Z(n469) );
  AO31D1 U286 ( .A1(n803), .A2(n857), .A3(n683), .B(n719), .Z(n462) );
  AO21D1 U297 ( .A1(n427), .A2(n833), .B(n736), .Z(n461) );
  OAI221D1 U1 ( .A1(n440), .A2(n733), .B1(n706), .B2(n720), .C(n695), .ZN(n701) );
  ND2D1 U2 ( .A1(n830), .A2(n837), .ZN(n627) );
  ND2D1 U3 ( .A1(n433), .A2(a[3]), .ZN(n752) );
  CKBD4 U4 ( .I(a[4]), .Z(n433) );
  OAI222D1 U5 ( .A1(n811), .A2(n633), .B1(n556), .B2(n536), .C1(n535), .C2(
        n782), .ZN(n542) );
  AOI221D2 U6 ( .A1(n694), .A2(n746), .B1(n442), .B2(n852), .C(n558), .ZN(n562) );
  CKND3 U7 ( .I(n439), .ZN(n437) );
  CKND4 U8 ( .I(a[0]), .ZN(n439) );
  NR2D1 U9 ( .A1(n441), .A2(a[3]), .ZN(n673) );
  CKND1 U10 ( .I(n437), .ZN(n441) );
  OAI222D1 U11 ( .A1(n726), .A2(n536), .B1(n490), .B2(n753), .C1(n489), .C2(
        n757), .ZN(n494) );
  AOI211D1 U12 ( .A1(n839), .A2(n809), .B(n488), .C(n487), .ZN(n489) );
  OAI222D1 U13 ( .A1(n644), .A2(n226), .B1(n762), .B2(n764), .C1(n643), .C2(
        n774), .ZN(n645) );
  AOI221D1 U14 ( .A1(n857), .A2(n646), .B1(n854), .B2(n803), .C(n645), .ZN(
        n663) );
  OAI31D1 U15 ( .A1(n706), .A2(n434), .A3(n442), .B(n639), .ZN(n558) );
  ND2D1 U16 ( .A1(n850), .A2(n440), .ZN(n639) );
  OAI31D2 U17 ( .A1(n673), .A2(n800), .A3(n816), .B(n672), .ZN(n674) );
  OAI22D1 U18 ( .A1(n445), .A2(n633), .B1(n632), .B2(n745), .ZN(n634) );
  AOI221D0 U19 ( .A1(n840), .A2(n655), .B1(n843), .B2(n654), .C(n653), .ZN(
        n662) );
  ND2D0 U20 ( .A1(n840), .A2(n672), .ZN(n733) );
  INVD2 U21 ( .I(n782), .ZN(n840) );
  ND2D1 U22 ( .A1(n310), .A2(n442), .ZN(n584) );
  AOI211XD0 U23 ( .A1(n860), .A2(n520), .B(n519), .C(n518), .ZN(n547) );
  OAI222D1 U24 ( .A1(n531), .A2(n777), .B1(n726), .B2(n627), .C1(n720), .C2(
        n530), .ZN(n543) );
  AOI211XD1 U25 ( .A1(n827), .A2(n589), .B(n587), .C(n588), .ZN(n590) );
  ND2D2 U26 ( .A1(n434), .A2(n817), .ZN(n767) );
  ND2D1 U27 ( .A1(n846), .A2(n830), .ZN(n638) );
  AOI221D1 U29 ( .A1(n806), .A2(n539), .B1(n843), .B2(n538), .C(n537), .ZN(
        n540) );
  AOI221XD4 U30 ( .A1(n845), .A2(n440), .B1(n855), .B2(n442), .C(n642), .ZN(
        n643) );
  INVD4 U31 ( .I(n444), .ZN(n443) );
  AN2D1 U32 ( .A1(n438), .A2(n444), .Z(n427) );
  ND2D2 U33 ( .A1(n440), .A2(n444), .ZN(n746) );
  CKND2 U34 ( .I(a[1]), .ZN(n444) );
  CKBD4 U36 ( .I(a[5]), .Z(n434) );
  ND2D3 U37 ( .A1(n442), .A2(n440), .ZN(n740) );
  CKND2 U38 ( .I(n444), .ZN(n442) );
  INVD4 U39 ( .I(n437), .ZN(n440) );
  OAI32D2 U40 ( .A1(n586), .A2(n746), .A3(n687), .B1(n585), .B2(n767), .ZN(
        n587) );
  NR2XD1 U41 ( .A1(n831), .A2(n827), .ZN(n675) );
  INVD2 U42 ( .I(n748), .ZN(n827) );
  AOI21D2 U43 ( .A1(n813), .A2(n442), .B(n804), .ZN(n585) );
  OAI222D1 U44 ( .A1(n732), .A2(n721), .B1(n699), .B2(n440), .C1(n698), .C2(
        n775), .ZN(n700) );
  NR2D0 U45 ( .A1(n753), .A2(n771), .ZN(n694) );
  CKND2D2 U46 ( .A1(n832), .A2(n837), .ZN(n753) );
  INVD4 U47 ( .I(n434), .ZN(n825) );
  CKND2D1 U48 ( .A1(a[3]), .A2(n445), .ZN(n679) );
  BUFFD4 U49 ( .I(n799), .Z(n436) );
  INVD1 U50 ( .I(n613), .ZN(n828) );
  INVD1 U51 ( .I(n753), .ZN(n843) );
  NR4D0 U52 ( .A1(n534), .A2(n533), .A3(n532), .A4(n596), .ZN(n535) );
  AOI22D1 U53 ( .A1(n828), .A2(n48), .B1(n806), .B2(n825), .ZN(n560) );
  INVD2 U54 ( .I(n754), .ZN(n801) );
  ND2D1 U55 ( .A1(a[3]), .A2(n817), .ZN(n751) );
  INVD2 U56 ( .I(n787), .ZN(n803) );
  INVD1 U57 ( .I(n48), .ZN(n226) );
  INVD1 U58 ( .I(n749), .ZN(n808) );
  ND2D2 U59 ( .A1(n435), .A2(a[6]), .ZN(n706) );
  ND3D2 U60 ( .A1(n51), .A2(n53), .A3(n844), .ZN(n670) );
  OR2D1 U61 ( .A1(n667), .A2(n666), .Z(n53) );
  ND2D1 U62 ( .A1(a[3]), .A2(n825), .ZN(n748) );
  ND2D1 U63 ( .A1(a[6]), .A2(n837), .ZN(n782) );
  NR2D1 U64 ( .A1(n800), .A2(n427), .ZN(n691) );
  ND2D1 U65 ( .A1(n436), .A2(n446), .ZN(n686) );
  INVD1 U66 ( .I(n657), .ZN(n834) );
  INVD2 U67 ( .I(n439), .ZN(n438) );
  ND2D2 U68 ( .A1(n438), .A2(n432), .ZN(n762) );
  INVD1 U69 ( .I(n686), .ZN(n813) );
  ND2D1 U70 ( .A1(n433), .A2(n446), .ZN(n711) );
  OAI222D0 U71 ( .A1(n465), .A2(n751), .B1(n687), .B2(n516), .C1(n464), .C2(
        n440), .ZN(n466) );
  OAI222D1 U72 ( .A1(n570), .A2(n711), .B1(n569), .B2(n745), .C1(n442), .C2(
        n568), .ZN(n571) );
  AOI21D1 U73 ( .A1(n859), .A2(n48), .B(n853), .ZN(n568) );
  INVD1 U74 ( .I(a[3]), .ZN(n446) );
  AN2XD1 U75 ( .A1(a[3]), .A2(n432), .Z(n48) );
  ND2D1 U76 ( .A1(n435), .A2(n825), .ZN(n729) );
  OAI33D0 U77 ( .A1(n657), .A2(n438), .A3(n436), .B1(n486), .B2(n729), .B3(
        n762), .ZN(n487) );
  NR2XD0 U78 ( .A1(n830), .A2(n310), .ZN(n517) );
  OAI31D0 U79 ( .A1(n801), .A2(n427), .A3(n310), .B(n858), .ZN(n491) );
  AOI31D0 U80 ( .A1(n433), .A2(n832), .A3(n310), .B(n696), .ZN(n474) );
  CKND2D1 U81 ( .A1(n825), .A2(n832), .ZN(n657) );
  INVD2 U82 ( .I(n726), .ZN(n800) );
  ND2D3 U83 ( .A1(n438), .A2(n436), .ZN(n726) );
  INVD1 U84 ( .I(n559), .ZN(n802) );
  ND2D2 U85 ( .A1(n828), .A2(n846), .ZN(n732) );
  OAI221D1 U86 ( .A1(n617), .A2(n767), .B1(n752), .B2(n762), .C(n496), .ZN(
        n499) );
  AN2XD1 U87 ( .A1(n814), .A2(n603), .Z(n72) );
  CKND2D0 U89 ( .A1(n828), .A2(n857), .ZN(n678) );
  AOI211XD0 U90 ( .A1(n857), .A2(n495), .B(n494), .C(n493), .ZN(n509) );
  OAI221D1 U91 ( .A1(n686), .A2(n676), .B1(n675), .B2(n787), .C(n674), .ZN(
        n677) );
  AOI221D1 U92 ( .A1(n859), .A2(n444), .B1(n841), .B2(n720), .C(n528), .ZN(
        n531) );
  INVD2 U93 ( .I(n770), .ZN(n831) );
  OA222D1 U94 ( .A1(n666), .A2(n770), .B1(n437), .B2(n560), .C1(n752), .C2(
        n559), .Z(n429) );
  AOI221D1 U95 ( .A1(n798), .A2(n689), .B1(n831), .B2(n800), .C(n688), .ZN(
        n690) );
  OAI222D1 U96 ( .A1(n785), .A2(n584), .B1(n777), .B2(n639), .C1(n497), .C2(
        n765), .ZN(n498) );
  CKND2D1 U97 ( .A1(n843), .A2(n830), .ZN(n785) );
  ND2D1 U98 ( .A1(n827), .A2(n846), .ZN(n599) );
  NR2XD0 U99 ( .A1(n817), .A2(n825), .ZN(n672) );
  ND2D0 U100 ( .A1(n438), .A2(n444), .ZN(n745) );
  AOI221D1 U101 ( .A1(n843), .A2(n459), .B1(n458), .B2(n440), .C(n457), .ZN(
        n482) );
  NR2D0 U102 ( .A1(n708), .A2(n711), .ZN(n719) );
  OAI22D1 U103 ( .A1(n470), .A2(n711), .B1(n469), .B2(n762), .ZN(n471) );
  AOI222D1 U104 ( .A1(n808), .A2(n828), .B1(n806), .B2(n485), .C1(n802), .C2(
        n831), .ZN(n490) );
  AOI221D1 U105 ( .A1(n820), .A2(n857), .B1(n310), .B2(n830), .C(n529), .ZN(
        n530) );
  AOI221D1 U106 ( .A1(n463), .A2(n808), .B1(n850), .B2(n815), .C(n462), .ZN(
        n464) );
  ND2D0 U107 ( .A1(n434), .A2(n446), .ZN(n770) );
  AOI221D1 U108 ( .A1(n427), .A2(n684), .B1(n683), .B2(n806), .C(n682), .ZN(
        n685) );
  AOI22D1 U109 ( .A1(n836), .A2(n806), .B1(n809), .B2(n835), .ZN(n470) );
  INVD2 U110 ( .I(n666), .ZN(n806) );
  CKND2D1 U111 ( .A1(a[3]), .A2(n434), .ZN(n687) );
  OAI21D0 U112 ( .A1(n437), .A2(n687), .B(n751), .ZN(n485) );
  INVD0 U113 ( .I(n687), .ZN(n829) );
  CKND2D1 U114 ( .A1(a[6]), .A2(n825), .ZN(n775) );
  INVD4 U115 ( .I(n435), .ZN(n837) );
  ND4D2 U116 ( .A1(n718), .A2(n717), .A3(n716), .A4(n715), .ZN(d[1]) );
  OAI222D1 U117 ( .A1(n226), .A2(n637), .B1(n592), .B2(n591), .C1(n590), .C2(
        n759), .ZN(n593) );
  ND2D1 U118 ( .A1(n672), .A2(n857), .ZN(n776) );
  CKND2D1 U119 ( .A1(n447), .A2(n817), .ZN(n757) );
  NR2D0 U120 ( .A1(n757), .A2(n556), .ZN(n426) );
  AOI221D1 U121 ( .A1(n833), .A2(n796), .B1(n594), .B2(n444), .C(n736), .ZN(
        n595) );
  INVD2 U122 ( .I(n638), .ZN(n852) );
  NR2D0 U123 ( .A1(n638), .A2(n723), .ZN(n742) );
  AOI21D1 U124 ( .A1(n831), .A2(n840), .B(n849), .ZN(n667) );
  OAI221D1 U125 ( .A1(n612), .A2(n586), .B1(a[3]), .B2(n776), .C(n703), .ZN(
        n529) );
  CKND2D1 U126 ( .A1(n828), .A2(n840), .ZN(n724) );
  CKND0 U127 ( .I(n729), .ZN(n856) );
  OA221D1 U128 ( .A1(n751), .A2(n428), .B1(n687), .B2(n749), .C(n429), .Z(n561) );
  ND2D1 U129 ( .A1(n443), .A2(n432), .ZN(n749) );
  OAI222D1 U130 ( .A1(n747), .A2(n720), .B1(n771), .B2(n584), .C1(n752), .C2(
        n762), .ZN(n588) );
  CKND2D1 U131 ( .A1(n817), .A2(n825), .ZN(n771) );
  OAI221D1 U132 ( .A1(n740), .A2(n686), .B1(n748), .B2(n705), .C(n685), .ZN(
        n693) );
  OA21D0 U133 ( .A1(n686), .A2(n441), .B(n616), .Z(n620) );
  ND2D1 U134 ( .A1(n443), .A2(n437), .ZN(n720) );
  AOI211XD0 U135 ( .A1(n804), .A2(n821), .B(n824), .C(n697), .ZN(n698) );
  NR4D1 U136 ( .A1(n789), .A2(n790), .A3(n791), .A4(n788), .ZN(n792) );
  OAI222D1 U137 ( .A1(n783), .A2(n782), .B1(a[3]), .B2(n838), .C1(n781), .C2(
        n440), .ZN(n789) );
  AOI22D1 U138 ( .A1(n440), .A2(n815), .B1(n447), .B2(n805), .ZN(n592) );
  AOI211XD0 U139 ( .A1(n861), .A2(n809), .B(n483), .C(n665), .ZN(n510) );
  OA221D1 U140 ( .A1(n633), .A2(n762), .B1(n430), .B2(n787), .C(n431), .Z(n718) );
  BUFFD4 U141 ( .I(a[7]), .Z(n435) );
  ND2D4 U142 ( .A1(n443), .A2(n436), .ZN(n787) );
  ND2D2 U143 ( .A1(n445), .A2(n436), .ZN(n754) );
  NR4D1 U144 ( .A1(n543), .A2(n544), .A3(n542), .A4(n541), .ZN(n545) );
  OAI33D0 U145 ( .A1(n757), .A2(n436), .A3(n729), .B1(n657), .B2(n442), .B3(
        n656), .ZN(n660) );
  CKND1 U146 ( .I(n785), .ZN(n845) );
  CKND2D0 U147 ( .A1(n726), .A2(n754), .ZN(n526) );
  AOI221D1 U148 ( .A1(n801), .A2(n822), .B1(n809), .B2(n829), .C(n768), .ZN(
        n783) );
  AOI221D1 U149 ( .A1(n702), .A2(n856), .B1(n48), .B2(n701), .C(n700), .ZN(
        n716) );
  OAI222D1 U150 ( .A1(n563), .A2(n759), .B1(n686), .B2(n562), .C1(n561), .C2(
        n753), .ZN(n564) );
  INVD6 U151 ( .I(n433), .ZN(n817) );
  AOI221D1 U152 ( .A1(n834), .A2(n822), .B1(n820), .B2(n573), .C(n849), .ZN(
        n497) );
  AOI221D1 U153 ( .A1(n840), .A2(n499), .B1(n802), .B2(n512), .C(n498), .ZN(
        n508) );
  AOI221D1 U154 ( .A1(n858), .A2(n440), .B1(n850), .B2(n808), .C(n634), .ZN(
        n664) );
  AOI221D1 U155 ( .A1(n802), .A2(n848), .B1(n796), .B2(n861), .C(n593), .ZN(
        n626) );
  AOI221D1 U156 ( .A1(n854), .A2(n796), .B1(n857), .B2(n693), .C(n692), .ZN(
        n717) );
  OR2XD1 U157 ( .A1(n668), .A2(n679), .Z(n51) );
  NR2XD1 U158 ( .A1(n841), .A2(n852), .ZN(n668) );
  ND2D2 U159 ( .A1(n432), .A2(n445), .ZN(n666) );
  INR4D2 U160 ( .A1(n671), .B1(n670), .B2(n669), .B3(n853), .ZN(n681) );
  CKAN2D1 U161 ( .A1(n442), .A2(n467), .Z(n68) );
  CKAN2D1 U162 ( .A1(n824), .A2(n834), .Z(n70) );
  NR3D0 U163 ( .A1(n68), .A2(n70), .A3(n466), .ZN(n481) );
  CKAN2D1 U164 ( .A1(n840), .A2(n602), .Z(n187) );
  NR3D1 U165 ( .A1(n72), .A2(n187), .A3(n601), .ZN(n625) );
  AOI221D1 U166 ( .A1(n812), .A2(n573), .B1(n572), .B2(n820), .C(n571), .ZN(
        n581) );
  AOI221D1 U167 ( .A1(n827), .A2(n798), .B1(n819), .B2(n806), .C(n677), .ZN(
        n680) );
  AOI221D1 U168 ( .A1(n437), .A2(n566), .B1(n840), .B2(n565), .C(n564), .ZN(
        n582) );
  OAI211D0 U169 ( .A1(n825), .A2(n757), .B(n774), .C(n752), .ZN(n684) );
  BUFFD8 U170 ( .I(a[2]), .Z(n432) );
  CKAN2D1 U171 ( .A1(a[3]), .A2(n436), .Z(n310) );
  NR2D0 U172 ( .A1(n726), .A2(n751), .ZN(n424) );
  NR2D0 U173 ( .A1(n691), .A2(n687), .ZN(n425) );
  OR3D1 U174 ( .A1(n424), .A2(n425), .A3(n426), .Z(n534) );
  ND2D0 U175 ( .A1(n432), .A2(n446), .ZN(n777) );
  AOI21D1 U176 ( .A1(n818), .A2(n860), .B(n847), .ZN(n569) );
  INR2D0 U177 ( .A1(n763), .B1(n501), .ZN(n502) );
  CKND2D0 U178 ( .A1(n432), .A2(n740), .ZN(n738) );
  CKND2D0 U179 ( .A1(n860), .A2(n822), .ZN(n786) );
  CKND2D0 U180 ( .A1(n784), .A2(n686), .ZN(n525) );
  CKND2D0 U181 ( .A1(n833), .A2(n822), .ZN(n536) );
  NR2D0 U182 ( .A1(n808), .A2(n796), .ZN(n616) );
  CKND0 U183 ( .I(n722), .ZN(n842) );
  NR2XD0 U184 ( .A1(n835), .A2(n846), .ZN(n641) );
  OAI22D1 U185 ( .A1(n746), .A2(n708), .B1(n641), .B2(n740), .ZN(n642) );
  CKND2D0 U186 ( .A1(n765), .A2(n762), .ZN(n750) );
  CKND2D0 U187 ( .A1(n672), .A2(n846), .ZN(n591) );
  CKND0 U188 ( .I(n704), .ZN(n860) );
  NR2XD0 U189 ( .A1(n858), .A2(n512), .ZN(n513) );
  ND2D0 U190 ( .A1(n432), .A2(n817), .ZN(n628) );
  ND2D0 U191 ( .A1(n434), .A2(n837), .ZN(n708) );
  CKND2D0 U192 ( .A1(n442), .A2(a[6]), .ZN(n486) );
  AOI22D0 U193 ( .A1(n859), .A2(n803), .B1(n815), .B2(n845), .ZN(n550) );
  NR2D0 U194 ( .A1(n441), .A2(n761), .ZN(n743) );
  NR2D0 U195 ( .A1(n805), .A2(n801), .ZN(n475) );
  NR2D0 U196 ( .A1(n800), .A2(n797), .ZN(n617) );
  ND2D0 U197 ( .A1(n310), .A2(n852), .ZN(n567) );
  NR2D0 U198 ( .A1(n719), .A2(n855), .ZN(n727) );
  CKND2D0 U200 ( .A1(n784), .A2(n556), .ZN(n557) );
  NR2D0 U201 ( .A1(n732), .A2(a[3]), .ZN(n696) );
  OAI22D0 U202 ( .A1(n745), .A2(n757), .B1(n604), .B2(n746), .ZN(n611) );
  NR2D0 U203 ( .A1(n823), .A2(n828), .ZN(n604) );
  AOI22D0 U204 ( .A1(n808), .A2(n437), .B1(n442), .B2(n48), .ZN(n484) );
  CKND0 U205 ( .I(n746), .ZN(n797) );
  CKND2D0 U206 ( .A1(n808), .A2(n440), .ZN(n707) );
  CKND2D0 U207 ( .A1(n438), .A2(n806), .ZN(n730) );
  AOI31D0 U208 ( .A1(n733), .A2(n732), .A3(n731), .B(n730), .ZN(n734) );
  NR2D0 U210 ( .A1(n48), .A2(n821), .ZN(n656) );
  ND2D0 U211 ( .A1(n820), .A2(n860), .ZN(n763) );
  CKND2D0 U212 ( .A1(n819), .A2(n843), .ZN(n671) );
  NR2D0 U213 ( .A1(n810), .A2(n808), .ZN(n468) );
  ND2D0 U214 ( .A1(n798), .A2(n857), .ZN(n516) );
  CKND0 U216 ( .I(n584), .ZN(n812) );
  AOI22D0 U217 ( .A1(n809), .A2(n856), .B1(n801), .B2(n835), .ZN(n570) );
  CKND2D0 U218 ( .A1(n828), .A2(n444), .ZN(n676) );
  OAI21D0 U219 ( .A1(n753), .A2(n613), .B(n722), .ZN(n594) );
  NR2D0 U220 ( .A1(n859), .A2(n845), .ZN(n460) );
  CKND2D0 U221 ( .A1(n48), .A2(n817), .ZN(n605) );
  OAI22D0 U222 ( .A1(n440), .A2(n722), .B1(n445), .B2(n733), .ZN(n528) );
  CKND0 U223 ( .I(n639), .ZN(n851) );
  AOI211XD0 U224 ( .A1(n841), .A2(n438), .B(n640), .C(n851), .ZN(n644) );
  CKND1 U225 ( .I(n665), .ZN(n844) );
  OAI32D0 U226 ( .A1(n559), .A2(n759), .A3(n748), .B1(n517), .B2(n516), .ZN(
        n518) );
  OAI22D0 U227 ( .A1(n787), .A2(n786), .B1(n785), .B2(n784), .ZN(n788) );
  CKND2D1 U228 ( .A1(n492), .A2(n491), .ZN(n493) );
  CKND2D0 U229 ( .A1(n440), .A2(n436), .ZN(n765) );
  CKND2D0 U230 ( .A1(a[3]), .A2(n436), .ZN(n774) );
  OAI31D0 U231 ( .A1(n740), .A2(n821), .A3(n753), .B(n739), .ZN(n744) );
  AOI31D0 U232 ( .A1(n846), .A2(n738), .A3(n821), .B(n737), .ZN(n739) );
  ND2D0 U233 ( .A1(n825), .A2(n837), .ZN(n612) );
  OAI22D0 U234 ( .A1(n767), .A2(n777), .B1(n442), .B2(n766), .ZN(n768) );
  AOI22D0 U235 ( .A1(n310), .A2(n830), .B1(n813), .B2(n825), .ZN(n766) );
  AOI32D0 U236 ( .A1(n801), .A2(n440), .A3(n831), .B1(n798), .B2(n552), .ZN(
        n554) );
  NR2D0 U237 ( .A1(n628), .A2(n720), .ZN(n702) );
  OAI21D0 U238 ( .A1(n752), .A2(n612), .B(n637), .ZN(n512) );
  AOI21D0 U239 ( .A1(n613), .A2(n657), .B(n686), .ZN(n501) );
  CKND2D0 U240 ( .A1(n683), .A2(n846), .ZN(n633) );
  ND2D0 U241 ( .A1(n436), .A2(n817), .ZN(n555) );
  CKND2D0 U242 ( .A1(n826), .A2(n846), .ZN(n637) );
  CKND2D0 U243 ( .A1(n797), .A2(n446), .ZN(n723) );
  CKND2D0 U244 ( .A1(n687), .A2(n751), .ZN(n689) );
  CKND2D0 U245 ( .A1(n829), .A2(n846), .ZN(n764) );
  AOI211D0 U246 ( .A1(n816), .A2(n438), .B(n48), .C(n810), .ZN(n606) );
  NR2XD0 U247 ( .A1(n648), .A2(n769), .ZN(n607) );
  CKND2D0 U248 ( .A1(n820), .A2(n846), .ZN(n608) );
  CKND1 U249 ( .I(n797), .ZN(n428) );
  CKND0 U250 ( .I(n694), .ZN(n430) );
  CKND2D0 U251 ( .A1(n800), .A2(n830), .ZN(n647) );
  AOI21D0 U252 ( .A1(n845), .A2(n48), .B(n755), .ZN(n756) );
  OAI21D0 U253 ( .A1(n226), .A2(n732), .B(n786), .ZN(n473) );
  CKND2D1 U254 ( .A1(n598), .A2(n597), .ZN(n602) );
  AOI21D0 U255 ( .A1(n807), .A2(n843), .B(n572), .ZN(n514) );
  NR2D0 U256 ( .A1(n810), .A2(a[3]), .ZN(n619) );
  OAI211D0 U257 ( .A1(n704), .A2(n679), .B(n551), .C(n550), .ZN(n566) );
  AOI21D0 U258 ( .A1(n820), .A2(n856), .B(n696), .ZN(n504) );
  CKND0 U259 ( .I(n769), .ZN(n838) );
  CKND2D0 U260 ( .A1(n720), .A2(n446), .ZN(n575) );
  AOI21D0 U261 ( .A1(n855), .A2(n815), .B(n696), .ZN(n699) );
  ND4D0 U262 ( .A1(n427), .A2(n834), .A3(n433), .A4(n435), .ZN(n728) );
  OAI22D0 U263 ( .A1(n767), .A2(n686), .B1(n691), .B2(n711), .ZN(n454) );
  AOI21D0 U264 ( .A1(n686), .A2(n586), .B(n745), .ZN(n453) );
  AOI211D0 U265 ( .A1(n778), .A2(n657), .B(n586), .C(n745), .ZN(n476) );
  OAI31D0 U266 ( .A1(n749), .A2(n778), .A3(n751), .B(n615), .ZN(n622) );
  AOI33D0 U267 ( .A1(n614), .A2(n832), .A3(n803), .B1(n852), .B2(n446), .B3(
        n798), .ZN(n615) );
  OAI22D0 U268 ( .A1(a[3]), .A2(n613), .B1(n440), .B2(n612), .ZN(n614) );
  OAI33D0 U269 ( .A1(n226), .A2(n435), .A3(n771), .B1(n704), .B2(n436), .B3(
        n752), .ZN(n537) );
  OAI21D0 U270 ( .A1(n657), .A2(n751), .B(n731), .ZN(n539) );
  CKND0 U272 ( .I(n612), .ZN(n839) );
  AOI21D0 U273 ( .A1(a[3]), .A2(n857), .B(n816), .ZN(n772) );
  OAI22D0 U274 ( .A1(n832), .A2(n711), .B1(n817), .B2(n657), .ZN(n649) );
  OAI22D0 U275 ( .A1(n435), .A2(n657), .B1(n752), .B2(n729), .ZN(n450) );
  NR2D0 U276 ( .A1(n855), .A2(n694), .ZN(n452) );
  OAI32D0 U277 ( .A1(n770), .A2(n475), .A3(n706), .B1(n474), .B2(n740), .ZN(
        n478) );
  CKND2D0 U278 ( .A1(n433), .A2(n436), .ZN(n586) );
  AOI21D0 U279 ( .A1(n854), .A2(n442), .B(n694), .ZN(n695) );
  CKND2D1 U280 ( .A1(n775), .A2(n729), .ZN(n573) );
  OAI21D0 U281 ( .A1(n710), .A2(n740), .B(n709), .ZN(n714) );
  OA33D0 U282 ( .A1(n708), .A2(n752), .A3(n745), .B1(n707), .B2(n706), .B3(
        n770), .Z(n709) );
  CKND2D0 U283 ( .A1(n434), .A2(a[6]), .ZN(n778) );
  AOI32D0 U284 ( .A1(n433), .A2(n837), .A3(n814), .B1(n48), .B2(n549), .ZN(
        n551) );
  CKND1 U285 ( .I(a[6]), .ZN(n832) );
  INVD1 U287 ( .I(n556), .ZN(n804) );
  INVD1 U288 ( .I(n567), .ZN(n853) );
  INVD1 U289 ( .I(n720), .ZN(n796) );
  INVD1 U290 ( .I(n784), .ZN(n815) );
  INVD1 U291 ( .I(n678), .ZN(n859) );
  INVD1 U292 ( .I(n740), .ZN(n798) );
  ND2D1 U293 ( .A1(n803), .A2(n440), .ZN(n556) );
  INVD1 U294 ( .I(n707), .ZN(n809) );
  ND2D1 U295 ( .A1(n730), .A2(n740), .ZN(n589) );
  INVD1 U296 ( .I(n730), .ZN(n807) );
  INVD1 U298 ( .I(n786), .ZN(n861) );
  INVD1 U299 ( .I(n600), .ZN(n824) );
  AOI222D0 U300 ( .A1(n808), .A2(n822), .B1(n820), .B2(n800), .C1(n829), .C2(
        n806), .ZN(n553) );
  ND2D1 U301 ( .A1(n442), .A2(a[3]), .ZN(n784) );
  NR2D1 U302 ( .A1(n761), .A2(n438), .ZN(n713) );
  INVD1 U303 ( .I(n591), .ZN(n855) );
  NR2D1 U304 ( .A1(n627), .A2(n745), .ZN(n769) );
  INVD1 U305 ( .I(n765), .ZN(n805) );
  INVD1 U306 ( .I(n757), .ZN(n819) );
  INVD1 U307 ( .I(n599), .ZN(n849) );
  INVD1 U308 ( .I(n637), .ZN(n854) );
  INVD1 U309 ( .I(n732), .ZN(n850) );
  INVD1 U310 ( .I(n679), .ZN(n816) );
  INVD1 U311 ( .I(n771), .ZN(n826) );
  INVD1 U312 ( .I(n724), .ZN(n841) );
  ND2D1 U313 ( .A1(n814), .A2(n442), .ZN(n721) );
  AO221D0 U314 ( .A1(n801), .A2(n831), .B1(n798), .B2(n814), .C(n702), .Z(n654) );
  ND2D1 U315 ( .A1(n796), .A2(n823), .ZN(n600) );
  ND2D1 U316 ( .A1(n801), .A2(n437), .ZN(n559) );
  INVD1 U317 ( .I(n608), .ZN(n847) );
  ND2D1 U318 ( .A1(n818), .A2(n834), .ZN(n703) );
  AOI221D0 U319 ( .A1(n804), .A2(n831), .B1(n826), .B2(n557), .C(n702), .ZN(
        n563) );
  INVD1 U320 ( .I(n555), .ZN(n818) );
  OAI222D0 U321 ( .A1(n727), .A2(n726), .B1(n725), .B2(n724), .C1(n723), .C2(
        n722), .ZN(n795) );
  OAI222D0 U322 ( .A1(n754), .A2(n687), .B1(n484), .B2(n767), .C1(n442), .C2(
        n752), .ZN(n495) );
  OAI222D0 U323 ( .A1(n748), .A2(n556), .B1(n226), .B2(n720), .C1(n749), .C2(
        n687), .ZN(n455) );
  NR4D0 U324 ( .A1(n711), .A2(n765), .A3(n759), .A4(n825), .ZN(n737) );
  OAI221D0 U325 ( .A1(n460), .A2(n777), .B1(n722), .B2(n774), .C(n567), .ZN(
        n467) );
  OAI222D0 U326 ( .A1(n759), .A2(n628), .B1(a[3]), .B2(n627), .C1(n753), .C2(
        n770), .ZN(n631) );
  OAI222D0 U327 ( .A1(n765), .A2(n764), .B1(n763), .B2(n762), .C1(n442), .C2(
        n761), .ZN(n790) );
  OAI222D0 U328 ( .A1(n760), .A2(n759), .B1(n758), .B2(n757), .C1(n438), .C2(
        n756), .ZN(n791) );
  OAI222D0 U329 ( .A1(n762), .A2(n770), .B1(n784), .B2(n647), .C1(n751), .C2(
        n707), .ZN(n655) );
  OAI221D0 U330 ( .A1(n449), .A2(n613), .B1(n777), .B2(n720), .C(n448), .ZN(
        n459) );
  AOI221D0 U331 ( .A1(n801), .A2(n856), .B1(n810), .B2(n835), .C(n461), .ZN(
        n465) );
  ND2D1 U332 ( .A1(n840), .A2(n826), .ZN(n722) );
  ND2D1 U333 ( .A1(n752), .A2(n747), .ZN(n552) );
  NR3D0 U334 ( .A1(n720), .A2(n817), .A3(n731), .ZN(n577) );
  NR3D0 U335 ( .A1(n740), .A2(a[3]), .A3(n767), .ZN(n533) );
  INVD1 U336 ( .I(n767), .ZN(n830) );
  ND2D1 U337 ( .A1(n683), .A2(n843), .ZN(n731) );
  NR3D0 U338 ( .A1(n511), .A2(n752), .A3(n787), .ZN(n477) );
  INVD1 U339 ( .I(n711), .ZN(n822) );
  INVD1 U340 ( .I(n777), .ZN(n814) );
  INVD1 U341 ( .I(n752), .ZN(n821) );
  NR2D1 U342 ( .A1(n704), .A2(n746), .ZN(n736) );
  INVD1 U343 ( .I(n705), .ZN(n823) );
  OAI222D0 U344 ( .A1(n638), .A2(n436), .B1(n612), .B2(n605), .C1(a[3]), .C2(
        n722), .ZN(n610) );
  AOI221D0 U345 ( .A1(n796), .A2(n813), .B1(n802), .B2(n827), .C(n596), .ZN(
        n597) );
  INVD1 U346 ( .I(n759), .ZN(n857) );
  INVD1 U347 ( .I(n511), .ZN(n833) );
  INVD1 U348 ( .I(n738), .ZN(n811) );
  NR4D0 U349 ( .A1(n455), .A2(n454), .A3(n532), .A4(n453), .ZN(n456) );
  AOI222D0 U350 ( .A1(n803), .A2(n819), .B1(n821), .B2(n805), .C1(n807), .C2(
        n434), .ZN(n598) );
  OAI222D0 U351 ( .A1(n729), .A2(n600), .B1(n726), .B2(n764), .C1(n616), .C2(
        n599), .ZN(n601) );
  OAI221D0 U352 ( .A1(n740), .A2(n733), .B1(n706), .B2(n746), .C(n595), .ZN(
        n603) );
  NR4D0 U353 ( .A1(n631), .A2(n630), .A3(n847), .A4(n629), .ZN(n632) );
  OAI221D0 U354 ( .A1(n452), .A2(n226), .B1(n774), .B2(n733), .C(n451), .ZN(
        n458) );
  NR4D0 U355 ( .A1(n443), .A2(n837), .A3(n765), .A4(n757), .ZN(n697) );
  OAI222D0 U356 ( .A1(n435), .A2(n773), .B1(n772), .B2(n771), .C1(n782), .C2(
        n770), .ZN(n780) );
  OAI222D0 U357 ( .A1(n432), .A2(n652), .B1(n651), .B2(n786), .C1(n650), .C2(
        n785), .ZN(n653) );
  AOI21D1 U358 ( .A1(n796), .A2(n649), .B(n648), .ZN(n652) );
  NR3D0 U359 ( .A1(n673), .A2(n801), .A3(n814), .ZN(n650) );
  NR2XD0 U360 ( .A1(n780), .A2(n779), .ZN(n781) );
  OAI222D0 U361 ( .A1(n515), .A2(n745), .B1(n514), .B2(n752), .C1(n513), .C2(
        n765), .ZN(n519) );
  NR2D1 U362 ( .A1(n433), .A2(n832), .ZN(n463) );
  OAI211D1 U363 ( .A1(n555), .A2(n720), .B(n554), .C(n553), .ZN(n565) );
  OAI222D0 U364 ( .A1(n576), .A2(n776), .B1(n785), .B2(n575), .C1(n574), .C2(
        n778), .ZN(n579) );
  OAI221D0 U365 ( .A1(n752), .A2(n754), .B1(n711), .B2(n787), .C(n636), .ZN(
        n646) );
  OAI221D0 U366 ( .A1(n442), .A2(n671), .B1(n723), .B2(n678), .C(n527), .ZN(
        n544) );
  OAI222D0 U367 ( .A1(n707), .A2(n733), .B1(n437), .B2(n540), .C1(n787), .C2(
        n776), .ZN(n541) );
  AOI221D0 U368 ( .A1(n473), .A2(n444), .B1(n819), .B2(n472), .C(n471), .ZN(
        n480) );
  OAI222D0 U369 ( .A1(n475), .A2(n708), .B1(n468), .B2(n706), .C1(n729), .C2(
        n730), .ZN(n472) );
  NR3D0 U370 ( .A1(n740), .A2(n433), .A3(n612), .ZN(n648) );
  ND2D1 U371 ( .A1(n433), .A2(n825), .ZN(n613) );
  NR4D0 U372 ( .A1(n438), .A2(n832), .A3(n771), .A4(n777), .ZN(n578) );
  NR3D0 U373 ( .A1(n777), .A2(n435), .A3(n433), .ZN(n669) );
  OAI221D0 U374 ( .A1(n740), .A2(n729), .B1(n443), .B2(n785), .C(n728), .ZN(
        n735) );
  NR3D0 U375 ( .A1(n441), .A2(n433), .A3(n687), .ZN(n596) );
  OAI222D0 U376 ( .A1(n442), .A2(n778), .B1(n746), .B2(n759), .C1(n753), .C2(
        n749), .ZN(n488) );
  NR3D0 U377 ( .A1(n706), .A2(n825), .A3(n711), .ZN(n523) );
  ND2D1 U378 ( .A1(n435), .A2(n832), .ZN(n759) );
  NR3D0 U379 ( .A1(n721), .A2(n433), .A3(n837), .ZN(n659) );
  ND2D1 U380 ( .A1(n434), .A2(n435), .ZN(n704) );
  INVD1 U381 ( .I(n775), .ZN(n835) );
  INVD1 U382 ( .I(n706), .ZN(n846) );
  ND2D1 U383 ( .A1(n434), .A2(n832), .ZN(n511) );
  ND2D1 U384 ( .A1(n433), .A2(n432), .ZN(n705) );
  OAI222D0 U385 ( .A1(n504), .A2(n746), .B1(n817), .B2(n503), .C1(n502), .C2(
        n720), .ZN(n506) );
  ND2D1 U386 ( .A1(n435), .A2(n500), .ZN(n503) );
  INVD1 U387 ( .I(n778), .ZN(n836) );
  OAI222D0 U388 ( .A1(n620), .A2(n776), .B1(n619), .B2(n724), .C1(n618), .C2(
        n757), .ZN(n621) );
  OA22D0 U389 ( .A1(n778), .A2(n745), .B1(n729), .B2(n617), .Z(n618) );
  INVD1 U390 ( .I(n432), .ZN(n799) );
  INVD1 U391 ( .I(a[1]), .ZN(n445) );
  INVD1 U392 ( .I(a[3]), .ZN(n447) );
  NR4D0 U393 ( .A1(a[6]), .A2(n447), .A3(n729), .A4(n762), .ZN(n505) );
  ND3D1 U394 ( .A1(n545), .A2(n546), .A3(n547), .ZN(d[5]) );
  INR4D0 U395 ( .A1(n761), .B1(n524), .B2(n742), .B3(n712), .ZN(n546) );
  ND4D1 U396 ( .A1(n626), .A2(n625), .A3(n624), .A4(n623), .ZN(d[3]) );
  NR2D1 U397 ( .A1(n622), .A2(n621), .ZN(n623) );
  AOI221D0 U398 ( .A1(n843), .A2(n611), .B1(n610), .B2(n440), .C(n609), .ZN(
        n624) );
  AOI221D0 U399 ( .A1(n736), .A2(n814), .B1(n813), .B2(n735), .C(n734), .ZN(
        n794) );
  NR4D0 U400 ( .A1(n744), .A2(n743), .A3(n742), .A4(n741), .ZN(n793) );
  ND4D1 U401 ( .A1(n664), .A2(n663), .A3(n662), .A4(n661), .ZN(d[2]) );
  NR4D0 U402 ( .A1(n660), .A2(n659), .A3(n658), .A4(n743), .ZN(n661) );
  ND4D1 U403 ( .A1(n480), .A2(n481), .A3(n482), .A4(n479), .ZN(d[7]) );
  NR4D0 U404 ( .A1(n478), .A2(n477), .A3(n713), .A4(n476), .ZN(n479) );
  ND4D1 U405 ( .A1(n510), .A2(n509), .A3(n508), .A4(n507), .ZN(d[6]) );
  NR4D0 U406 ( .A1(n506), .A2(n505), .A3(n521), .A4(n522), .ZN(n507) );
  NR4D0 U407 ( .A1(n579), .A2(n578), .A3(n577), .A4(n741), .ZN(n580) );
  NR4D0 U408 ( .A1(n714), .A2(n737), .A3(n713), .A4(n712), .ZN(n715) );
  NR2D1 U409 ( .A1(n804), .A2(n807), .ZN(n576) );
  OAI31D0 U410 ( .A1(n446), .A2(n804), .A3(n810), .B(n694), .ZN(n492) );
  AOI221D0 U411 ( .A1(n310), .A2(n842), .B1(n850), .B2(n815), .C(n548), .ZN(
        n583) );
  NR2D1 U412 ( .A1(n310), .A2(n805), .ZN(n449) );
  OAI22D1 U413 ( .A1(n226), .A2(n745), .B1(n746), .B2(n774), .ZN(n500) );
  OAI222D0 U414 ( .A1(n778), .A2(n787), .B1(n777), .B2(n776), .C1(n775), .C2(
        n774), .ZN(n779) );
  AOI22D0 U415 ( .A1(n803), .A2(n834), .B1(n310), .B2(n817), .ZN(n773) );
  OAI22D0 U416 ( .A1(n757), .A2(n754), .B1(n656), .B2(n740), .ZN(n520) );
  OAI222D0 U417 ( .A1(n754), .A2(n608), .B1(n607), .B2(n436), .C1(n606), .C2(
        n678), .ZN(n609) );
  OAI33D0 U418 ( .A1(n754), .A2(n753), .A3(n752), .B1(n775), .B2(n436), .B3(
        n751), .ZN(n755) );
  OAI22D1 U419 ( .A1(n724), .A2(n754), .B1(n436), .B2(n731), .ZN(n665) );
  INR2XD0 U420 ( .A1(n523), .B1(n666), .ZN(n712) );
  NR2XD0 U421 ( .A1(n511), .A2(n666), .ZN(n572) );
  OAI222D0 U422 ( .A1(n226), .A2(n724), .B1(n592), .B2(n733), .C1(n638), .C2(
        n666), .ZN(n483) );
  IND4D1 U423 ( .A1(n795), .B1(n794), .B2(n793), .B3(n792), .ZN(d[0]) );
  INVD1 U424 ( .I(n776), .ZN(n858) );
  AN4D1 U425 ( .A1(n672), .A2(n815), .A3(n438), .A4(n843), .Z(n521) );
  ND3D1 U426 ( .A1(n48), .A2(n672), .A3(n843), .ZN(n761) );
  OAI222D0 U427 ( .A1(n754), .A2(n763), .B1(n691), .B2(n722), .C1(n690), .C2(
        n782), .ZN(n692) );
  OAI222D0 U428 ( .A1(n726), .A2(n599), .B1(n733), .B2(n679), .C1(n638), .C2(
        n762), .ZN(n548) );
  OAI22D0 U429 ( .A1(n445), .A2(n722), .B1(n442), .B2(n638), .ZN(n640) );
  OA222D0 U430 ( .A1(n749), .A2(n748), .B1(n747), .B2(n746), .C1(n751), .C2(
        n745), .Z(n760) );
  OAI22D0 U431 ( .A1(n748), .A2(n754), .B1(n767), .B2(n787), .ZN(n688) );
  AOI22D0 U432 ( .A1(n823), .A2(n797), .B1(n821), .B2(n432), .ZN(n574) );
  AOI31D0 U433 ( .A1(n432), .A2(n825), .A3(n427), .B(n824), .ZN(n496) );
  AOI21D0 U434 ( .A1(n732), .A2(n671), .B(n432), .ZN(n630) );
  ND2D1 U435 ( .A1(n432), .A2(n434), .ZN(n747) );
  AOI22D0 U436 ( .A1(n850), .A2(n526), .B1(n694), .B2(n525), .ZN(n527) );
  AOI32D1 U437 ( .A1(n434), .A2(n440), .A3(n815), .B1(n826), .B2(n635), .ZN(
        n636) );
  OAI22D0 U438 ( .A1(a[6]), .A2(n433), .B1(n434), .B2(n759), .ZN(n549) );
  OAI211D0 U439 ( .A1(n434), .A2(n784), .B(n628), .C(n751), .ZN(n538) );
  NR2D1 U440 ( .A1(a[3]), .A2(n434), .ZN(n683) );
  NR3D0 U441 ( .A1(n825), .A2(n443), .A3(n726), .ZN(n532) );
  AOI21D0 U442 ( .A1(n687), .A2(n767), .B(n726), .ZN(n682) );
  NR4D0 U443 ( .A1(n771), .A2(n759), .A3(n666), .A4(a[3]), .ZN(n741) );
  AOI22D0 U444 ( .A1(n827), .A2(n806), .B1(n803), .B2(n829), .ZN(n448) );
  AOI22D0 U445 ( .A1(n834), .A2(n750), .B1(n836), .B2(n806), .ZN(n758) );
  AOI32D1 U446 ( .A1(n435), .A2(n817), .A3(n801), .B1(n806), .B2(n450), .ZN(
        n451) );
  NR2D1 U447 ( .A1(n797), .A2(n806), .ZN(n651) );
  INVD1 U448 ( .I(n751), .ZN(n820) );
  OA222D1 U449 ( .A1(n437), .A2(n681), .B1(n753), .B2(n680), .C1(n679), .C2(
        n678), .Z(n431) );
  INVD1 U450 ( .I(n633), .ZN(n848) );
  INVD1 U451 ( .I(n762), .ZN(n810) );
  ND4D1 U452 ( .A1(n582), .A2(n583), .A3(n581), .A4(n580), .ZN(d[4]) );
  OAI22D0 U453 ( .A1(n456), .A2(n782), .B1(n749), .B2(n637), .ZN(n457) );
  AOI21D0 U454 ( .A1(n777), .A2(n747), .B(n782), .ZN(n629) );
  NR4D0 U455 ( .A1(n687), .A2(n754), .A3(n782), .A4(n817), .ZN(n658) );
endmodule


module aes_sbox_2 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n51, n65, n70, n72, n142, n192, n277, n304, n305, n306, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852;

  AN2XD1 U28 ( .A1(n711), .A2(n710), .Z(n715) );
  OA21D1 U35 ( .A1(n695), .A2(n694), .B(n693), .Z(n700) );
  OR3D1 U88 ( .A1(n663), .A2(n801), .A3(n436), .Z(n624) );
  OR4D1 U199 ( .A1(n648), .A2(n567), .A3(n514), .A4(n513), .Z(n516) );
  MAOI22D1 U209 ( .A1(n846), .A2(n439), .B1(n617), .B2(n764), .ZN(n507) );
  AN2XD1 U215 ( .A1(n515), .A2(n799), .Z(n514) );
  AN4XD1 U217 ( .A1(n662), .A2(n806), .A3(n431), .A4(n834), .Z(n513) );
  AO31D1 U286 ( .A1(n792), .A2(n848), .A3(n673), .B(n709), .Z(n454) );
  OAI222D0 U1 ( .A1(n425), .A2(n528), .B1(n482), .B2(n742), .C1(n481), .C2(
        n746), .ZN(n486) );
  AOI221D1 U2 ( .A1(n787), .A2(n674), .B1(n673), .B2(n795), .C(n672), .ZN(n675) );
  ND2D1 U3 ( .A1(n429), .A2(n823), .ZN(n748) );
  INVD3 U4 ( .I(a[6]), .ZN(n823) );
  INR4D1 U5 ( .A1(n661), .B1(n844), .B2(n659), .B3(n660), .ZN(n670) );
  INVD3 U6 ( .I(n427), .ZN(n789) );
  AN2D2 U7 ( .A1(n431), .A2(n789), .Z(n306) );
  CKND2D1 U8 ( .A1(n789), .A2(n438), .ZN(n676) );
  CKND2D0 U9 ( .A1(n789), .A2(n808), .ZN(n547) );
  CKND2D0 U10 ( .A1(n431), .A2(n789), .ZN(n424) );
  CKND2D2 U11 ( .A1(n428), .A2(n437), .ZN(n741) );
  AOI221D1 U12 ( .A1(n790), .A2(n813), .B1(n798), .B2(n820), .C(n757), .ZN(
        n772) );
  NR4D1 U13 ( .A1(n778), .A2(n779), .A3(n780), .A4(n777), .ZN(n781) );
  ND2D2 U14 ( .A1(n433), .A2(n436), .ZN(n735) );
  CKND0 U15 ( .I(n735), .ZN(n786) );
  AOI221D1 U16 ( .A1(n684), .A2(n735), .B1(n434), .B2(n843), .C(n550), .ZN(
        n555) );
  OAI21D1 U17 ( .A1(n742), .A2(n602), .B(n712), .ZN(n583) );
  CKND4 U18 ( .I(a[1]), .ZN(n436) );
  ND2D1 U19 ( .A1(n811), .A2(n837), .ZN(n597) );
  INVD2 U20 ( .I(n740), .ZN(n811) );
  AOI221D2 U21 ( .A1(n811), .A2(n786), .B1(n820), .B2(n797), .C(n553), .ZN(
        n554) );
  AOI221D1 U22 ( .A1(n825), .A2(n813), .B1(n811), .B2(n563), .C(n840), .ZN(
        n489) );
  CKND2D2 U23 ( .A1(n823), .A2(n828), .ZN(n742) );
  INVD4 U24 ( .I(n429), .ZN(n828) );
  ND2D1 U25 ( .A1(n437), .A2(n808), .ZN(n740) );
  INVD2 U26 ( .I(n748), .ZN(n848) );
  ND2D1 U27 ( .A1(a[6]), .A2(n828), .ZN(n771) );
  CKND2D2 U29 ( .A1(n435), .A2(n430), .ZN(n710) );
  ND2D1 U30 ( .A1(n439), .A2(n808), .ZN(n746) );
  ND2D2 U31 ( .A1(n434), .A2(n433), .ZN(n729) );
  INVD1 U32 ( .I(n742), .ZN(n834) );
  INVD1 U33 ( .I(n668), .ZN(n807) );
  OAI31D1 U34 ( .A1(n663), .A2(n306), .A3(n807), .B(n662), .ZN(n664) );
  ND2D2 U36 ( .A1(a[5]), .A2(n808), .ZN(n756) );
  NR2D1 U37 ( .A1(n808), .A2(n816), .ZN(n662) );
  ND2D1 U38 ( .A1(n792), .A2(n433), .ZN(n548) );
  INVD1 U39 ( .I(n548), .ZN(n793) );
  NR2D0 U40 ( .A1(n432), .A2(n437), .ZN(n663) );
  INVD1 U41 ( .I(n743), .ZN(n790) );
  CKND2D1 U42 ( .A1(n437), .A2(a[5]), .ZN(n677) );
  INVD1 U43 ( .I(n738), .ZN(n797) );
  INVD2 U44 ( .I(a[5]), .ZN(n816) );
  INVD2 U45 ( .I(n304), .ZN(n305) );
  INVD2 U46 ( .I(n656), .ZN(n795) );
  ND2D2 U47 ( .A1(n436), .A2(n789), .ZN(n743) );
  INVD2 U48 ( .I(n432), .ZN(n431) );
  CKND2D0 U49 ( .A1(n433), .A2(n789), .ZN(n754) );
  CKND2D1 U50 ( .A1(n434), .A2(n437), .ZN(n773) );
  INVD3 U51 ( .I(n436), .ZN(n435) );
  ND4D1 U52 ( .A1(n615), .A2(n614), .A3(n613), .A4(n612), .ZN(d[3]) );
  AOI221D1 U53 ( .A1(n455), .A2(n797), .B1(n841), .B2(n806), .C(n454), .ZN(
        n456) );
  NR4D0 U54 ( .A1(n526), .A2(n525), .A3(n524), .A4(n585), .ZN(n527) );
  ND2D1 U55 ( .A1(n818), .A2(n837), .ZN(n588) );
  AOI21D1 U56 ( .A1(n803), .A2(n434), .B(n793), .ZN(n575) );
  OAI222D0 U57 ( .A1(n736), .A2(n710), .B1(n760), .B2(n574), .C1(n741), .C2(
        n751), .ZN(n578) );
  NR2D1 U58 ( .A1(n822), .A2(n818), .ZN(n665) );
  ND2D1 U59 ( .A1(n437), .A2(n436), .ZN(n668) );
  ND2D1 U60 ( .A1(a[6]), .A2(n816), .ZN(n764) );
  AOI221D0 U61 ( .A1(n788), .A2(n679), .B1(n822), .B2(n306), .C(n678), .ZN(
        n680) );
  ND2D1 U62 ( .A1(n837), .A2(n821), .ZN(n627) );
  ND2D1 U63 ( .A1(n808), .A2(n816), .ZN(n760) );
  INVD1 U64 ( .I(n676), .ZN(n803) );
  AOI221D0 U65 ( .A1(n824), .A2(n785), .B1(n583), .B2(n436), .C(n725), .ZN(
        n584) );
  ND2D1 U66 ( .A1(n831), .A2(n817), .ZN(n712) );
  INVD4 U67 ( .I(n430), .ZN(n433) );
  OAI22D1 U68 ( .A1(n436), .A2(n622), .B1(n621), .B2(n734), .ZN(n623) );
  ND2D1 U69 ( .A1(n831), .A2(n662), .ZN(n722) );
  CKAN2D0 U70 ( .A1(n528), .A2(n722), .Z(n461) );
  AOI221D0 U71 ( .A1(n850), .A2(n436), .B1(n832), .B2(n710), .C(n520), .ZN(
        n523) );
  OAI31D2 U72 ( .A1(n696), .A2(a[5]), .A3(n434), .B(n628), .ZN(n550) );
  AOI21D1 U73 ( .A1(n850), .A2(n805), .B(n844), .ZN(n558) );
  NR2D1 U74 ( .A1(n694), .A2(n735), .ZN(n725) );
  OAI222D2 U75 ( .A1(n656), .A2(n759), .B1(n430), .B2(n552), .C1(n741), .C2(
        n551), .ZN(n553) );
  INVD2 U76 ( .I(a[3]), .ZN(n438) );
  INVD1 U77 ( .I(n655), .ZN(n835) );
  INVD4 U78 ( .I(n432), .ZN(n430) );
  INVD3 U79 ( .I(a[0]), .ZN(n432) );
  AOI22D1 U80 ( .A1(n827), .A2(n795), .B1(n798), .B2(n826), .ZN(n462) );
  OR2XD1 U81 ( .A1(n522), .A2(n710), .Z(n277) );
  AOI22D2 U82 ( .A1(n819), .A2(n805), .B1(n795), .B2(n816), .ZN(n552) );
  ND2D2 U83 ( .A1(n427), .A2(n436), .ZN(n656) );
  ND2D1 U84 ( .A1(n797), .A2(n433), .ZN(n697) );
  OAI22D0 U85 ( .A1(n462), .A2(n305), .B1(n461), .B2(n751), .ZN(n463) );
  OAI221D1 U86 ( .A1(n601), .A2(n576), .B1(n437), .B2(n765), .C(n693), .ZN(
        n521) );
  ND2D1 U87 ( .A1(n662), .A2(n848), .ZN(n765) );
  OAI222D1 U89 ( .A1(n800), .A2(n622), .B1(n548), .B2(n528), .C1(n527), .C2(
        n771), .ZN(n534) );
  OAI221D1 U90 ( .A1(n658), .A2(n668), .B1(n657), .B2(n656), .C(n835), .ZN(
        n660) );
  OAI222D1 U91 ( .A1(n425), .A2(n740), .B1(n681), .B2(n677), .C1(n746), .C2(
        n548), .ZN(n526) );
  NR2XD0 U92 ( .A1(n306), .A2(n787), .ZN(n681) );
  OAI22D1 U93 ( .A1(n756), .A2(n766), .B1(n434), .B2(n755), .ZN(n757) );
  CKND2D1 U94 ( .A1(n429), .A2(n816), .ZN(n718) );
  AOI221D1 U95 ( .A1(n834), .A2(n451), .B1(n450), .B2(n433), .C(n449), .ZN(
        n474) );
  ND2D2 U96 ( .A1(n437), .A2(n427), .ZN(n633) );
  AOI211XD0 U97 ( .A1(n807), .A2(n431), .B(n805), .C(n799), .ZN(n595) );
  OA221D1 U98 ( .A1(n551), .A2(n622), .B1(n710), .B2(n775), .C(n51), .Z(n615)
         );
  OA222D1 U99 ( .A1(n633), .A2(n626), .B1(n582), .B2(n581), .C1(n580), .C2(
        n748), .Z(n51) );
  CKND1 U100 ( .I(n710), .ZN(n785) );
  CKND2D1 U101 ( .A1(n816), .A2(n823), .ZN(n647) );
  INVD3 U102 ( .I(n436), .ZN(n434) );
  AOI221D1 U103 ( .A1(n790), .A2(n847), .B1(n799), .B2(n826), .C(n453), .ZN(
        n457) );
  AO21D0 U104 ( .A1(n787), .A2(n824), .B(n725), .Z(n453) );
  OAI222D1 U105 ( .A1(n721), .A2(n711), .B1(n689), .B2(n433), .C1(n688), .C2(
        n764), .ZN(n690) );
  INVD2 U106 ( .I(n696), .ZN(n837) );
  ND2D2 U107 ( .A1(n429), .A2(a[6]), .ZN(n696) );
  ND2D2 U108 ( .A1(n819), .A2(n837), .ZN(n721) );
  NR2D1 U109 ( .A1(n826), .A2(n837), .ZN(n630) );
  ND2D1 U110 ( .A1(n817), .A2(n837), .ZN(n626) );
  AOI221D1 U111 ( .A1(n831), .A2(n491), .B1(n791), .B2(n504), .C(n490), .ZN(
        n500) );
  ND4D2 U112 ( .A1(n572), .A2(n573), .A3(n571), .A4(n570), .ZN(d[4]) );
  ND2D0 U113 ( .A1(a[5]), .A2(n438), .ZN(n759) );
  OA221D1 U114 ( .A1(n432), .A2(n65), .B1(n771), .B2(n70), .C(n72), .Z(n572)
         );
  OA211D0 U115 ( .A1(n694), .A2(n668), .B(n543), .C(n542), .Z(n65) );
  OA211D0 U116 ( .A1(n547), .A2(n710), .B(n546), .C(n545), .Z(n70) );
  OA222D1 U117 ( .A1(n556), .A2(n748), .B1(n676), .B2(n555), .C1(n742), .C2(
        n554), .Z(n72) );
  INVD2 U118 ( .I(n771), .ZN(n831) );
  AOI211XD0 U119 ( .A1(n852), .A2(n798), .B(n475), .C(n655), .ZN(n502) );
  ND2D2 U120 ( .A1(n841), .A2(n433), .ZN(n628) );
  AOI221D1 U121 ( .A1(n845), .A2(n785), .B1(n848), .B2(n683), .C(n682), .ZN(
        n707) );
  AOI222D1 U122 ( .A1(n797), .A2(n819), .B1(n795), .B2(n477), .C1(n791), .C2(
        n822), .ZN(n482) );
  OA221D1 U123 ( .A1(n676), .A2(n666), .B1(n665), .B2(n776), .C(n664), .Z(n426) );
  OA21D0 U124 ( .A1(n676), .A2(n433), .B(n605), .Z(n609) );
  OAI22D1 U125 ( .A1(n714), .A2(n743), .B1(n789), .B2(n720), .ZN(n655) );
  OAI222D1 U126 ( .A1(n457), .A2(n740), .B1(n677), .B2(n508), .C1(n433), .C2(
        n456), .ZN(n458) );
  ND2D2 U127 ( .A1(n790), .A2(n430), .ZN(n551) );
  CKND0 U128 ( .I(n718), .ZN(n847) );
  OAI33D0 U129 ( .A1(n647), .A2(n431), .A3(n789), .B1(n478), .B2(n718), .B3(
        n751), .ZN(n479) );
  AOI221D1 U130 ( .A1(n836), .A2(n433), .B1(n846), .B2(n434), .C(n631), .ZN(
        n632) );
  OAI22D0 U131 ( .A1(n735), .A2(n698), .B1(n630), .B2(n729), .ZN(n631) );
  CKND1 U132 ( .I(n774), .ZN(n836) );
  OAI211D0 U133 ( .A1(n816), .A2(n746), .B(n763), .C(n741), .ZN(n674) );
  OAI222D1 U134 ( .A1(n772), .A2(n771), .B1(n437), .B2(n829), .C1(n770), .C2(
        n433), .ZN(n778) );
  INVD0 U135 ( .I(n751), .ZN(n799) );
  ND2D1 U136 ( .A1(n431), .A2(n427), .ZN(n751) );
  INVD2 U137 ( .I(n633), .ZN(n805) );
  AOI221D1 U138 ( .A1(n811), .A2(n848), .B1(n801), .B2(n821), .C(n521), .ZN(
        n522) );
  INVD4 U139 ( .I(n776), .ZN(n792) );
  ND2D4 U140 ( .A1(n435), .A2(n789), .ZN(n776) );
  AOI211XD1 U141 ( .A1(n818), .A2(n579), .B(n577), .C(n578), .ZN(n580) );
  INVD6 U142 ( .I(n428), .ZN(n808) );
  INVD2 U143 ( .I(n756), .ZN(n821) );
  AOI221D1 U144 ( .A1(n802), .A2(n563), .B1(n562), .B2(n811), .C(n561), .ZN(
        n571) );
  OAI222D1 U145 ( .A1(n634), .A2(n633), .B1(n751), .B2(n753), .C1(n632), .C2(
        n763), .ZN(n635) );
  AOI211XD0 U146 ( .A1(n793), .A2(n812), .B(n815), .C(n687), .ZN(n688) );
  INVD4 U147 ( .I(n438), .ZN(n437) );
  ND2D2 U148 ( .A1(n437), .A2(n816), .ZN(n737) );
  ND2D2 U149 ( .A1(n437), .A2(n789), .ZN(n763) );
  OAI222D1 U150 ( .A1(n430), .A2(n670), .B1(n669), .B2(n742), .C1(n668), .C2(
        n667), .ZN(n671) );
  AOI221D1 U151 ( .A1(n834), .A2(n600), .B1(n599), .B2(n433), .C(n598), .ZN(
        n613) );
  OA221D1 U152 ( .A1(n737), .A2(n729), .B1(n746), .B2(n656), .C(n426), .Z(n669) );
  OR2XD1 U153 ( .A1(n523), .A2(n766), .Z(n142) );
  OR2D0 U154 ( .A1(n424), .A2(n616), .Z(n192) );
  ND3D1 U155 ( .A1(n142), .A2(n192), .A3(n277), .ZN(n535) );
  ND2D1 U156 ( .A1(n821), .A2(n828), .ZN(n616) );
  NR4D1 U157 ( .A1(n536), .A2(n535), .A3(n534), .A4(n533), .ZN(n537) );
  AOI221D1 U158 ( .A1(n434), .A2(n459), .B1(n815), .B2(n825), .C(n458), .ZN(
        n473) );
  INVD1 U159 ( .I(n701), .ZN(n304) );
  AOI221D1 U160 ( .A1(n848), .A2(n636), .B1(n845), .B2(n792), .C(n635), .ZN(
        n653) );
  AOI221D1 U161 ( .A1(n592), .A2(n804), .B1(n831), .B2(n591), .C(n590), .ZN(
        n614) );
  AOI221D1 U162 ( .A1(n839), .A2(n799), .B1(n684), .B2(n792), .C(n671), .ZN(
        n708) );
  NR2D0 U163 ( .A1(n503), .A2(n656), .ZN(n562) );
  ND2D0 U164 ( .A1(n816), .A2(n828), .ZN(n601) );
  ND2D0 U165 ( .A1(a[5]), .A2(n828), .ZN(n698) );
  CKND2D0 U166 ( .A1(n434), .A2(a[6]), .ZN(n478) );
  ND2D0 U167 ( .A1(n819), .A2(n848), .ZN(n667) );
  OAI22D0 U168 ( .A1(n436), .A2(n712), .B1(n434), .B2(n627), .ZN(n629) );
  AOI211XD0 U169 ( .A1(n848), .A2(n487), .B(n486), .C(n485), .ZN(n501) );
  BUFFD4 U170 ( .I(a[7]), .Z(n429) );
  ND2D1 U171 ( .A1(n801), .A2(n434), .ZN(n574) );
  NR2D0 U172 ( .A1(n616), .A2(n734), .ZN(n758) );
  CKND2D0 U173 ( .A1(n788), .A2(n848), .ZN(n508) );
  CKND0 U174 ( .I(n712), .ZN(n833) );
  CKND2D0 U175 ( .A1(n677), .A2(n740), .ZN(n679) );
  CKND2D0 U176 ( .A1(n754), .A2(n751), .ZN(n739) );
  CKND2D0 U177 ( .A1(n673), .A2(n837), .ZN(n622) );
  CKND2D0 U178 ( .A1(n662), .A2(n837), .ZN(n581) );
  CKND0 U179 ( .I(n694), .ZN(n851) );
  NR2XD0 U180 ( .A1(n849), .A2(n504), .ZN(n505) );
  NR2D0 U181 ( .A1(n799), .A2(n797), .ZN(n460) );
  INR2D0 U182 ( .A1(n752), .B1(n493), .ZN(n494) );
  ND2D0 U183 ( .A1(a[5]), .A2(n823), .ZN(n503) );
  OAI31D0 U184 ( .A1(n790), .A2(n787), .A3(n801), .B(n849), .ZN(n483) );
  AOI22D0 U185 ( .A1(n850), .A2(n792), .B1(n806), .B2(n836), .ZN(n542) );
  NR2D0 U186 ( .A1(n433), .A2(n750), .ZN(n732) );
  NR2D0 U187 ( .A1(n794), .A2(n790), .ZN(n467) );
  ND2D0 U188 ( .A1(n801), .A2(n843), .ZN(n557) );
  NR2D0 U189 ( .A1(n801), .A2(n794), .ZN(n441) );
  CKND0 U190 ( .I(n551), .ZN(n791) );
  NR2D0 U191 ( .A1(n709), .A2(n846), .ZN(n716) );
  OAI22D0 U192 ( .A1(n433), .A2(n712), .B1(n436), .B2(n722), .ZN(n520) );
  CKND2D0 U193 ( .A1(n773), .A2(n548), .ZN(n549) );
  ND3D0 U194 ( .A1(n805), .A2(n662), .A3(n834), .ZN(n750) );
  OAI22D0 U195 ( .A1(n746), .A2(n743), .B1(n646), .B2(n729), .ZN(n512) );
  CKND2D0 U196 ( .A1(n773), .A2(n676), .ZN(n517) );
  CKND2D0 U197 ( .A1(n424), .A2(n743), .ZN(n518) );
  NR2D0 U198 ( .A1(n721), .A2(n437), .ZN(n686) );
  OAI22D0 U200 ( .A1(n734), .A2(n746), .B1(n593), .B2(n735), .ZN(n600) );
  NR2D0 U201 ( .A1(n814), .A2(n819), .ZN(n593) );
  AOI22D0 U202 ( .A1(n433), .A2(n806), .B1(n439), .B2(n794), .ZN(n582) );
  ND2D0 U203 ( .A1(n834), .A2(n821), .ZN(n774) );
  AOI22D0 U204 ( .A1(n797), .A2(n430), .B1(n434), .B2(n805), .ZN(n476) );
  CKND2D0 U205 ( .A1(n431), .A2(n795), .ZN(n719) );
  NR2D0 U206 ( .A1(n805), .A2(n812), .ZN(n646) );
  AOI31D0 U207 ( .A1(n722), .A2(n721), .A3(n720), .B(n719), .ZN(n723) );
  CKND2D0 U208 ( .A1(n804), .A2(n434), .ZN(n711) );
  AOI22D0 U210 ( .A1(n818), .A2(n795), .B1(n792), .B2(n820), .ZN(n440) );
  NR2D0 U211 ( .A1(n627), .A2(n713), .ZN(n731) );
  NR2D0 U212 ( .A1(n797), .A2(n785), .ZN(n605) );
  CKND2D0 U213 ( .A1(n851), .A2(n813), .ZN(n775) );
  ND2D0 U214 ( .A1(n811), .A2(n851), .ZN(n752) );
  NR2D0 U216 ( .A1(n306), .A2(n786), .ZN(n606) );
  CKND2D0 U218 ( .A1(n810), .A2(n834), .ZN(n661) );
  ND2D0 U219 ( .A1(n819), .A2(n436), .ZN(n666) );
  CKND2D0 U220 ( .A1(n824), .A2(n813), .ZN(n528) );
  NR2D0 U221 ( .A1(n786), .A2(n795), .ZN(n641) );
  NR2D0 U222 ( .A1(n846), .A2(n684), .ZN(n444) );
  CKND2D0 U223 ( .A1(n306), .A2(n821), .ZN(n637) );
  AOI211XD0 U224 ( .A1(n832), .A2(n431), .B(n629), .C(n842), .ZN(n634) );
  CKND2D0 U225 ( .A1(n719), .A2(n729), .ZN(n579) );
  CKND0 U226 ( .I(n574), .ZN(n802) );
  NR2D0 U227 ( .A1(n850), .A2(n836), .ZN(n452) );
  OAI22D0 U228 ( .A1(n756), .A2(n676), .B1(n681), .B2(n305), .ZN(n446) );
  AOI21D0 U229 ( .A1(n676), .A2(n576), .B(n734), .ZN(n445) );
  CKND2D0 U230 ( .A1(n805), .A2(n808), .ZN(n594) );
  OAI22D0 U231 ( .A1(n737), .A2(n743), .B1(n756), .B2(n776), .ZN(n678) );
  OAI33D0 U232 ( .A1(n746), .A2(n789), .A3(n718), .B1(n647), .B2(n434), .B3(
        n646), .ZN(n650) );
  NR2D0 U233 ( .A1(n742), .A2(n760), .ZN(n684) );
  OAI32D0 U234 ( .A1(n551), .A2(n748), .A3(n737), .B1(n509), .B2(n508), .ZN(
        n510) );
  NR2D0 U235 ( .A1(n821), .A2(n801), .ZN(n509) );
  OAI22D0 U236 ( .A1(n776), .A2(n775), .B1(n774), .B2(n773), .ZN(n777) );
  CKND2D1 U237 ( .A1(n484), .A2(n483), .ZN(n485) );
  AOI22D0 U238 ( .A1(n801), .A2(n821), .B1(n803), .B2(n816), .ZN(n755) );
  AOI32D0 U239 ( .A1(n790), .A2(n433), .A3(n822), .B1(n788), .B2(n544), .ZN(
        n546) );
  OAI31D0 U240 ( .A1(n729), .A2(n812), .A3(n742), .B(n728), .ZN(n733) );
  OAI21D0 U241 ( .A1(n741), .A2(n601), .B(n626), .ZN(n504) );
  AOI21D0 U242 ( .A1(n602), .A2(n647), .B(n676), .ZN(n493) );
  AOI22D0 U243 ( .A1(n825), .A2(n739), .B1(n827), .B2(n795), .ZN(n747) );
  AOI22D0 U244 ( .A1(n798), .A2(n847), .B1(n790), .B2(n826), .ZN(n560) );
  CKND0 U245 ( .I(a[3]), .ZN(n439) );
  CKND2D0 U246 ( .A1(n820), .A2(n837), .ZN(n753) );
  NR2XD0 U247 ( .A1(n638), .A2(n758), .ZN(n596) );
  AOI32D0 U248 ( .A1(a[5]), .A2(n433), .A3(n806), .B1(n817), .B2(n624), .ZN(
        n625) );
  AOI21D0 U249 ( .A1(n796), .A2(n834), .B(n562), .ZN(n506) );
  NR2D0 U250 ( .A1(n799), .A2(n437), .ZN(n608) );
  AOI21D0 U251 ( .A1(n811), .A2(n847), .B(n686), .ZN(n496) );
  CKND2D1 U252 ( .A1(n429), .A2(n492), .ZN(n495) );
  CKND0 U253 ( .I(n758), .ZN(n829) );
  NR2XD0 U254 ( .A1(n769), .A2(n768), .ZN(n770) );
  NR2D0 U255 ( .A1(n793), .A2(n796), .ZN(n566) );
  OAI21D0 U256 ( .A1(n647), .A2(n740), .B(n720), .ZN(n531) );
  AOI21D0 U257 ( .A1(n846), .A2(n806), .B(n686), .ZN(n689) );
  AOI21D0 U258 ( .A1(n845), .A2(n434), .B(n684), .ZN(n685) );
  ND4D0 U259 ( .A1(n787), .A2(n825), .A3(n428), .A4(n429), .ZN(n717) );
  CKND2D0 U260 ( .A1(n428), .A2(n438), .ZN(n701) );
  OAI32D0 U261 ( .A1(n759), .A2(n467), .A3(n696), .B1(n466), .B2(n729), .ZN(
        n470) );
  AOI31D0 U262 ( .A1(n428), .A2(n823), .A3(n801), .B(n686), .ZN(n466) );
  AOI211D0 U263 ( .A1(n767), .A2(n647), .B(n576), .C(n734), .ZN(n468) );
  NR2D0 U264 ( .A1(n437), .A2(a[5]), .ZN(n673) );
  AOI211XD0 U265 ( .A1(n830), .A2(n798), .B(n480), .C(n479), .ZN(n481) );
  CKND0 U266 ( .I(n601), .ZN(n830) );
  AOI32D0 U267 ( .A1(n429), .A2(n808), .A3(n790), .B1(n795), .B2(n442), .ZN(
        n443) );
  OAI22D0 U268 ( .A1(n429), .A2(n647), .B1(n741), .B2(n718), .ZN(n442) );
  CKND2D0 U269 ( .A1(n428), .A2(n789), .ZN(n576) );
  AOI22D0 U270 ( .A1(n792), .A2(n825), .B1(n801), .B2(n808), .ZN(n762) );
  CKND2D1 U271 ( .A1(n587), .A2(n586), .ZN(n591) );
  AOI21D0 U272 ( .A1(n836), .A2(n805), .B(n744), .ZN(n745) );
  OAI33D0 U273 ( .A1(n743), .A2(n742), .A3(n741), .B1(n764), .B2(n789), .B3(
        n740), .ZN(n744) );
  AOI21D0 U274 ( .A1(n785), .A2(n639), .B(n638), .ZN(n642) );
  OAI22D0 U275 ( .A1(n823), .A2(n305), .B1(n808), .B2(n647), .ZN(n639) );
  CKND2D1 U276 ( .A1(n764), .A2(n718), .ZN(n563) );
  OAI21D0 U277 ( .A1(n700), .A2(n729), .B(n699), .ZN(n704) );
  OA33D0 U278 ( .A1(n698), .A2(n741), .A3(n734), .B1(n697), .B2(n696), .B3(
        n759), .Z(n699) );
  NR2D0 U279 ( .A1(n428), .A2(n823), .ZN(n455) );
  CKND2D0 U280 ( .A1(a[5]), .A2(a[6]), .ZN(n767) );
  AOI32D0 U281 ( .A1(n428), .A2(n828), .A3(n804), .B1(n805), .B2(n541), .ZN(
        n543) );
  OAI22D0 U282 ( .A1(a[6]), .A2(n428), .B1(a[5]), .B2(n748), .ZN(n541) );
  BUFFD4 U283 ( .I(a[4]), .Z(n428) );
  BUFFD4 U284 ( .I(a[2]), .Z(n427) );
  INVD1 U285 ( .I(n773), .ZN(n806) );
  INVD1 U287 ( .I(n557), .ZN(n844) );
  INVD1 U288 ( .I(n697), .ZN(n798) );
  INVD1 U289 ( .I(n667), .ZN(n850) );
  INVD1 U290 ( .I(n734), .ZN(n787) );
  INVD1 U291 ( .I(n765), .ZN(n849) );
  INVD1 U292 ( .I(n719), .ZN(n796) );
  INVD1 U293 ( .I(n589), .ZN(n815) );
  INVD1 U294 ( .I(n775), .ZN(n852) );
  AOI222D0 U295 ( .A1(n797), .A2(n813), .B1(n811), .B2(n306), .C1(n820), .C2(
        n795), .ZN(n545) );
  INVD1 U296 ( .I(n628), .ZN(n842) );
  INVD1 U297 ( .I(n763), .ZN(n801) );
  INVD1 U298 ( .I(n581), .ZN(n846) );
  INVD1 U299 ( .I(n626), .ZN(n845) );
  NR2D1 U300 ( .A1(n750), .A2(n431), .ZN(n703) );
  NR3D0 U301 ( .A1(n663), .A2(n790), .A3(n804), .ZN(n640) );
  INVD1 U302 ( .I(n754), .ZN(n794) );
  ND2D1 U303 ( .A1(n431), .A2(n436), .ZN(n734) );
  INVD1 U304 ( .I(n588), .ZN(n840) );
  INVD1 U305 ( .I(n714), .ZN(n832) );
  INVD1 U306 ( .I(n760), .ZN(n817) );
  ND2D1 U307 ( .A1(n785), .A2(n814), .ZN(n589) );
  INVD1 U308 ( .I(n721), .ZN(n841) );
  INVD1 U309 ( .I(n627), .ZN(n843) );
  ND2D1 U310 ( .A1(n809), .A2(n825), .ZN(n693) );
  INVD1 U311 ( .I(n737), .ZN(n818) );
  INVD1 U312 ( .I(n547), .ZN(n809) );
  INVD1 U313 ( .I(n597), .ZN(n838) );
  INVD1 U314 ( .I(n622), .ZN(n839) );
  OAI222D0 U315 ( .A1(n716), .A2(n424), .B1(n715), .B2(n714), .C1(n713), .C2(
        n712), .ZN(n784) );
  NR4D0 U316 ( .A1(n447), .A2(n446), .A3(n524), .A4(n445), .ZN(n448) );
  OAI222D0 U317 ( .A1(n560), .A2(n305), .B1(n559), .B2(n734), .C1(n434), .C2(
        n558), .ZN(n561) );
  AOI21D1 U318 ( .A1(n809), .A2(n851), .B(n838), .ZN(n559) );
  OAI222D0 U319 ( .A1(n425), .A2(n588), .B1(n722), .B2(n668), .C1(n627), .C2(
        n751), .ZN(n540) );
  OAI21D1 U320 ( .A1(n430), .A2(n677), .B(n740), .ZN(n477) );
  OAI222D0 U321 ( .A1(n749), .A2(n748), .B1(n747), .B2(n746), .C1(n431), .C2(
        n745), .ZN(n780) );
  NR2XD0 U322 ( .A1(n832), .A2(n843), .ZN(n658) );
  AOI21D1 U323 ( .A1(n822), .A2(n831), .B(n840), .ZN(n657) );
  NR4D0 U324 ( .A1(n305), .A2(n754), .A3(n748), .A4(n816), .ZN(n726) );
  AOI221D0 U325 ( .A1(n785), .A2(n803), .B1(n791), .B2(n818), .C(n585), .ZN(
        n586) );
  INVD1 U326 ( .I(n759), .ZN(n822) );
  ND2D1 U327 ( .A1(n741), .A2(n736), .ZN(n544) );
  OAI222D0 U328 ( .A1(n743), .A2(n677), .B1(n476), .B2(n756), .C1(n434), .C2(
        n741), .ZN(n487) );
  INVD1 U329 ( .I(n647), .ZN(n825) );
  INVD1 U330 ( .I(n305), .ZN(n813) );
  NR3D0 U331 ( .A1(n710), .A2(n808), .A3(n720), .ZN(n567) );
  NR3D0 U332 ( .A1(n729), .A2(n437), .A3(n756), .ZN(n525) );
  INVD1 U333 ( .I(n602), .ZN(n819) );
  ND2D1 U334 ( .A1(n819), .A2(n831), .ZN(n714) );
  INVD1 U335 ( .I(n677), .ZN(n820) );
  ND2D1 U336 ( .A1(n673), .A2(n834), .ZN(n720) );
  NR3D0 U337 ( .A1(n503), .A2(n741), .A3(n776), .ZN(n469) );
  INVD1 U338 ( .I(n741), .ZN(n812) );
  NR2D1 U339 ( .A1(n698), .A2(n305), .ZN(n709) );
  INVD1 U340 ( .I(n503), .ZN(n824) );
  OAI222D0 U341 ( .A1(n743), .A2(n597), .B1(n596), .B2(n789), .C1(n595), .C2(
        n667), .ZN(n598) );
  OAI221D0 U342 ( .A1(n606), .A2(n756), .B1(n741), .B2(n751), .C(n488), .ZN(
        n491) );
  AOI221D0 U343 ( .A1(n831), .A2(n645), .B1(n834), .B2(n644), .C(n643), .ZN(
        n652) );
  AO221D0 U344 ( .A1(n790), .A2(n822), .B1(n788), .B2(n804), .C(n692), .Z(n644) );
  OAI222D0 U345 ( .A1(n427), .A2(n642), .B1(n641), .B2(n775), .C1(n640), .C2(
        n774), .ZN(n643) );
  OAI221D0 U346 ( .A1(n729), .A2(n722), .B1(n696), .B2(n735), .C(n584), .ZN(
        n592) );
  OAI222D0 U347 ( .A1(n718), .A2(n589), .B1(n425), .B2(n753), .C1(n605), .C2(
        n588), .ZN(n590) );
  NR4D0 U348 ( .A1(n435), .A2(n828), .A3(n754), .A4(n746), .ZN(n687) );
  OAI222D0 U349 ( .A1(n467), .A2(n698), .B1(n460), .B2(n696), .C1(n718), .C2(
        n719), .ZN(n464) );
  OAI222D0 U350 ( .A1(n429), .A2(n762), .B1(n761), .B2(n760), .C1(n771), .C2(
        n759), .ZN(n769) );
  AOI222D0 U351 ( .A1(n792), .A2(n810), .B1(n812), .B2(n794), .C1(n796), .C2(
        a[5]), .ZN(n587) );
  OAI222D0 U352 ( .A1(n507), .A2(n734), .B1(n506), .B2(n741), .C1(n505), .C2(
        n754), .ZN(n511) );
  OAI222D0 U353 ( .A1(n609), .A2(n765), .B1(n608), .B2(n714), .C1(n607), .C2(
        n746), .ZN(n610) );
  OA22D0 U354 ( .A1(n767), .A2(n734), .B1(n718), .B2(n606), .Z(n607) );
  OAI222D0 U355 ( .A1(n496), .A2(n735), .B1(n808), .B2(n495), .C1(n494), .C2(
        n710), .ZN(n498) );
  NR3D0 U356 ( .A1(n433), .A2(n428), .A3(n677), .ZN(n585) );
  OAI222D0 U357 ( .A1(n697), .A2(n722), .B1(n430), .B2(n532), .C1(n776), .C2(
        n765), .ZN(n533) );
  AOI221D0 U358 ( .A1(n795), .A2(n531), .B1(n834), .B2(n530), .C(n529), .ZN(
        n532) );
  OAI221D0 U359 ( .A1(n729), .A2(n718), .B1(n435), .B2(n774), .C(n717), .ZN(
        n724) );
  OAI221D0 U360 ( .A1(n433), .A2(n722), .B1(n696), .B2(n710), .C(n685), .ZN(
        n691) );
  OAI221D0 U361 ( .A1(n741), .A2(n743), .B1(n305), .B2(n776), .C(n625), .ZN(
        n636) );
  OAI221D0 U362 ( .A1(n434), .A2(n661), .B1(n713), .B2(n667), .C(n519), .ZN(
        n536) );
  OAI221D0 U363 ( .A1(n441), .A2(n602), .B1(n766), .B2(n710), .C(n440), .ZN(
        n451) );
  NR3D0 U364 ( .A1(n729), .A2(n428), .A3(n601), .ZN(n638) );
  NR4D0 U365 ( .A1(n431), .A2(n823), .A3(n760), .A4(n766), .ZN(n568) );
  NR4D0 U366 ( .A1(n620), .A2(n619), .A3(n838), .A4(n618), .ZN(n621) );
  OAI222D0 U367 ( .A1(n434), .A2(n767), .B1(n735), .B2(n748), .C1(n742), .C2(
        n738), .ZN(n480) );
  NR3D0 U368 ( .A1(n696), .A2(n816), .A3(n305), .ZN(n515) );
  NR3D0 U369 ( .A1(n711), .A2(n428), .A3(n828), .ZN(n649) );
  ND2D1 U370 ( .A1(a[5]), .A2(n429), .ZN(n694) );
  INVD1 U371 ( .I(n764), .ZN(n826) );
  ND2D1 U372 ( .A1(n428), .A2(n816), .ZN(n602) );
  INVD1 U373 ( .I(n767), .ZN(n827) );
  OAI221D0 U374 ( .A1(n729), .A2(n676), .B1(n737), .B2(n695), .C(n675), .ZN(
        n683) );
  OAI222D0 U375 ( .A1(n743), .A2(n752), .B1(n681), .B2(n712), .C1(n680), .C2(
        n771), .ZN(n682) );
  NR4D0 U376 ( .A1(a[6]), .A2(n439), .A3(n718), .A4(n751), .ZN(n497) );
  ND3D1 U377 ( .A1(n539), .A2(n538), .A3(n537), .ZN(d[5]) );
  AOI211D1 U378 ( .A1(n851), .A2(n512), .B(n511), .C(n510), .ZN(n539) );
  INR4D0 U379 ( .A1(n750), .B1(n516), .B2(n731), .B3(n702), .ZN(n538) );
  NR2D1 U380 ( .A1(n611), .A2(n610), .ZN(n612) );
  NR4D0 U381 ( .A1(n470), .A2(n469), .A3(n703), .A4(n468), .ZN(n471) );
  AOI221D0 U382 ( .A1(n465), .A2(n436), .B1(n810), .B2(n464), .C(n463), .ZN(
        n472) );
  NR4D0 U383 ( .A1(n733), .A2(n732), .A3(n731), .A4(n730), .ZN(n782) );
  AOI221D0 U384 ( .A1(n725), .A2(n804), .B1(n803), .B2(n724), .C(n723), .ZN(
        n783) );
  ND4D1 U385 ( .A1(n654), .A2(n653), .A3(n652), .A4(n651), .ZN(d[2]) );
  NR4D0 U386 ( .A1(n650), .A2(n649), .A3(n648), .A4(n732), .ZN(n651) );
  AOI221D0 U387 ( .A1(n849), .A2(n433), .B1(n841), .B2(n797), .C(n623), .ZN(
        n654) );
  ND4D1 U388 ( .A1(n708), .A2(n707), .A3(n706), .A4(n705), .ZN(d[1]) );
  NR4D0 U389 ( .A1(n704), .A2(n726), .A3(n703), .A4(n702), .ZN(n705) );
  AOI221D0 U390 ( .A1(n692), .A2(n847), .B1(n805), .B2(n691), .C(n690), .ZN(
        n706) );
  ND4D1 U391 ( .A1(n502), .A2(n501), .A3(n500), .A4(n499), .ZN(d[6]) );
  NR4D0 U392 ( .A1(n498), .A2(n497), .A3(n513), .A4(n514), .ZN(n499) );
  AOI221D0 U393 ( .A1(n801), .A2(n833), .B1(n841), .B2(n806), .C(n540), .ZN(
        n573) );
  NR4D0 U394 ( .A1(n569), .A2(n568), .A3(n567), .A4(n730), .ZN(n570) );
  ND4D1 U395 ( .A1(n473), .A2(n474), .A3(n472), .A4(n471), .ZN(d[7]) );
  OAI22D0 U396 ( .A1(n437), .A2(n602), .B1(n433), .B2(n601), .ZN(n603) );
  OAI222D0 U397 ( .A1(n627), .A2(n789), .B1(n601), .B2(n594), .C1(n437), .C2(
        n712), .ZN(n599) );
  AOI21D1 U398 ( .A1(n437), .A2(n848), .B(n807), .ZN(n761) );
  OAI222D0 U399 ( .A1(n748), .A2(n617), .B1(n437), .B2(n616), .C1(n742), .C2(
        n759), .ZN(n620) );
  ND2D1 U400 ( .A1(n435), .A2(n427), .ZN(n738) );
  ND2D0 U401 ( .A1(n428), .A2(n427), .ZN(n695) );
  AOI31D1 U402 ( .A1(n427), .A2(n816), .A3(n787), .B(n815), .ZN(n488) );
  ND2D0 U403 ( .A1(n427), .A2(n808), .ZN(n617) );
  ND2D1 U404 ( .A1(n427), .A2(n729), .ZN(n727) );
  ND2D1 U405 ( .A1(n427), .A2(a[5]), .ZN(n736) );
  AOI22D0 U406 ( .A1(n814), .A2(n786), .B1(n812), .B2(n427), .ZN(n564) );
  AOI21D0 U407 ( .A1(n721), .A2(n661), .B(n427), .ZN(n619) );
  OAI222D0 U408 ( .A1(n633), .A2(n714), .B1(n582), .B2(n722), .C1(n627), .C2(
        n656), .ZN(n475) );
  OAI221D0 U409 ( .A1(n444), .A2(n633), .B1(n763), .B2(n722), .C(n443), .ZN(
        n450) );
  OAI222D0 U410 ( .A1(n737), .A2(n548), .B1(n633), .B2(n710), .C1(n738), .C2(
        n677), .ZN(n447) );
  OAI33D0 U411 ( .A1(n633), .A2(n429), .A3(n760), .B1(n694), .B2(n789), .B3(
        n741), .ZN(n529) );
  OAI222D0 U412 ( .A1(n754), .A2(n753), .B1(n752), .B2(n751), .C1(n434), .C2(
        n750), .ZN(n779) );
  OAI222D0 U413 ( .A1(n751), .A2(n759), .B1(n773), .B2(n637), .C1(n740), .C2(
        n697), .ZN(n645) );
  OA222D0 U414 ( .A1(n738), .A2(n737), .B1(n736), .B2(n735), .C1(n740), .C2(
        n734), .Z(n749) );
  OAI31D1 U415 ( .A1(n738), .A2(n767), .A3(n740), .B(n604), .ZN(n611) );
  INVD1 U416 ( .I(n695), .ZN(n814) );
  NR2D1 U417 ( .A1(n617), .A2(n710), .ZN(n692) );
  OAI211D1 U418 ( .A1(a[5]), .A2(n773), .B(n617), .C(n740), .ZN(n530) );
  INVD1 U419 ( .I(n727), .ZN(n800) );
  AOI31D1 U420 ( .A1(n837), .A2(n727), .A3(n812), .B(n726), .ZN(n728) );
  OAI222D0 U421 ( .A1(n566), .A2(n765), .B1(n774), .B2(n565), .C1(n564), .C2(
        n767), .ZN(n569) );
  INVD1 U422 ( .I(n766), .ZN(n804) );
  NR3D0 U423 ( .A1(n766), .A2(n429), .A3(n428), .ZN(n659) );
  OAI222D0 U424 ( .A1(n774), .A2(n574), .B1(n766), .B2(n628), .C1(n489), .C2(
        n754), .ZN(n490) );
  OAI221D0 U425 ( .A1(n452), .A2(n766), .B1(n712), .B2(n763), .C(n557), .ZN(
        n459) );
  OAI222D0 U426 ( .A1(n767), .A2(n776), .B1(n766), .B2(n765), .C1(n764), .C2(
        n763), .ZN(n768) );
  NR4D0 U427 ( .A1(n760), .A2(n748), .A3(n656), .A4(n437), .ZN(n730) );
  INR2D1 U428 ( .A1(n515), .B1(n656), .ZN(n702) );
  IND4D1 U429 ( .A1(n784), .B1(n783), .B2(n782), .B3(n781), .ZN(d[0]) );
  CKND2D0 U430 ( .A1(n431), .A2(n789), .ZN(n425) );
  CKND2D0 U431 ( .A1(n710), .A2(n438), .ZN(n565) );
  CKND2D0 U432 ( .A1(n786), .A2(n438), .ZN(n713) );
  AOI33D0 U433 ( .A1(n603), .A2(n823), .A3(n792), .B1(n843), .B2(n438), .B3(
        n788), .ZN(n604) );
  CKND2D1 U434 ( .A1(n427), .A2(n438), .ZN(n766) );
  OAI21D0 U435 ( .A1(n633), .A2(n721), .B(n775), .ZN(n465) );
  OAI22D0 U436 ( .A1(n633), .A2(n734), .B1(n735), .B2(n763), .ZN(n492) );
  INVD1 U437 ( .I(n729), .ZN(n788) );
  INVD1 U438 ( .I(n746), .ZN(n810) );
  AOI22D0 U439 ( .A1(n841), .A2(n518), .B1(n684), .B2(n517), .ZN(n519) );
  AOI221D0 U440 ( .A1(n793), .A2(n822), .B1(n817), .B2(n549), .C(n692), .ZN(
        n556) );
  OAI31D0 U441 ( .A1(n438), .A2(n793), .A3(n799), .B(n684), .ZN(n484) );
  OAI32D1 U442 ( .A1(n576), .A2(n735), .A3(n677), .B1(n575), .B2(n756), .ZN(
        n577) );
  AOI21D0 U443 ( .A1(n677), .A2(n756), .B(n424), .ZN(n672) );
  NR3D0 U444 ( .A1(n816), .A2(n435), .A3(n425), .ZN(n524) );
  OAI22D0 U445 ( .A1(n448), .A2(n771), .B1(n738), .B2(n626), .ZN(n449) );
  AOI21D0 U446 ( .A1(n766), .A2(n736), .B(n771), .ZN(n618) );
  NR4D0 U447 ( .A1(n677), .A2(n743), .A3(n771), .A4(n808), .ZN(n648) );
endmodule


module aes_sbox_1 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n51, n65, n68, n70, n71, n72, n123, n142, n148, n187, n192, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863;

  AN2XD1 U28 ( .A1(n725), .A2(n430), .Z(n729) );
  OA21D1 U35 ( .A1(n710), .A2(n709), .B(n708), .Z(n715) );
  OR4D1 U199 ( .A1(n664), .A2(n582), .A3(n526), .A4(n525), .Z(n528) );
  MAOI22D1 U209 ( .A1(n857), .A2(n451), .B1(n633), .B2(n777), .ZN(n519) );
  AN2XD1 U215 ( .A1(n527), .A2(n810), .Z(n526) );
  AN2XD1 U271 ( .A1(n540), .A2(n736), .Z(n473) );
  AO21D1 U297 ( .A1(n123), .A2(n835), .B(n739), .Z(n465) );
  OAI222D1 U1 ( .A1(n432), .A2(n753), .B1(n696), .B2(n692), .C1(n759), .C2(
        n560), .ZN(n538) );
  CKND2 U2 ( .I(a[1]), .ZN(n448) );
  OAI222D1 U3 ( .A1(n787), .A2(n589), .B1(n779), .B2(n644), .C1(n501), .C2(
        n767), .ZN(n502) );
  AOI21D2 U4 ( .A1(n814), .A2(n447), .B(n804), .ZN(n590) );
  ND4D2 U5 ( .A1(n723), .A2(n722), .A3(n721), .A4(n720), .ZN(d[1]) );
  OAI222D1 U6 ( .A1(n469), .A2(n753), .B1(n692), .B2(n520), .C1(n468), .C2(
        n445), .ZN(n470) );
  AOI211XD1 U7 ( .A1(n829), .A2(n594), .B(n593), .C(n592), .ZN(n595) );
  AOI222D1 U8 ( .A1(n808), .A2(n830), .B1(n806), .B2(n489), .C1(n802), .C2(
        n833), .ZN(n494) );
  AOI211D1 U9 ( .A1(n859), .A2(n499), .B(n498), .C(n497), .ZN(n513) );
  INVD2 U10 ( .I(n750), .ZN(n829) );
  INR4D2 U11 ( .A1(n677), .B1(n676), .B2(n675), .B3(n855), .ZN(n686) );
  INVD2 U12 ( .I(n563), .ZN(n802) );
  OAI32D1 U13 ( .A1(n591), .A2(n748), .A3(n692), .B1(n590), .B2(n769), .ZN(
        n592) );
  NR3D1 U14 ( .A1(n434), .A2(n435), .A3(n569), .ZN(n587) );
  OAI222D1 U15 ( .A1(n568), .A2(n761), .B1(n567), .B2(n691), .C1(n566), .C2(
        n755), .ZN(n569) );
  INVD4 U16 ( .I(a[0]), .ZN(n444) );
  INVD2 U17 ( .I(n769), .ZN(n832) );
  OAI222D1 U18 ( .A1(n756), .A2(n613), .B1(n612), .B2(n800), .C1(n611), .C2(
        n683), .ZN(n614) );
  AOI211XD0 U19 ( .A1(n818), .A2(n443), .B(n816), .C(n810), .ZN(n611) );
  CKND4 U20 ( .I(n142), .ZN(n430) );
  AOI21D2 U21 ( .A1(n861), .A2(n816), .B(n855), .ZN(n573) );
  INVD1 U22 ( .I(n431), .ZN(n51) );
  INVD1 U23 ( .I(n51), .ZN(n65) );
  INVD2 U24 ( .I(n51), .ZN(n68) );
  ND3D2 U25 ( .A1(n187), .A2(n192), .A3(n846), .ZN(n676) );
  INVD1 U26 ( .I(n618), .ZN(n70) );
  CKND2 U27 ( .I(n70), .ZN(n71) );
  AOI221D1 U29 ( .A1(n801), .A2(n858), .B1(n810), .B2(n837), .C(n465), .ZN(
        n469) );
  ND2D1 U30 ( .A1(n440), .A2(n819), .ZN(n769) );
  ND2D2 U31 ( .A1(n819), .A2(n827), .ZN(n773) );
  CKND2D0 U32 ( .A1(n800), .A2(n819), .ZN(n559) );
  NR2D0 U33 ( .A1(n819), .A2(n827), .ZN(n678) );
  INVD6 U34 ( .I(n439), .ZN(n819) );
  OAI21D1 U36 ( .A1(n755), .A2(n71), .B(n726), .ZN(n599) );
  INVD2 U37 ( .I(n71), .ZN(n830) );
  ND2D0 U38 ( .A1(n439), .A2(n827), .ZN(n618) );
  CKND2D0 U39 ( .A1(a[3]), .A2(n449), .ZN(n684) );
  CKND2D1 U40 ( .A1(a[3]), .A2(n827), .ZN(n750) );
  CKND6 U41 ( .I(n444), .ZN(n442) );
  INVD3 U42 ( .I(n444), .ZN(n443) );
  CKND2D1 U43 ( .A1(n443), .A2(n438), .ZN(n764) );
  ND2D2 U44 ( .A1(a[1]), .A2(n800), .ZN(n789) );
  AOI221D0 U45 ( .A1(n806), .A2(n543), .B1(n845), .B2(n542), .C(n541), .ZN(
        n544) );
  ND2D1 U46 ( .A1(n803), .A2(n445), .ZN(n560) );
  BUFFD6 U47 ( .I(a[5]), .Z(n440) );
  INVD1 U48 ( .I(a[6]), .ZN(n834) );
  CKND2D1 U49 ( .A1(a[3]), .A2(n819), .ZN(n753) );
  INVD1 U50 ( .I(n772), .ZN(n833) );
  ND2D2 U51 ( .A1(n441), .A2(a[6]), .ZN(n711) );
  BUFFD6 U52 ( .I(a[4]), .Z(n439) );
  ND2D1 U53 ( .A1(n688), .A2(n845), .ZN(n734) );
  INVD3 U54 ( .I(n442), .ZN(n445) );
  INVD1 U55 ( .I(n776), .ZN(n812) );
  ND2D1 U56 ( .A1(n827), .A2(n834), .ZN(n663) );
  OAI31D1 U57 ( .A1(n679), .A2(n72), .A3(n818), .B(n678), .ZN(n680) );
  INVD1 U58 ( .I(n691), .ZN(n814) );
  ND2D1 U59 ( .A1(n428), .A2(n429), .ZN(n671) );
  OAI222D0 U60 ( .A1(n811), .A2(n638), .B1(n560), .B2(n540), .C1(n539), .C2(
        n784), .ZN(n546) );
  AOI221D0 U61 ( .A1(n835), .A2(n142), .B1(n599), .B2(n448), .C(n739), .ZN(
        n600) );
  AN2XD1 U62 ( .A1(n859), .A2(n652), .Z(n424) );
  OAI221D0 U63 ( .A1(n743), .A2(n691), .B1(n750), .B2(n710), .C(n690), .ZN(
        n698) );
  AOI221D0 U64 ( .A1(n799), .A2(n694), .B1(n833), .B2(n72), .C(n693), .ZN(n695) );
  ND2D1 U65 ( .A1(n842), .A2(n828), .ZN(n726) );
  OAI222D0 U66 ( .A1(n762), .A2(n761), .B1(n760), .B2(n759), .C1(n443), .C2(
        n758), .ZN(n793) );
  ND2D1 U67 ( .A1(n439), .A2(n450), .ZN(n716) );
  AOI22D1 U68 ( .A1(n812), .A2(n832), .B1(n814), .B2(n827), .ZN(n768) );
  AN2XD1 U69 ( .A1(n443), .A2(n800), .Z(n72) );
  ND2D1 U70 ( .A1(n449), .A2(n800), .ZN(n756) );
  INVD2 U71 ( .I(a[3]), .ZN(n450) );
  INVD1 U72 ( .I(n72), .ZN(n432) );
  AN2XD1 U73 ( .A1(n443), .A2(n448), .Z(n123) );
  AN2XD1 U74 ( .A1(a[1]), .A2(n442), .Z(n142) );
  AN3XD1 U75 ( .A1(n586), .A2(n588), .A3(n585), .Z(n148) );
  INVD2 U76 ( .I(n438), .ZN(n800) );
  ND2D1 U77 ( .A1(n438), .A2(n450), .ZN(n779) );
  ND2D0 U78 ( .A1(n678), .A2(n848), .ZN(n596) );
  OAI22D1 U79 ( .A1(n460), .A2(n784), .B1(n751), .B2(n642), .ZN(n461) );
  ND2D1 U80 ( .A1(n808), .A2(n445), .ZN(n712) );
  NR4D0 U81 ( .A1(n791), .A2(n792), .A3(n793), .A4(n790), .ZN(n794) );
  ND2D1 U82 ( .A1(n439), .A2(a[3]), .ZN(n754) );
  OAI222D1 U83 ( .A1(n672), .A2(n772), .B1(n442), .B2(n564), .C1(n754), .C2(
        n563), .ZN(n565) );
  ND2D0 U84 ( .A1(n754), .A2(n749), .ZN(n556) );
  OAI222D1 U85 ( .A1(n432), .A2(n540), .B1(n494), .B2(n755), .C1(n493), .C2(
        n759), .ZN(n498) );
  AOI221D1 U86 ( .A1(n467), .A2(n808), .B1(n852), .B2(n817), .C(n466), .ZN(
        n468) );
  OAI222D1 U87 ( .A1(n575), .A2(n716), .B1(n574), .B2(n68), .C1(n447), .C2(
        n573), .ZN(n576) );
  OAI222D1 U88 ( .A1(n650), .A2(n649), .B1(n764), .B2(n766), .C1(n648), .C2(
        n776), .ZN(n651) );
  CKND2D1 U89 ( .A1(a[3]), .A2(n440), .ZN(n692) );
  AOI221D1 U90 ( .A1(n847), .A2(n445), .B1(n857), .B2(n447), .C(n647), .ZN(
        n648) );
  ND2D0 U91 ( .A1(n447), .A2(n438), .ZN(n751) );
  AOI22D1 U92 ( .A1(n809), .A2(n858), .B1(n801), .B2(n837), .ZN(n575) );
  ND2D1 U93 ( .A1(n845), .A2(n832), .ZN(n787) );
  AOI221D1 U94 ( .A1(n845), .A2(n463), .B1(n462), .B2(n445), .C(n461), .ZN(
        n486) );
  AOI221D1 U95 ( .A1(n845), .A2(n616), .B1(n615), .B2(n445), .C(n614), .ZN(
        n629) );
  INVD2 U96 ( .I(n755), .ZN(n845) );
  INVD4 U97 ( .I(n784), .ZN(n842) );
  ND2D2 U98 ( .A1(a[6]), .A2(n839), .ZN(n784) );
  AOI22D1 U99 ( .A1(n838), .A2(n806), .B1(n809), .B2(n837), .ZN(n474) );
  OAI22D1 U100 ( .A1(n474), .A2(n716), .B1(n473), .B2(n764), .ZN(n475) );
  CKND2D2 U101 ( .A1(n834), .A2(n839), .ZN(n755) );
  CKND1 U102 ( .I(n716), .ZN(n824) );
  ND2D2 U103 ( .A1(a[3]), .A2(n800), .ZN(n776) );
  AOI221D1 U104 ( .A1(n123), .A2(n689), .B1(n688), .B2(n806), .C(n687), .ZN(
        n690) );
  ND2D1 U105 ( .A1(n441), .A2(n827), .ZN(n732) );
  OA221D1 U106 ( .A1(n750), .A2(n743), .B1(n759), .B2(n672), .C(n433), .Z(n685) );
  ND2D1 U107 ( .A1(n800), .A2(n450), .ZN(n691) );
  OA21D0 U108 ( .A1(n691), .A2(n446), .B(n621), .Z(n625) );
  ND2D1 U109 ( .A1(n440), .A2(n450), .ZN(n772) );
  AOI21D1 U110 ( .A1(n833), .A2(n842), .B(n851), .ZN(n673) );
  AO221D1 U111 ( .A1(n801), .A2(n833), .B1(n799), .B2(n815), .C(n707), .Z(n660) );
  INVD4 U112 ( .I(n441), .ZN(n839) );
  ND2D1 U113 ( .A1(n852), .A2(n445), .ZN(n644) );
  AOI221D1 U114 ( .A1(n836), .A2(n824), .B1(n822), .B2(n578), .C(n851), .ZN(
        n501) );
  NR4D1 U115 ( .A1(n548), .A2(n547), .A3(n546), .A4(n545), .ZN(n549) );
  OAI222D1 U116 ( .A1(n535), .A2(n779), .B1(n432), .B2(n632), .C1(n534), .C2(
        n430), .ZN(n547) );
  OAI33D0 U117 ( .A1(n756), .A2(n755), .A3(n754), .B1(n777), .B2(n800), .B3(
        n753), .ZN(n757) );
  OA222D0 U118 ( .A1(n751), .A2(n750), .B1(n749), .B2(n748), .C1(n753), .C2(
        n65), .Z(n762) );
  AOI221D1 U119 ( .A1(n860), .A2(n445), .B1(n852), .B2(n808), .C(n639), .ZN(
        n670) );
  AOI221D1 U120 ( .A1(n699), .A2(n748), .B1(n447), .B2(n854), .C(n562), .ZN(
        n567) );
  INVD1 U121 ( .I(n761), .ZN(n859) );
  ND2D2 U122 ( .A1(n441), .A2(n834), .ZN(n761) );
  AOI221D1 U123 ( .A1(n856), .A2(n142), .B1(n859), .B2(n698), .C(n697), .ZN(
        n722) );
  INVD1 U124 ( .I(n560), .ZN(n804) );
  OAI222D1 U125 ( .A1(n649), .A2(n642), .B1(n597), .B2(n596), .C1(n761), .C2(
        n595), .ZN(n598) );
  OA221D1 U126 ( .A1(n638), .A2(n764), .B1(n436), .B2(n789), .C(n437), .Z(n723) );
  INVD6 U127 ( .I(n440), .ZN(n827) );
  OAI221D1 U128 ( .A1(n617), .A2(n591), .B1(a[3]), .B2(n778), .C(n708), .ZN(
        n533) );
  AOI22D1 U129 ( .A1(n830), .A2(n816), .B1(n806), .B2(n827), .ZN(n564) );
  INVD1 U130 ( .I(n649), .ZN(n816) );
  ND2D2 U131 ( .A1(n801), .A2(n442), .ZN(n563) );
  AOI221D1 U132 ( .A1(n822), .A2(n798), .B1(n831), .B2(n808), .C(n565), .ZN(
        n566) );
  ND2D1 U133 ( .A1(a[3]), .A2(n438), .ZN(n649) );
  OAI222D1 U134 ( .A1(n749), .A2(n430), .B1(n773), .B2(n589), .C1(n754), .C2(
        n764), .ZN(n593) );
  NR2D0 U135 ( .A1(n832), .A2(n812), .ZN(n521) );
  CKND2D1 U136 ( .A1(n832), .A2(n839), .ZN(n632) );
  ND2D2 U137 ( .A1(n848), .A2(n832), .ZN(n643) );
  AOI221D1 U138 ( .A1(n801), .A2(n824), .B1(n809), .B2(n831), .C(n770), .ZN(
        n785) );
  OA221D1 U139 ( .A1(n691), .A2(n682), .B1(n681), .B2(n789), .C(n680), .Z(n433) );
  INVD2 U140 ( .I(n711), .ZN(n848) );
  ND2D0 U141 ( .A1(n445), .A2(n800), .ZN(n767) );
  AOI221D1 U142 ( .A1(n707), .A2(n858), .B1(n816), .B2(n706), .C(n705), .ZN(
        n721) );
  ND3D0 U143 ( .A1(n816), .A2(n678), .A3(n845), .ZN(n763) );
  CKND2D1 U144 ( .A1(n438), .A2(n440), .ZN(n749) );
  CKND2D0 U145 ( .A1(n440), .A2(n834), .ZN(n515) );
  CKND2D1 U146 ( .A1(n440), .A2(n441), .ZN(n709) );
  CKND2D1 U147 ( .A1(n842), .A2(n678), .ZN(n736) );
  ND2D0 U148 ( .A1(n827), .A2(n839), .ZN(n617) );
  CKND2D1 U149 ( .A1(n678), .A2(n859), .ZN(n778) );
  CKND2D1 U150 ( .A1(n440), .A2(n839), .ZN(n713) );
  ND2D0 U151 ( .A1(a[6]), .A2(n827), .ZN(n777) );
  AOI221D1 U152 ( .A1(n813), .A2(n578), .B1(n577), .B2(n822), .C(n576), .ZN(
        n586) );
  AOI221D1 U153 ( .A1(n842), .A2(n503), .B1(n802), .B2(n516), .C(n502), .ZN(
        n512) );
  OAI33D0 U154 ( .A1(n663), .A2(n443), .A3(n800), .B1(n490), .B2(n732), .B3(
        n764), .ZN(n491) );
  CKND1 U155 ( .I(n732), .ZN(n858) );
  BUFFD8 U156 ( .I(a[2]), .Z(n438) );
  AOI221D1 U157 ( .A1(n815), .A2(n608), .B1(n842), .B2(n607), .C(n606), .ZN(
        n630) );
  OAI222D1 U158 ( .A1(n785), .A2(n784), .B1(a[3]), .B2(n840), .C1(n783), .C2(
        n445), .ZN(n791) );
  NR2XD0 U159 ( .A1(n812), .A2(n805), .ZN(n453) );
  OAI211D0 U160 ( .A1(n827), .A2(n759), .B(n776), .C(n754), .ZN(n689) );
  OR2D0 U161 ( .A1(n674), .A2(n684), .Z(n187) );
  OR2D0 U162 ( .A1(n673), .A2(n672), .Z(n192) );
  NR2D0 U163 ( .A1(n843), .A2(n854), .ZN(n674) );
  INVD1 U164 ( .I(n671), .ZN(n846) );
  CKAN2D1 U165 ( .A1(n856), .A2(n803), .Z(n425) );
  NR3D1 U166 ( .A1(n424), .A2(n425), .A3(n651), .ZN(n669) );
  INVD2 U167 ( .I(n789), .ZN(n803) );
  CKAN2D1 U168 ( .A1(n447), .A2(n471), .Z(n426) );
  CKAN2D1 U169 ( .A1(n826), .A2(n836), .Z(n427) );
  NR3D0 U170 ( .A1(n426), .A2(n427), .A3(n470), .ZN(n485) );
  INVD2 U171 ( .I(n448), .ZN(n447) );
  OR2XD1 U172 ( .A1(n728), .A2(n756), .Z(n428) );
  OR2D0 U173 ( .A1(n800), .A2(n734), .Z(n429) );
  AOI211XD0 U174 ( .A1(n863), .A2(n809), .B(n487), .C(n671), .ZN(n514) );
  OAI33D0 U175 ( .A1(n759), .A2(n800), .A3(n732), .B1(n663), .B2(n447), .B3(
        n662), .ZN(n666) );
  CKND2D0 U176 ( .A1(n815), .A2(n447), .ZN(n725) );
  AOI21D0 U177 ( .A1(n856), .A2(n447), .B(n699), .ZN(n700) );
  OAI31D0 U178 ( .A1(n711), .A2(n440), .A3(n447), .B(n644), .ZN(n562) );
  OAI22D0 U179 ( .A1(n769), .A2(n779), .B1(n447), .B2(n768), .ZN(n770) );
  ND2D0 U180 ( .A1(n812), .A2(n447), .ZN(n589) );
  ND2D0 U181 ( .A1(n447), .A2(a[3]), .ZN(n786) );
  AOI221D1 U182 ( .A1(n802), .A2(n850), .B1(n142), .B2(n863), .C(n598), .ZN(
        n631) );
  CKND0 U183 ( .I(n123), .ZN(n431) );
  OAI33D0 U184 ( .A1(n649), .A2(n441), .A3(n773), .B1(n709), .B2(n800), .B3(
        n754), .ZN(n541) );
  OAI22D0 U185 ( .A1(n649), .A2(n68), .B1(n748), .B2(n776), .ZN(n504) );
  NR2XD0 U186 ( .A1(n798), .A2(n806), .ZN(n657) );
  CKND2D0 U187 ( .A1(n72), .A2(n832), .ZN(n653) );
  CKND2D0 U188 ( .A1(n822), .A2(n848), .ZN(n613) );
  CKND2D1 U189 ( .A1(n830), .A2(n848), .ZN(n735) );
  CKND2D0 U190 ( .A1(n828), .A2(n848), .ZN(n642) );
  ND2D0 U191 ( .A1(n830), .A2(n859), .ZN(n683) );
  BUFFD4 U192 ( .I(a[7]), .Z(n441) );
  CKND2D0 U193 ( .A1(n786), .A2(n691), .ZN(n529) );
  NR2D0 U194 ( .A1(n632), .A2(n68), .ZN(n771) );
  NR2D0 U195 ( .A1(n808), .A2(n142), .ZN(n621) );
  NR2D0 U196 ( .A1(n643), .A2(n727), .ZN(n745) );
  CKND2D0 U197 ( .A1(n799), .A2(n859), .ZN(n520) );
  CKND2D0 U198 ( .A1(n496), .A2(n495), .ZN(n497) );
  CKND2D0 U200 ( .A1(n692), .A2(n753), .ZN(n694) );
  NR2D1 U201 ( .A1(n713), .A2(n716), .ZN(n724) );
  CKND2D0 U202 ( .A1(n767), .A2(n764), .ZN(n752) );
  CKND2D0 U203 ( .A1(n688), .A2(n848), .ZN(n638) );
  ND2D0 U204 ( .A1(n830), .A2(n448), .ZN(n682) );
  AOI211XD0 U205 ( .A1(n843), .A2(n443), .B(n645), .C(n853), .ZN(n650) );
  NR2D0 U206 ( .A1(n810), .A2(n808), .ZN(n472) );
  AOI211XD0 U207 ( .A1(n841), .A2(n809), .B(n492), .C(n491), .ZN(n493) );
  CKND2D1 U208 ( .A1(n777), .A2(n732), .ZN(n578) );
  CKND2D0 U210 ( .A1(n447), .A2(a[6]), .ZN(n490) );
  NR2D0 U211 ( .A1(n446), .A2(n763), .ZN(n746) );
  NR2D0 U212 ( .A1(n805), .A2(n801), .ZN(n479) );
  CKND2D0 U213 ( .A1(n733), .A2(n743), .ZN(n594) );
  NR2D0 U214 ( .A1(n72), .A2(n798), .ZN(n622) );
  ND2D0 U216 ( .A1(n812), .A2(n854), .ZN(n572) );
  CKND0 U217 ( .I(n778), .ZN(n860) );
  CKND0 U218 ( .I(n589), .ZN(n813) );
  OAI22D0 U219 ( .A1(n759), .A2(n756), .B1(n662), .B2(n743), .ZN(n524) );
  OAI22D0 U220 ( .A1(n68), .A2(n759), .B1(n609), .B2(n748), .ZN(n616) );
  NR2D0 U221 ( .A1(n825), .A2(n830), .ZN(n609) );
  NR2D0 U222 ( .A1(n816), .A2(n823), .ZN(n662) );
  AOI22D0 U223 ( .A1(n852), .A2(n530), .B1(n699), .B2(n529), .ZN(n531) );
  CKND2D0 U224 ( .A1(n862), .A2(n824), .ZN(n788) );
  ND2D0 U225 ( .A1(n822), .A2(n862), .ZN(n765) );
  CKND2D0 U226 ( .A1(n821), .A2(n845), .ZN(n677) );
  CKND2D0 U227 ( .A1(n835), .A2(n824), .ZN(n540) );
  NR2D0 U228 ( .A1(n857), .A2(n699), .ZN(n456) );
  NR2D0 U229 ( .A1(n724), .A2(n857), .ZN(n730) );
  NR2D0 U230 ( .A1(n861), .A2(n847), .ZN(n464) );
  OAI22D0 U231 ( .A1(n769), .A2(n691), .B1(n696), .B2(n716), .ZN(n458) );
  AOI21D0 U232 ( .A1(n691), .A2(n591), .B(n65), .ZN(n457) );
  ND2D0 U233 ( .A1(n816), .A2(n819), .ZN(n610) );
  NR2XD0 U234 ( .A1(n837), .A2(n848), .ZN(n646) );
  OAI22D0 U235 ( .A1(n750), .A2(n756), .B1(n769), .B2(n789), .ZN(n693) );
  OAI22D0 U236 ( .A1(n445), .A2(n726), .B1(n449), .B2(n736), .ZN(n532) );
  NR2D0 U237 ( .A1(n755), .A2(n773), .ZN(n699) );
  CKND2D1 U238 ( .A1(n445), .A2(n448), .ZN(n748) );
  OAI32D0 U239 ( .A1(n563), .A2(n761), .A3(n750), .B1(n521), .B2(n520), .ZN(
        n522) );
  OAI22D0 U240 ( .A1(n789), .A2(n788), .B1(n787), .B2(n786), .ZN(n790) );
  OAI31D0 U241 ( .A1(n743), .A2(n823), .A3(n755), .B(n742), .ZN(n747) );
  AOI31D0 U242 ( .A1(n848), .A2(n741), .A3(n823), .B(n740), .ZN(n742) );
  OAI31D0 U243 ( .A1(n450), .A2(n804), .A3(n810), .B(n699), .ZN(n496) );
  OAI21D0 U244 ( .A1(n754), .A2(n617), .B(n642), .ZN(n516) );
  AOI22D0 U245 ( .A1(n445), .A2(n817), .B1(n451), .B2(n805), .ZN(n597) );
  NR2D0 U246 ( .A1(n633), .A2(n430), .ZN(n707) );
  AOI22D0 U247 ( .A1(n808), .A2(n442), .B1(n447), .B2(n816), .ZN(n488) );
  AOI21D0 U248 ( .A1(n71), .A2(n663), .B(n691), .ZN(n505) );
  INR2D0 U249 ( .A1(n527), .B1(n672), .ZN(n717) );
  AOI22D0 U250 ( .A1(n836), .A2(n752), .B1(n838), .B2(n806), .ZN(n760) );
  AOI21D0 U251 ( .A1(n692), .A2(n769), .B(n432), .ZN(n687) );
  OAI21D0 U252 ( .A1(n442), .A2(n692), .B(n753), .ZN(n489) );
  CKND0 U253 ( .I(n709), .ZN(n862) );
  CKND2D0 U254 ( .A1(n798), .A2(n450), .ZN(n727) );
  OAI21D0 U255 ( .A1(n649), .A2(n735), .B(n788), .ZN(n477) );
  CKND2D0 U256 ( .A1(n831), .A2(n848), .ZN(n766) );
  OAI22D0 U257 ( .A1(n449), .A2(n726), .B1(n447), .B2(n643), .ZN(n645) );
  AOI32D0 U258 ( .A1(n801), .A2(n445), .A3(n833), .B1(n799), .B2(n556), .ZN(
        n558) );
  AOI31D0 U259 ( .A1(n736), .A2(n735), .A3(n734), .B(n733), .ZN(n737) );
  AOI32D0 U260 ( .A1(n440), .A2(n445), .A3(n817), .B1(n828), .B2(n640), .ZN(
        n641) );
  CKND2D1 U261 ( .A1(n603), .A2(n602), .ZN(n607) );
  AOI21D0 U262 ( .A1(n807), .A2(n845), .B(n577), .ZN(n518) );
  CKND0 U263 ( .I(n617), .ZN(n841) );
  NR2D0 U264 ( .A1(n810), .A2(a[3]), .ZN(n624) );
  AOI21D0 U265 ( .A1(n822), .A2(n858), .B(n701), .ZN(n508) );
  INR2XD0 U266 ( .A1(n765), .B1(n505), .ZN(n506) );
  CKND0 U267 ( .I(n771), .ZN(n840) );
  AOI211D0 U268 ( .A1(n804), .A2(n823), .B(n826), .C(n702), .ZN(n703) );
  AOI21D0 U269 ( .A1(n857), .A2(n817), .B(n701), .ZN(n704) );
  AOI21D0 U270 ( .A1(n847), .A2(n816), .B(n757), .ZN(n758) );
  OAI21D0 U272 ( .A1(n663), .A2(n753), .B(n734), .ZN(n543) );
  OAI211D0 U273 ( .A1(n440), .A2(n786), .B(n633), .C(n753), .ZN(n542) );
  OAI22D0 U274 ( .A1(n449), .A2(n638), .B1(n637), .B2(n68), .ZN(n639) );
  OAI31D0 U275 ( .A1(n751), .A2(n780), .A3(n753), .B(n620), .ZN(n627) );
  AOI33D0 U276 ( .A1(n619), .A2(n834), .A3(n803), .B1(n854), .B2(n450), .B3(
        n799), .ZN(n620) );
  OAI22D0 U277 ( .A1(a[3]), .A2(n71), .B1(n445), .B2(n617), .ZN(n619) );
  AOI211D0 U278 ( .A1(n780), .A2(n663), .B(n591), .C(n68), .ZN(n480) );
  NR2D0 U279 ( .A1(a[3]), .A2(n440), .ZN(n688) );
  AOI21D0 U280 ( .A1(a[3]), .A2(n859), .B(n818), .ZN(n774) );
  NR2D0 U281 ( .A1(n804), .A2(n807), .ZN(n581) );
  CKND2D0 U282 ( .A1(n430), .A2(n450), .ZN(n580) );
  AOI32D0 U283 ( .A1(n441), .A2(n819), .A3(n801), .B1(n806), .B2(n454), .ZN(
        n455) );
  OAI22D0 U284 ( .A1(n441), .A2(n663), .B1(n754), .B2(n732), .ZN(n454) );
  CKND2D0 U285 ( .A1(n438), .A2(n819), .ZN(n633) );
  OAI21D0 U286 ( .A1(n715), .A2(n743), .B(n714), .ZN(n719) );
  CKND2D0 U287 ( .A1(n438), .A2(n743), .ZN(n741) );
  OAI22D0 U288 ( .A1(n834), .A2(n716), .B1(n819), .B2(n663), .ZN(n655) );
  AO31D0 U289 ( .A1(n803), .A2(n859), .A3(n688), .B(n724), .Z(n466) );
  AOI22D0 U290 ( .A1(n861), .A2(n803), .B1(n817), .B2(n847), .ZN(n554) );
  CKND2D0 U291 ( .A1(n440), .A2(a[6]), .ZN(n780) );
  INVD1 U292 ( .I(n572), .ZN(n855) );
  INVD1 U293 ( .I(n786), .ZN(n817) );
  INVD1 U294 ( .I(n787), .ZN(n847) );
  INVD1 U295 ( .I(n683), .ZN(n861) );
  INVD1 U296 ( .I(n712), .ZN(n809) );
  INVD1 U298 ( .I(n605), .ZN(n826) );
  INVD1 U299 ( .I(n733), .ZN(n807) );
  INVD1 U300 ( .I(n788), .ZN(n863) );
  ND2D1 U301 ( .A1(n432), .A2(n756), .ZN(n530) );
  INVD1 U302 ( .I(n753), .ZN(n822) );
  NR2D1 U303 ( .A1(n763), .A2(n443), .ZN(n718) );
  NR2D1 U304 ( .A1(n446), .A2(a[3]), .ZN(n679) );
  NR2D1 U305 ( .A1(n735), .A2(a[3]), .ZN(n701) );
  INVD1 U306 ( .I(n596), .ZN(n857) );
  INVD1 U307 ( .I(n773), .ZN(n828) );
  ND2D1 U308 ( .A1(n447), .A2(n445), .ZN(n743) );
  INVD1 U309 ( .I(n642), .ZN(n856) );
  INVD1 U310 ( .I(n735), .ZN(n852) );
  ND2D1 U311 ( .A1(n443), .A2(n806), .ZN(n733) );
  NR3D0 U312 ( .A1(n679), .A2(n801), .A3(n815), .ZN(n656) );
  INVD1 U313 ( .I(n767), .ZN(n805) );
  INVD1 U314 ( .I(n643), .ZN(n854) );
  ND2D1 U315 ( .A1(n142), .A2(n825), .ZN(n605) );
  INVD1 U316 ( .I(n604), .ZN(n851) );
  INVD1 U317 ( .I(n748), .ZN(n798) );
  INVD1 U318 ( .I(n756), .ZN(n801) );
  INVD1 U319 ( .I(n684), .ZN(n818) );
  ND2D1 U320 ( .A1(n820), .A2(n836), .ZN(n708) );
  INVD1 U321 ( .I(n559), .ZN(n820) );
  INVD1 U322 ( .I(n726), .ZN(n844) );
  INVD1 U323 ( .I(n613), .ZN(n849) );
  INVD1 U324 ( .I(n442), .ZN(n446) );
  NR2D1 U325 ( .A1(n654), .A2(n771), .ZN(n612) );
  AOI221D0 U326 ( .A1(n861), .A2(n448), .B1(n843), .B2(n430), .C(n532), .ZN(
        n535) );
  AOI221D0 U327 ( .A1(n822), .A2(n859), .B1(n812), .B2(n832), .C(n533), .ZN(
        n534) );
  NR4D0 U328 ( .A1(n716), .A2(n767), .A3(n761), .A4(n827), .ZN(n740) );
  AOI21D1 U329 ( .A1(n820), .A2(n862), .B(n849), .ZN(n574) );
  OAI222D0 U330 ( .A1(n756), .A2(n692), .B1(n488), .B2(n769), .C1(n447), .C2(
        n754), .ZN(n499) );
  OAI222D0 U331 ( .A1(n761), .A2(n633), .B1(a[3]), .B2(n632), .C1(n755), .C2(
        n772), .ZN(n636) );
  AOI221D0 U332 ( .A1(n804), .A2(n833), .B1(n828), .B2(n561), .C(n707), .ZN(
        n568) );
  OAI222D0 U333 ( .A1(n432), .A2(n604), .B1(n736), .B2(n684), .C1(n643), .C2(
        n764), .ZN(n552) );
  NR2D1 U334 ( .A1(n709), .A2(n748), .ZN(n739) );
  NR4D0 U335 ( .A1(n773), .A2(n761), .A3(n672), .A4(a[3]), .ZN(n744) );
  OAI221D0 U336 ( .A1(n464), .A2(n779), .B1(n726), .B2(n776), .C(n572), .ZN(
        n471) );
  OAI22D1 U337 ( .A1(n748), .A2(n713), .B1(n646), .B2(n743), .ZN(n647) );
  INVD1 U338 ( .I(n672), .ZN(n806) );
  NR3D0 U339 ( .A1(n827), .A2(a[1]), .A3(n432), .ZN(n536) );
  INVD1 U340 ( .I(n663), .ZN(n836) );
  OAI222D0 U341 ( .A1(n767), .A2(n766), .B1(n765), .B2(n764), .C1(n447), .C2(
        n763), .ZN(n792) );
  NR4D0 U342 ( .A1(n459), .A2(n458), .A3(n536), .A4(n457), .ZN(n460) );
  INVD1 U343 ( .I(n644), .ZN(n853) );
  NR4D0 U344 ( .A1(n538), .A2(n537), .A3(n536), .A4(n601), .ZN(n539) );
  NR3D0 U345 ( .A1(n743), .A2(a[3]), .A3(n769), .ZN(n537) );
  NR3D0 U346 ( .A1(n430), .A2(n819), .A3(n734), .ZN(n582) );
  NR3D0 U347 ( .A1(n515), .A2(n754), .A3(n789), .ZN(n481) );
  INVD1 U348 ( .I(n754), .ZN(n823) );
  INVD1 U349 ( .I(n779), .ZN(n815) );
  ND2D1 U350 ( .A1(n830), .A2(n842), .ZN(n728) );
  INVD1 U351 ( .I(n751), .ZN(n808) );
  INVD1 U352 ( .I(n699), .ZN(n436) );
  ND2D1 U353 ( .A1(n451), .A2(n819), .ZN(n759) );
  INVD1 U354 ( .I(n515), .ZN(n835) );
  INVD1 U355 ( .I(n710), .ZN(n825) );
  ND2D1 U356 ( .A1(n829), .A2(n848), .ZN(n604) );
  INVD1 U357 ( .I(n692), .ZN(n831) );
  OAI222D0 U358 ( .A1(n643), .A2(n800), .B1(n617), .B2(n610), .C1(a[3]), .C2(
        n726), .ZN(n615) );
  AOI221D0 U359 ( .A1(n142), .A2(n814), .B1(n802), .B2(n829), .C(n601), .ZN(
        n602) );
  INVD1 U360 ( .I(n741), .ZN(n811) );
  OAI222D0 U361 ( .A1(n732), .A2(n605), .B1(n432), .B2(n766), .C1(n621), .C2(
        n604), .ZN(n606) );
  OAI221D0 U362 ( .A1(n743), .A2(n736), .B1(n711), .B2(n748), .C(n600), .ZN(
        n608) );
  OAI221D0 U363 ( .A1(n622), .A2(n769), .B1(n754), .B2(n764), .C(n500), .ZN(
        n503) );
  OAI222D0 U364 ( .A1(n735), .A2(n725), .B1(n704), .B2(n445), .C1(n703), .C2(
        n777), .ZN(n705) );
  OAI222D0 U365 ( .A1(n625), .A2(n778), .B1(n624), .B2(n728), .C1(n623), .C2(
        n759), .ZN(n626) );
  OA22D0 U366 ( .A1(n780), .A2(n68), .B1(n732), .B2(n622), .Z(n623) );
  AOI222D0 U367 ( .A1(n803), .A2(n821), .B1(n823), .B2(n805), .C1(n807), .C2(
        n440), .ZN(n603) );
  OAI222D0 U368 ( .A1(n441), .A2(n775), .B1(n774), .B2(n773), .C1(n784), .C2(
        n772), .ZN(n782) );
  AOI221D0 U369 ( .A1(n842), .A2(n661), .B1(n845), .B2(n660), .C(n659), .ZN(
        n668) );
  OAI222D0 U370 ( .A1(n764), .A2(n772), .B1(n786), .B2(n653), .C1(n753), .C2(
        n712), .ZN(n661) );
  OAI222D0 U371 ( .A1(n438), .A2(n658), .B1(n657), .B2(n788), .C1(n656), .C2(
        n787), .ZN(n659) );
  OAI222D0 U372 ( .A1(n447), .A2(n780), .B1(n748), .B2(n761), .C1(n755), .C2(
        n751), .ZN(n492) );
  OAI222D0 U373 ( .A1(n581), .A2(n778), .B1(n787), .B2(n580), .C1(n579), .C2(
        n780), .ZN(n584) );
  OAI221D0 U374 ( .A1(n754), .A2(n756), .B1(n716), .B2(n789), .C(n641), .ZN(
        n652) );
  OAI221D0 U375 ( .A1(n453), .A2(n71), .B1(n779), .B2(n430), .C(n452), .ZN(
        n463) );
  OAI221D0 U376 ( .A1(n456), .A2(n649), .B1(n776), .B2(n736), .C(n455), .ZN(
        n462) );
  OAI222D0 U377 ( .A1(n756), .A2(n765), .B1(n696), .B2(n726), .C1(n695), .C2(
        n784), .ZN(n697) );
  OAI221D0 U378 ( .A1(n447), .A2(n677), .B1(n727), .B2(n683), .C(n531), .ZN(
        n548) );
  OAI222D0 U379 ( .A1(n712), .A2(n736), .B1(n442), .B2(n544), .C1(n789), .C2(
        n778), .ZN(n545) );
  NR4D0 U380 ( .A1(n636), .A2(n635), .A3(n849), .A4(n634), .ZN(n637) );
  AOI221D0 U381 ( .A1(n739), .A2(n815), .B1(n814), .B2(n738), .C(n737), .ZN(
        n796) );
  OAI221D0 U382 ( .A1(n743), .A2(n732), .B1(a[1]), .B2(n787), .C(n731), .ZN(
        n738) );
  OAI221D0 U383 ( .A1(n445), .A2(n736), .B1(n711), .B2(n430), .C(n700), .ZN(
        n706) );
  NR4D0 U384 ( .A1(n443), .A2(n834), .A3(n773), .A4(n779), .ZN(n583) );
  OAI222D0 U385 ( .A1(n519), .A2(n68), .B1(n518), .B2(n754), .C1(n517), .C2(
        n767), .ZN(n523) );
  NR2D1 U386 ( .A1(n860), .A2(n516), .ZN(n517) );
  INVD1 U387 ( .I(n777), .ZN(n837) );
  AOI21D1 U388 ( .A1(n142), .A2(n655), .B(n654), .ZN(n658) );
  OAI222D0 U389 ( .A1(n508), .A2(n748), .B1(n819), .B2(n507), .C1(n506), .C2(
        n430), .ZN(n510) );
  ND2D1 U390 ( .A1(n441), .A2(n504), .ZN(n507) );
  INVD1 U391 ( .I(n780), .ZN(n838) );
  OAI222D0 U392 ( .A1(n479), .A2(n713), .B1(n472), .B2(n711), .C1(n732), .C2(
        n733), .ZN(n476) );
  OAI222D0 U393 ( .A1(n780), .A2(n789), .B1(n779), .B2(n778), .C1(n777), .C2(
        n776), .ZN(n781) );
  INVD1 U394 ( .I(a[1]), .ZN(n449) );
  INVD1 U395 ( .I(a[3]), .ZN(n451) );
  ND4D1 U396 ( .A1(n514), .A2(n513), .A3(n512), .A4(n511), .ZN(d[6]) );
  NR4D0 U397 ( .A1(n510), .A2(n509), .A3(n525), .A4(n526), .ZN(n511) );
  NR4D0 U398 ( .A1(n747), .A2(n746), .A3(n745), .A4(n744), .ZN(n795) );
  OAI222D0 U399 ( .A1(n730), .A2(n432), .B1(n729), .B2(n728), .C1(n727), .C2(
        n726), .ZN(n797) );
  ND3D1 U400 ( .A1(n551), .A2(n550), .A3(n549), .ZN(d[5]) );
  INR4D0 U401 ( .A1(n763), .B1(n528), .B2(n745), .B3(n717), .ZN(n550) );
  AOI211D1 U402 ( .A1(n862), .A2(n524), .B(n523), .C(n522), .ZN(n551) );
  ND4D1 U403 ( .A1(n670), .A2(n669), .A3(n668), .A4(n667), .ZN(d[2]) );
  NR4D0 U404 ( .A1(n666), .A2(n665), .A3(n664), .A4(n746), .ZN(n667) );
  ND4D1 U405 ( .A1(n484), .A2(n485), .A3(n486), .A4(n483), .ZN(d[7]) );
  NR4D0 U406 ( .A1(n482), .A2(n481), .A3(n718), .A4(n480), .ZN(n483) );
  AOI221D0 U407 ( .A1(n477), .A2(n448), .B1(n821), .B2(n476), .C(n475), .ZN(
        n484) );
  NR4D0 U408 ( .A1(n719), .A2(n740), .A3(n718), .A4(n717), .ZN(n720) );
  ND4D1 U409 ( .A1(n631), .A2(n630), .A3(n629), .A4(n628), .ZN(d[3]) );
  NR2D1 U410 ( .A1(n627), .A2(n626), .ZN(n628) );
  INVD1 U411 ( .I(n743), .ZN(n799) );
  INVD1 U412 ( .I(n759), .ZN(n821) );
  OAI222D0 U413 ( .A1(n649), .A2(n728), .B1(n597), .B2(n736), .C1(n643), .C2(
        n672), .ZN(n487) );
  ND4D1 U414 ( .A1(n123), .A2(n836), .A3(n439), .A4(n441), .ZN(n731) );
  AN4D1 U415 ( .A1(n678), .A2(n817), .A3(n443), .A4(n845), .Z(n525) );
  NR3D0 U416 ( .A1(n779), .A2(n441), .A3(n439), .ZN(n675) );
  NR3D0 U417 ( .A1(n743), .A2(n439), .A3(n617), .ZN(n654) );
  NR2D1 U418 ( .A1(n439), .A2(n834), .ZN(n467) );
  NR3D0 U419 ( .A1(n446), .A2(n439), .A3(n692), .ZN(n601) );
  ND2D1 U420 ( .A1(n439), .A2(n800), .ZN(n591) );
  ND2D1 U421 ( .A1(n439), .A2(n438), .ZN(n710) );
  NR2D1 U422 ( .A1(n72), .A2(n123), .ZN(n696) );
  AOI222D0 U423 ( .A1(n808), .A2(n824), .B1(n822), .B2(n72), .C1(n831), .C2(
        n806), .ZN(n557) );
  IND4D1 U424 ( .A1(n797), .B1(n796), .B2(n795), .B3(n794), .ZN(d[0]) );
  OAI31D0 U425 ( .A1(n801), .A2(n123), .A3(n812), .B(n860), .ZN(n495) );
  AOI31D0 U426 ( .A1(n439), .A2(n834), .A3(n812), .B(n701), .ZN(n478) );
  OR3D0 U427 ( .A1(n679), .A2(n812), .A3(n449), .Z(n640) );
  AOI22D0 U428 ( .A1(n803), .A2(n836), .B1(n812), .B2(n819), .ZN(n775) );
  NR2D1 U429 ( .A1(n782), .A2(n781), .ZN(n783) );
  AOI32D0 U430 ( .A1(n439), .A2(n839), .A3(n815), .B1(n816), .B2(n553), .ZN(
        n555) );
  AOI31D0 U431 ( .A1(n438), .A2(n827), .A3(n123), .B(n826), .ZN(n500) );
  AOI21D0 U432 ( .A1(n735), .A2(n677), .B(n438), .ZN(n635) );
  AOI22D0 U433 ( .A1(n825), .A2(n798), .B1(n823), .B2(n438), .ZN(n579) );
  ND2D1 U434 ( .A1(n438), .A2(n449), .ZN(n672) );
  NR2XD0 U435 ( .A1(n833), .A2(n829), .ZN(n681) );
  CKND2D1 U436 ( .A1(n587), .A2(n148), .ZN(d[4]) );
  CKAN2D1 U437 ( .A1(n442), .A2(n571), .Z(n434) );
  CKAN2D1 U438 ( .A1(n842), .A2(n570), .Z(n435) );
  AOI221D0 U439 ( .A1(n812), .A2(n844), .B1(n852), .B2(n817), .C(n552), .ZN(
        n588) );
  NR4D0 U440 ( .A1(n584), .A2(n583), .A3(n582), .A4(n744), .ZN(n585) );
  OAI211D0 U441 ( .A1(n709), .A2(n684), .B(n555), .C(n554), .ZN(n571) );
  OAI211D1 U442 ( .A1(n559), .A2(n430), .B(n558), .C(n557), .ZN(n570) );
  NR3D0 U443 ( .A1(n725), .A2(n439), .A3(n839), .ZN(n665) );
  NR4D0 U444 ( .A1(n447), .A2(n839), .A3(n767), .A4(n759), .ZN(n702) );
  INVD1 U445 ( .I(n728), .ZN(n843) );
  CKND2D0 U446 ( .A1(n786), .A2(n560), .ZN(n561) );
  OAI222D0 U447 ( .A1(n750), .A2(n560), .B1(n649), .B2(n430), .C1(n751), .C2(
        n692), .ZN(n459) );
  AOI22D0 U448 ( .A1(n829), .A2(n806), .B1(n803), .B2(n831), .ZN(n452) );
  NR2D1 U449 ( .A1(n515), .A2(n672), .ZN(n577) );
  OAI32D1 U450 ( .A1(n772), .A2(n479), .A3(n711), .B1(n478), .B2(n743), .ZN(
        n482) );
  NR4D0 U451 ( .A1(a[6]), .A2(n451), .A3(n732), .A4(n764), .ZN(n509) );
  OA33D0 U452 ( .A1(n713), .A2(n754), .A3(n68), .B1(n712), .B2(n711), .B3(n772), .Z(n714) );
  NR3D0 U453 ( .A1(n711), .A2(n827), .A3(n716), .ZN(n527) );
  OAI22D0 U454 ( .A1(a[6]), .A2(n439), .B1(n440), .B2(n761), .ZN(n553) );
  AOI21D0 U455 ( .A1(n779), .A2(n749), .B(n784), .ZN(n634) );
  NR4D0 U456 ( .A1(n692), .A2(n756), .A3(n784), .A4(n819), .ZN(n664) );
  OA222D1 U457 ( .A1(n686), .A2(n442), .B1(n685), .B2(n755), .C1(n684), .C2(
        n683), .Z(n437) );
  INVD1 U458 ( .I(n638), .ZN(n850) );
  INVD1 U459 ( .I(n764), .ZN(n810) );
endmodule


module aes_rcon ( clk, kld, out );
  output [31:0] out;
  input clk, kld;
  wire   N44, N45, N46, N47, N48, N49, N51, N52, N53, N54, N55, n1, n2, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n3, n22;
  wire   [2:0] rcnt;

  DFQD1 rcnt_reg_0_ ( .D(N52), .CP(clk), .Q(rcnt[0]) );
  DFKCNQD1 rcnt_reg_1_ ( .CN(n22), .D(n13), .CP(clk), .Q(rcnt[1]) );
  DFKCNQD1 rcnt_reg_2_ ( .CN(n22), .D(n2), .CP(clk), .Q(rcnt[2]) );
  DFQD1 out_reg_24_ ( .D(N44), .CP(clk), .Q(out[24]) );
  DFD1 rcnt_reg_3_ ( .D(N55), .CP(clk), .QN(n5) );
  DFQD1 out_reg_31_ ( .D(N51), .CP(clk), .Q(out[31]) );
  DFQD1 out_reg_29_ ( .D(N49), .CP(clk), .Q(out[29]) );
  DFKCNQD1 out_reg_30_ ( .CN(n1), .D(n13), .CP(clk), .Q(out[30]) );
  DFQD1 out_reg_28_ ( .D(N48), .CP(clk), .Q(out[28]) );
  DFQD1 out_reg_27_ ( .D(N47), .CP(clk), .Q(out[27]) );
  DFQD1 out_reg_26_ ( .D(N46), .CP(clk), .Q(out[26]) );
  DFQD1 out_reg_25_ ( .D(N45), .CP(clk), .Q(out[25]) );
  INVD1 U3 ( .I(n11), .ZN(n1) );
  INVD1 U4 ( .I(n14), .ZN(n2) );
  CKXOR2D1 U33 ( .A1(n14), .A2(n4), .Z(n12) );
  XNR2D1 U42 ( .A1(n6), .A2(n18), .ZN(n14) );
  CKXOR2D1 U43 ( .A1(n19), .A2(n5), .Z(n16) );
  AO21D1 U48 ( .A1(n20), .A2(n21), .B(n3), .Z(N44) );
  CKXOR2D1 U49 ( .A1(n13), .A2(rcnt[2]), .Z(n21) );
  CKXOR2D1 U52 ( .A1(rcnt[0]), .A2(rcnt[1]), .Z(n13) );
  INVD1 U5 ( .I(n22), .ZN(n3) );
  INVD1 U6 ( .I(kld), .ZN(n22) );
  ND3D1 U7 ( .A1(n7), .A2(n4), .A3(n14), .ZN(n15) );
  NR2D1 U8 ( .A1(n14), .A2(n3), .ZN(N54) );
  OAI21D1 U9 ( .A1(n7), .A2(n6), .B(n18), .ZN(n20) );
  OAI31D1 U10 ( .A1(n20), .A2(n3), .A3(n21), .B(n10), .ZN(N45) );
  OAI22D1 U11 ( .A1(n3), .A2(n15), .B1(n13), .B2(n11), .ZN(N48) );
  OAI22D1 U12 ( .A1(n9), .A2(n15), .B1(n8), .B2(n17), .ZN(N46) );
  ND3D1 U13 ( .A1(n16), .A2(n14), .A3(N53), .ZN(n17) );
  NR2D1 U14 ( .A1(n7), .A2(n3), .ZN(N53) );
  INVD1 U15 ( .I(n13), .ZN(n7) );
  NR3D0 U16 ( .A1(n9), .A2(n12), .A3(n13), .ZN(N49) );
  INVD1 U17 ( .I(n16), .ZN(n4) );
  INVD1 U18 ( .I(N52), .ZN(n9) );
  OAI32D1 U19 ( .A1(n15), .A2(n3), .A3(n8), .B1(rcnt[0]), .B2(n17), .ZN(N47)
         );
  NR2D1 U20 ( .A1(n6), .A2(n18), .ZN(n19) );
  INR4D0 U21 ( .A1(N54), .B1(rcnt[0]), .B2(n7), .B3(n4), .ZN(N51) );
  IND4D1 U22 ( .A1(n3), .B1(n21), .B2(n20), .B3(n5), .ZN(n10) );
  ND3D1 U23 ( .A1(n16), .A2(rcnt[0]), .A3(N54), .ZN(n11) );
  ND2D1 U24 ( .A1(rcnt[0]), .A2(rcnt[1]), .ZN(n18) );
  NR2D1 U25 ( .A1(n3), .A2(rcnt[0]), .ZN(N52) );
  INVD1 U26 ( .I(rcnt[0]), .ZN(n8) );
  OAI21D1 U27 ( .A1(N44), .A2(n5), .B(n10), .ZN(N55) );
  INVD1 U28 ( .I(rcnt[2]), .ZN(n6) );
endmodule


module aes_key_expand_128 ( clk, kld, key, wo_0, wo_1, wo_2, wo_3 );
  input [127:0] key;
  output [31:0] wo_0;
  output [31:0] wo_1;
  output [31:0] wo_2;
  output [31:0] wo_3;
  input clk, kld;
  wire   n209, n210, n211, n212, n213, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n66, n67,
         n68, n69, n70, n72, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n88, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n120, n121, n122, n123, n124,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n65, n71, n73, n77, n87, n89, n103, n119, n125, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n198, n199, n201, n203, n205, n207, n208,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24;
  wire   [31:0] subword;
  wire   [31:24] rcon;

  aes_sbox_4 u0 ( .a(wo_3[23:16]), .d(subword[31:24]) );
  aes_sbox_3 u1 ( .a(wo_3[15:8]), .d(subword[23:16]) );
  aes_sbox_2 u2 ( .a(wo_3[7:0]), .d(subword[15:8]) );
  aes_sbox_1 u3 ( .a(wo_3[31:24]), .d(subword[7:0]) );
  aes_rcon r0 ( .clk(clk), .kld(n194), .out({rcon, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24}) );
  DFQD1 w_reg_0__8_ ( .D(N50), .CP(clk), .Q(wo_0[8]) );
  DFQD1 w_reg_2__8_ ( .D(N182), .CP(clk), .Q(wo_2[8]) );
  DFQD1 w_reg_1__8_ ( .D(N116), .CP(clk), .Q(wo_1[8]) );
  DFQD1 w_reg_0__9_ ( .D(N51), .CP(clk), .Q(wo_0[9]) );
  DFQD1 w_reg_2__9_ ( .D(N183), .CP(clk), .Q(wo_2[9]) );
  DFQD1 w_reg_1__9_ ( .D(N117), .CP(clk), .Q(wo_1[9]) );
  DFQD1 w_reg_0__10_ ( .D(N52), .CP(clk), .Q(wo_0[10]) );
  DFQD1 w_reg_2__10_ ( .D(N184), .CP(clk), .Q(wo_2[10]) );
  DFQD1 w_reg_1__10_ ( .D(N118), .CP(clk), .Q(wo_1[10]) );
  DFQD1 w_reg_0__11_ ( .D(N53), .CP(clk), .Q(wo_0[11]) );
  DFQD1 w_reg_2__11_ ( .D(N185), .CP(clk), .Q(wo_2[11]) );
  DFQD1 w_reg_1__11_ ( .D(N119), .CP(clk), .Q(wo_1[11]) );
  DFQD1 w_reg_0__12_ ( .D(N54), .CP(clk), .Q(wo_0[12]) );
  DFQD1 w_reg_2__12_ ( .D(N186), .CP(clk), .Q(wo_2[12]) );
  DFQD1 w_reg_1__12_ ( .D(N120), .CP(clk), .Q(wo_1[12]) );
  DFQD1 w_reg_0__13_ ( .D(N55), .CP(clk), .Q(wo_0[13]) );
  DFQD1 w_reg_2__13_ ( .D(N187), .CP(clk), .Q(wo_2[13]) );
  DFQD1 w_reg_1__13_ ( .D(N121), .CP(clk), .Q(wo_1[13]) );
  DFQD1 w_reg_0__14_ ( .D(N56), .CP(clk), .Q(wo_0[14]) );
  DFQD1 w_reg_2__14_ ( .D(N188), .CP(clk), .Q(wo_2[14]) );
  DFQD1 w_reg_1__14_ ( .D(N122), .CP(clk), .Q(wo_1[14]) );
  DFQD1 w_reg_0__15_ ( .D(N57), .CP(clk), .Q(wo_0[15]) );
  DFQD1 w_reg_2__15_ ( .D(N189), .CP(clk), .Q(wo_2[15]) );
  DFQD1 w_reg_0__16_ ( .D(N58), .CP(clk), .Q(wo_0[16]) );
  DFQD1 w_reg_2__16_ ( .D(N190), .CP(clk), .Q(wo_2[16]) );
  DFQD1 w_reg_1__16_ ( .D(N124), .CP(clk), .Q(wo_1[16]) );
  DFQD1 w_reg_0__17_ ( .D(N59), .CP(clk), .Q(wo_0[17]) );
  DFQD1 w_reg_2__17_ ( .D(N191), .CP(clk), .Q(wo_2[17]) );
  DFQD1 w_reg_0__18_ ( .D(N60), .CP(clk), .Q(wo_0[18]) );
  DFQD1 w_reg_2__18_ ( .D(N192), .CP(clk), .Q(wo_2[18]) );
  DFQD1 w_reg_1__18_ ( .D(N126), .CP(clk), .Q(wo_1[18]) );
  DFQD1 w_reg_0__19_ ( .D(N61), .CP(clk), .Q(wo_0[19]) );
  DFQD1 w_reg_2__19_ ( .D(N193), .CP(clk), .Q(wo_2[19]) );
  DFQD1 w_reg_1__19_ ( .D(N127), .CP(clk), .Q(wo_1[19]) );
  DFQD1 w_reg_0__20_ ( .D(N62), .CP(clk), .Q(wo_0[20]) );
  DFQD1 w_reg_2__20_ ( .D(N194), .CP(clk), .Q(wo_2[20]) );
  DFQD1 w_reg_0__21_ ( .D(N63), .CP(clk), .Q(wo_0[21]) );
  DFQD1 w_reg_2__21_ ( .D(N195), .CP(clk), .Q(wo_2[21]) );
  DFQD1 w_reg_3__21_ ( .D(N261), .CP(clk), .Q(wo_3[21]) );
  DFQD1 w_reg_1__21_ ( .D(N129), .CP(clk), .Q(wo_1[21]) );
  DFQD1 w_reg_0__22_ ( .D(N64), .CP(clk), .Q(wo_0[22]) );
  DFQD1 w_reg_2__22_ ( .D(N196), .CP(clk), .Q(wo_2[22]) );
  DFQD1 w_reg_1__22_ ( .D(N130), .CP(clk), .Q(wo_1[22]) );
  DFQD1 w_reg_0__23_ ( .D(N65), .CP(clk), .Q(wo_0[23]) );
  DFQD1 w_reg_2__23_ ( .D(N197), .CP(clk), .Q(wo_2[23]) );
  DFQD1 w_reg_3__23_ ( .D(N263), .CP(clk), .Q(wo_3[23]) );
  DFQD1 w_reg_0__24_ ( .D(N66), .CP(clk), .Q(wo_0[24]) );
  DFQD1 w_reg_2__24_ ( .D(N198), .CP(clk), .Q(wo_2[24]) );
  DFQD1 w_reg_1__24_ ( .D(N132), .CP(clk), .Q(wo_1[24]) );
  DFQD1 w_reg_0__25_ ( .D(N67), .CP(clk), .Q(wo_0[25]) );
  DFQD1 w_reg_2__25_ ( .D(N199), .CP(clk), .Q(wo_2[25]) );
  DFQD1 w_reg_1__25_ ( .D(N133), .CP(clk), .Q(wo_1[25]) );
  DFQD1 w_reg_0__26_ ( .D(N68), .CP(clk), .Q(wo_0[26]) );
  DFQD1 w_reg_2__26_ ( .D(N200), .CP(clk), .Q(wo_2[26]) );
  DFQD1 w_reg_1__26_ ( .D(N134), .CP(clk), .Q(wo_1[26]) );
  DFQD1 w_reg_0__27_ ( .D(N69), .CP(clk), .Q(wo_0[27]) );
  DFQD1 w_reg_2__27_ ( .D(N201), .CP(clk), .Q(wo_2[27]) );
  DFQD1 w_reg_1__27_ ( .D(N135), .CP(clk), .Q(wo_1[27]) );
  DFQD1 w_reg_0__28_ ( .D(N70), .CP(clk), .Q(wo_0[28]) );
  DFQD1 w_reg_2__28_ ( .D(N202), .CP(clk), .Q(wo_2[28]) );
  DFQD1 w_reg_1__28_ ( .D(N136), .CP(clk), .Q(wo_1[28]) );
  DFQD1 w_reg_0__29_ ( .D(N71), .CP(clk), .Q(wo_0[29]) );
  DFQD1 w_reg_2__29_ ( .D(N203), .CP(clk), .Q(wo_2[29]) );
  DFQD1 w_reg_1__29_ ( .D(N137), .CP(clk), .Q(wo_1[29]) );
  DFQD1 w_reg_0__30_ ( .D(N72), .CP(clk), .Q(wo_0[30]) );
  DFQD1 w_reg_2__30_ ( .D(N204), .CP(clk), .Q(wo_2[30]) );
  DFQD1 w_reg_1__30_ ( .D(N138), .CP(clk), .Q(wo_1[30]) );
  DFQD1 w_reg_0__31_ ( .D(N73), .CP(clk), .Q(wo_0[31]) );
  DFQD1 w_reg_2__31_ ( .D(N205), .CP(clk), .Q(wo_2[31]) );
  DFQD1 w_reg_3__31_ ( .D(N271), .CP(clk), .Q(wo_3[31]) );
  DFQD1 w_reg_0__0_ ( .D(N42), .CP(clk), .Q(wo_0[0]) );
  DFQD1 w_reg_2__0_ ( .D(N174), .CP(clk), .Q(wo_2[0]) );
  DFQD1 w_reg_1__0_ ( .D(N108), .CP(clk), .Q(wo_1[0]) );
  DFQD1 w_reg_0__1_ ( .D(N43), .CP(clk), .Q(wo_0[1]) );
  DFQD1 w_reg_2__1_ ( .D(N175), .CP(clk), .Q(wo_2[1]) );
  DFQD1 w_reg_1__1_ ( .D(N109), .CP(clk), .Q(wo_1[1]) );
  DFQD1 w_reg_0__2_ ( .D(N44), .CP(clk), .Q(wo_0[2]) );
  DFQD1 w_reg_2__2_ ( .D(N176), .CP(clk), .Q(wo_2[2]) );
  DFQD1 w_reg_1__2_ ( .D(N110), .CP(clk), .Q(wo_1[2]) );
  DFQD1 w_reg_0__3_ ( .D(N45), .CP(clk), .Q(wo_0[3]) );
  DFQD1 w_reg_2__3_ ( .D(N177), .CP(clk), .Q(wo_2[3]) );
  DFQD1 w_reg_1__3_ ( .D(N111), .CP(clk), .Q(wo_1[3]) );
  DFQD1 w_reg_0__4_ ( .D(N46), .CP(clk), .Q(wo_0[4]) );
  DFQD1 w_reg_2__4_ ( .D(N178), .CP(clk), .Q(wo_2[4]) );
  DFQD1 w_reg_1__4_ ( .D(N112), .CP(clk), .Q(wo_1[4]) );
  DFQD1 w_reg_0__5_ ( .D(N47), .CP(clk), .Q(wo_0[5]) );
  DFQD1 w_reg_2__5_ ( .D(N179), .CP(clk), .Q(wo_2[5]) );
  DFQD1 w_reg_1__5_ ( .D(N113), .CP(clk), .Q(wo_1[5]) );
  DFQD1 w_reg_0__6_ ( .D(N48), .CP(clk), .Q(wo_0[6]) );
  DFQD1 w_reg_2__6_ ( .D(N180), .CP(clk), .Q(wo_2[6]) );
  DFQD1 w_reg_1__6_ ( .D(N114), .CP(clk), .Q(wo_1[6]) );
  DFQD1 w_reg_0__7_ ( .D(N49), .CP(clk), .Q(wo_0[7]) );
  DFQD1 w_reg_2__7_ ( .D(N181), .CP(clk), .Q(wo_2[7]) );
  DFQD1 w_reg_1__7_ ( .D(N115), .CP(clk), .Q(wo_1[7]) );
  DFQD1 w_reg_1__31_ ( .D(N139), .CP(clk), .Q(wo_1[31]) );
  DFQD1 w_reg_1__23_ ( .D(N131), .CP(clk), .Q(wo_1[23]) );
  DFQD1 w_reg_1__15_ ( .D(N123), .CP(clk), .Q(wo_1[15]) );
  MOAI22D1 U3 ( .A1(n208), .A2(n1), .B1(n208), .B2(key[127]), .ZN(N73) );
  XNR2D1 U4 ( .A1(n2), .A2(rcon[31]), .ZN(n1) );
  MOAI22D1 U5 ( .A1(n208), .A2(n3), .B1(key[126]), .B2(n196), .ZN(N72) );
  XNR2D1 U6 ( .A1(n4), .A2(rcon[30]), .ZN(n3) );
  MOAI22D1 U7 ( .A1(n208), .A2(n5), .B1(key[125]), .B2(n196), .ZN(N71) );
  XNR2D1 U8 ( .A1(n6), .A2(rcon[29]), .ZN(n5) );
  MOAI22D1 U9 ( .A1(n208), .A2(n7), .B1(key[124]), .B2(n196), .ZN(N70) );
  XNR2D1 U10 ( .A1(n8), .A2(rcon[28]), .ZN(n7) );
  MOAI22D1 U11 ( .A1(n208), .A2(n9), .B1(key[123]), .B2(n196), .ZN(N69) );
  XNR2D1 U12 ( .A1(n10), .A2(rcon[27]), .ZN(n9) );
  MOAI22D1 U13 ( .A1(n208), .A2(n11), .B1(key[122]), .B2(n195), .ZN(N68) );
  XNR2D1 U14 ( .A1(n12), .A2(rcon[26]), .ZN(n11) );
  MOAI22D1 U15 ( .A1(n208), .A2(n13), .B1(key[121]), .B2(n195), .ZN(N67) );
  XNR2D1 U16 ( .A1(n14), .A2(rcon[25]), .ZN(n13) );
  MOAI22D1 U17 ( .A1(n195), .A2(n15), .B1(key[120]), .B2(n194), .ZN(N66) );
  XNR2D1 U18 ( .A1(n16), .A2(rcon[24]), .ZN(n15) );
  MOAI22D1 U19 ( .A1(n194), .A2(n17), .B1(key[119]), .B2(n195), .ZN(N65) );
  MOAI22D1 U21 ( .A1(n208), .A2(n19), .B1(key[118]), .B2(n195), .ZN(N64) );
  MOAI22D1 U23 ( .A1(n208), .A2(n21), .B1(key[117]), .B2(n194), .ZN(N63) );
  MOAI22D1 U25 ( .A1(n196), .A2(n23), .B1(key[116]), .B2(n195), .ZN(N62) );
  MOAI22D1 U27 ( .A1(n208), .A2(n25), .B1(key[115]), .B2(n196), .ZN(N61) );
  MOAI22D1 U29 ( .A1(n194), .A2(n27), .B1(key[114]), .B2(n196), .ZN(N60) );
  MOAI22D1 U31 ( .A1(n196), .A2(n29), .B1(key[113]), .B2(n196), .ZN(N59) );
  MOAI22D1 U33 ( .A1(n208), .A2(n31), .B1(key[112]), .B2(n195), .ZN(N58) );
  MOAI22D1 U35 ( .A1(n196), .A2(n33), .B1(key[111]), .B2(n194), .ZN(N57) );
  MOAI22D1 U37 ( .A1(n195), .A2(n35), .B1(key[110]), .B2(n195), .ZN(N56) );
  MOAI22D1 U39 ( .A1(n208), .A2(n37), .B1(key[109]), .B2(n194), .ZN(N55) );
  MOAI22D1 U41 ( .A1(n196), .A2(n39), .B1(key[108]), .B2(n194), .ZN(N54) );
  MOAI22D1 U43 ( .A1(n194), .A2(n41), .B1(key[107]), .B2(n194), .ZN(N53) );
  MOAI22D1 U45 ( .A1(n195), .A2(n43), .B1(key[106]), .B2(n194), .ZN(N52) );
  MOAI22D1 U47 ( .A1(n195), .A2(n45), .B1(key[105]), .B2(n194), .ZN(N51) );
  MOAI22D1 U49 ( .A1(n194), .A2(n47), .B1(key[104]), .B2(n194), .ZN(N50) );
  MOAI22D1 U51 ( .A1(n195), .A2(n49), .B1(key[103]), .B2(n194), .ZN(N49) );
  MOAI22D1 U53 ( .A1(n196), .A2(n51), .B1(key[102]), .B2(n194), .ZN(N48) );
  MOAI22D1 U55 ( .A1(n195), .A2(n53), .B1(key[101]), .B2(n194), .ZN(N47) );
  MOAI22D1 U57 ( .A1(n194), .A2(n55), .B1(key[100]), .B2(n194), .ZN(N46) );
  MOAI22D1 U59 ( .A1(n195), .A2(n57), .B1(key[99]), .B2(n194), .ZN(N45) );
  MOAI22D1 U61 ( .A1(n194), .A2(n59), .B1(key[98]), .B2(n194), .ZN(N44) );
  MOAI22D1 U63 ( .A1(n196), .A2(n61), .B1(key[97]), .B2(n194), .ZN(N43) );
  MOAI22D1 U65 ( .A1(n208), .A2(n63), .B1(key[96]), .B2(n194), .ZN(N42) );
  MOAI22D1 U69 ( .A1(n194), .A2(n67), .B1(key[30]), .B2(n194), .ZN(N270) );
  MOAI22D1 U71 ( .A1(n208), .A2(n69), .B1(key[29]), .B2(n194), .ZN(N269) );
  MOAI22D1 U77 ( .A1(n208), .A2(n75), .B1(key[26]), .B2(n194), .ZN(N266) );
  MOAI22D1 U81 ( .A1(n208), .A2(n79), .B1(key[24]), .B2(n194), .ZN(N264) );
  MOAI22D1 U85 ( .A1(n208), .A2(n83), .B1(key[22]), .B2(n194), .ZN(N262) );
  MOAI22D1 U87 ( .A1(n208), .A2(n85), .B1(key[21]), .B2(n195), .ZN(N261) );
  MOAI22D1 U93 ( .A1(n208), .A2(n91), .B1(key[18]), .B2(n195), .ZN(N258) );
  MOAI22D1 U97 ( .A1(n208), .A2(n95), .B1(key[16]), .B2(n195), .ZN(N256) );
  MOAI22D1 U99 ( .A1(n208), .A2(n97), .B1(key[15]), .B2(n196), .ZN(N255) );
  MOAI22D1 U101 ( .A1(n208), .A2(n99), .B1(key[14]), .B2(n195), .ZN(N254) );
  MOAI22D1 U103 ( .A1(n208), .A2(n101), .B1(key[13]), .B2(n196), .ZN(N253) );
  MOAI22D1 U109 ( .A1(n208), .A2(n107), .B1(key[10]), .B2(n195), .ZN(N250) );
  MOAI22D1 U113 ( .A1(n208), .A2(n111), .B1(key[8]), .B2(n195), .ZN(N248) );
  MOAI22D1 U117 ( .A1(n208), .A2(n115), .B1(key[6]), .B2(n195), .ZN(N246) );
  MOAI22D1 U119 ( .A1(n208), .A2(n117), .B1(key[5]), .B2(n196), .ZN(N245) );
  MOAI22D1 U123 ( .A1(n208), .A2(n121), .B1(key[3]), .B2(n196), .ZN(N243) );
  MOAI22D1 U125 ( .A1(n208), .A2(n123), .B1(key[2]), .B2(n195), .ZN(N242) );
  MOAI22D1 U129 ( .A1(n208), .A2(n127), .B1(key[0]), .B2(n195), .ZN(N240) );
  MOAI22D1 U131 ( .A1(n208), .A2(n129), .B1(key[63]), .B2(n196), .ZN(N205) );
  CKXOR2D1 U132 ( .A1(n66), .A2(wo_2[31]), .Z(n129) );
  MOAI22D1 U133 ( .A1(n208), .A2(n130), .B1(key[62]), .B2(n195), .ZN(N204) );
  CKXOR2D1 U134 ( .A1(n68), .A2(wo_2[30]), .Z(n130) );
  MOAI22D1 U135 ( .A1(n208), .A2(n131), .B1(key[61]), .B2(n196), .ZN(N203) );
  CKXOR2D1 U136 ( .A1(n70), .A2(wo_2[29]), .Z(n131) );
  MOAI22D1 U137 ( .A1(n208), .A2(n132), .B1(key[60]), .B2(n195), .ZN(N202) );
  CKXOR2D1 U138 ( .A1(n72), .A2(wo_2[28]), .Z(n132) );
  MOAI22D1 U139 ( .A1(n208), .A2(n133), .B1(key[59]), .B2(n196), .ZN(N201) );
  CKXOR2D1 U140 ( .A1(n74), .A2(wo_2[27]), .Z(n133) );
  MOAI22D1 U141 ( .A1(n208), .A2(n134), .B1(key[58]), .B2(n195), .ZN(N200) );
  CKXOR2D1 U142 ( .A1(n76), .A2(wo_2[26]), .Z(n134) );
  MOAI22D1 U143 ( .A1(n208), .A2(n135), .B1(key[57]), .B2(n196), .ZN(N199) );
  MOAI22D1 U145 ( .A1(n208), .A2(n136), .B1(key[56]), .B2(n195), .ZN(N198) );
  CKXOR2D1 U146 ( .A1(n80), .A2(wo_2[24]), .Z(n136) );
  MOAI22D1 U147 ( .A1(n208), .A2(n137), .B1(key[55]), .B2(n196), .ZN(N197) );
  CKXOR2D1 U148 ( .A1(n82), .A2(wo_2[23]), .Z(n137) );
  MOAI22D1 U149 ( .A1(n208), .A2(n138), .B1(key[54]), .B2(n195), .ZN(N196) );
  CKXOR2D1 U150 ( .A1(n84), .A2(wo_2[22]), .Z(n138) );
  MOAI22D1 U151 ( .A1(n208), .A2(n139), .B1(key[53]), .B2(n196), .ZN(N195) );
  CKXOR2D1 U152 ( .A1(n86), .A2(wo_2[21]), .Z(n139) );
  MOAI22D1 U153 ( .A1(n208), .A2(n140), .B1(key[52]), .B2(n195), .ZN(N194) );
  CKXOR2D1 U154 ( .A1(n168), .A2(wo_2[20]), .Z(n140) );
  MOAI22D1 U155 ( .A1(n208), .A2(n141), .B1(key[51]), .B2(n196), .ZN(N193) );
  MOAI22D1 U157 ( .A1(n208), .A2(n142), .B1(key[50]), .B2(n195), .ZN(N192) );
  CKXOR2D1 U158 ( .A1(n92), .A2(wo_2[18]), .Z(n142) );
  MOAI22D1 U159 ( .A1(n208), .A2(n143), .B1(key[49]), .B2(n196), .ZN(N191) );
  MOAI22D1 U161 ( .A1(n208), .A2(n144), .B1(key[48]), .B2(n195), .ZN(N190) );
  CKXOR2D1 U162 ( .A1(n96), .A2(wo_2[16]), .Z(n144) );
  MOAI22D1 U163 ( .A1(n208), .A2(n145), .B1(key[47]), .B2(n196), .ZN(N189) );
  CKXOR2D1 U164 ( .A1(n98), .A2(wo_2[15]), .Z(n145) );
  MOAI22D1 U165 ( .A1(n208), .A2(n146), .B1(key[46]), .B2(n195), .ZN(N188) );
  CKXOR2D1 U166 ( .A1(n100), .A2(wo_2[14]), .Z(n146) );
  MOAI22D1 U167 ( .A1(n208), .A2(n147), .B1(key[45]), .B2(n196), .ZN(N187) );
  CKXOR2D1 U168 ( .A1(n102), .A2(wo_2[13]), .Z(n147) );
  MOAI22D1 U169 ( .A1(n208), .A2(n148), .B1(key[44]), .B2(n195), .ZN(N186) );
  MOAI22D1 U171 ( .A1(n208), .A2(n149), .B1(key[43]), .B2(n196), .ZN(N185) );
  MOAI22D1 U173 ( .A1(n208), .A2(n150), .B1(key[42]), .B2(n195), .ZN(N184) );
  CKXOR2D1 U174 ( .A1(n108), .A2(wo_2[10]), .Z(n150) );
  MOAI22D1 U175 ( .A1(n208), .A2(n151), .B1(key[41]), .B2(n196), .ZN(N183) );
  CKXOR2D1 U176 ( .A1(n110), .A2(wo_2[9]), .Z(n151) );
  MOAI22D1 U177 ( .A1(n208), .A2(n152), .B1(key[40]), .B2(n195), .ZN(N182) );
  CKXOR2D1 U178 ( .A1(n112), .A2(wo_2[8]), .Z(n152) );
  MOAI22D1 U179 ( .A1(n208), .A2(n153), .B1(key[39]), .B2(n196), .ZN(N181) );
  CKXOR2D1 U180 ( .A1(n114), .A2(wo_2[7]), .Z(n153) );
  MOAI22D1 U181 ( .A1(n208), .A2(n154), .B1(key[38]), .B2(n195), .ZN(N180) );
  CKXOR2D1 U182 ( .A1(n116), .A2(wo_2[6]), .Z(n154) );
  MOAI22D1 U183 ( .A1(n208), .A2(n155), .B1(key[37]), .B2(n196), .ZN(N179) );
  CKXOR2D1 U184 ( .A1(n118), .A2(wo_2[5]), .Z(n155) );
  MOAI22D1 U185 ( .A1(n208), .A2(n156), .B1(key[36]), .B2(n196), .ZN(N178) );
  CKXOR2D1 U186 ( .A1(n120), .A2(wo_2[4]), .Z(n156) );
  MOAI22D1 U187 ( .A1(n208), .A2(n157), .B1(key[35]), .B2(n194), .ZN(N177) );
  MOAI22D1 U189 ( .A1(n208), .A2(n158), .B1(key[34]), .B2(n196), .ZN(N176) );
  CKXOR2D1 U190 ( .A1(n124), .A2(wo_2[2]), .Z(n158) );
  MOAI22D1 U191 ( .A1(n208), .A2(n159), .B1(key[33]), .B2(n194), .ZN(N175) );
  MOAI22D1 U193 ( .A1(n208), .A2(n160), .B1(key[32]), .B2(n195), .ZN(N174) );
  CKXOR2D1 U194 ( .A1(n128), .A2(wo_2[0]), .Z(n160) );
  MOAI22D1 U195 ( .A1(n208), .A2(n66), .B1(key[95]), .B2(n194), .ZN(N139) );
  CKXOR2D1 U197 ( .A1(subword[31]), .A2(wo_0[31]), .Z(n2) );
  MOAI22D1 U198 ( .A1(n208), .A2(n68), .B1(key[94]), .B2(n194), .ZN(N138) );
  CKXOR2D1 U200 ( .A1(subword[30]), .A2(wo_0[30]), .Z(n4) );
  CKXOR2D1 U203 ( .A1(wo_0[29]), .A2(subword[29]), .Z(n6) );
  MOAI22D1 U204 ( .A1(n208), .A2(n72), .B1(key[92]), .B2(n194), .ZN(N136) );
  CKXOR2D1 U209 ( .A1(subword[27]), .A2(wo_0[27]), .Z(n10) );
  MOAI22D1 U210 ( .A1(n208), .A2(n76), .B1(key[90]), .B2(n196), .ZN(N134) );
  CKXOR2D1 U212 ( .A1(subword[26]), .A2(wo_0[26]), .Z(n12) );
  MOAI22D1 U216 ( .A1(n208), .A2(n80), .B1(key[88]), .B2(n195), .ZN(N132) );
  CKXOR2D1 U218 ( .A1(subword[24]), .A2(wo_0[24]), .Z(n16) );
  MOAI22D1 U219 ( .A1(n208), .A2(n82), .B1(key[87]), .B2(n196), .ZN(N131) );
  CKXOR2D1 U221 ( .A1(wo_0[23]), .A2(subword[23]), .Z(n18) );
  MOAI22D1 U222 ( .A1(n208), .A2(n84), .B1(key[86]), .B2(n196), .ZN(N130) );
  CKXOR2D1 U224 ( .A1(wo_0[22]), .A2(subword[22]), .Z(n20) );
  MOAI22D1 U225 ( .A1(n208), .A2(n86), .B1(key[85]), .B2(n196), .ZN(N129) );
  CKXOR2D1 U227 ( .A1(wo_0[21]), .A2(subword[21]), .Z(n22) );
  CKXOR2D1 U230 ( .A1(subword[20]), .A2(wo_0[20]), .Z(n24) );
  MOAI22D1 U234 ( .A1(n208), .A2(n92), .B1(key[82]), .B2(n196), .ZN(N126) );
  CKXOR2D1 U236 ( .A1(wo_0[18]), .A2(subword[18]), .Z(n28) );
  CKXOR2D1 U239 ( .A1(subword[17]), .A2(wo_0[17]), .Z(n30) );
  MOAI22D1 U240 ( .A1(n208), .A2(n96), .B1(key[80]), .B2(n195), .ZN(N124) );
  CKXOR2D1 U242 ( .A1(subword[16]), .A2(wo_0[16]), .Z(n32) );
  MOAI22D1 U243 ( .A1(n208), .A2(n98), .B1(key[79]), .B2(n195), .ZN(N123) );
  CKXOR2D1 U245 ( .A1(subword[15]), .A2(wo_0[15]), .Z(n34) );
  MOAI22D1 U246 ( .A1(n208), .A2(n100), .B1(key[78]), .B2(n196), .ZN(N122) );
  CKXOR2D1 U248 ( .A1(wo_0[14]), .A2(subword[14]), .Z(n36) );
  MOAI22D1 U249 ( .A1(n208), .A2(n102), .B1(key[77]), .B2(n196), .ZN(N121) );
  CKXOR2D1 U251 ( .A1(wo_0[13]), .A2(subword[13]), .Z(n38) );
  CKXOR2D1 U254 ( .A1(subword[12]), .A2(wo_0[12]), .Z(n40) );
  CKXOR2D1 U257 ( .A1(wo_0[11]), .A2(subword[11]), .Z(n42) );
  MOAI22D1 U258 ( .A1(n208), .A2(n108), .B1(key[74]), .B2(n196), .ZN(N118) );
  CKXOR2D1 U260 ( .A1(wo_0[10]), .A2(subword[10]), .Z(n44) );
  MOAI22D1 U264 ( .A1(n208), .A2(n112), .B1(key[72]), .B2(n196), .ZN(N116) );
  CKXOR2D1 U266 ( .A1(wo_0[8]), .A2(subword[8]), .Z(n48) );
  MOAI22D1 U267 ( .A1(n208), .A2(n114), .B1(key[71]), .B2(n195), .ZN(N115) );
  CKXOR2D1 U269 ( .A1(wo_0[7]), .A2(subword[7]), .Z(n50) );
  MOAI22D1 U270 ( .A1(n208), .A2(n116), .B1(key[70]), .B2(n195), .ZN(N114) );
  CKXOR2D1 U272 ( .A1(wo_0[6]), .A2(subword[6]), .Z(n52) );
  MOAI22D1 U273 ( .A1(n208), .A2(n118), .B1(key[69]), .B2(n196), .ZN(N113) );
  CKXOR2D1 U275 ( .A1(wo_0[5]), .A2(subword[5]), .Z(n54) );
  MOAI22D1 U276 ( .A1(n208), .A2(n120), .B1(key[68]), .B2(n195), .ZN(N112) );
  CKXOR2D1 U278 ( .A1(wo_0[4]), .A2(subword[4]), .Z(n56) );
  CKXOR2D1 U281 ( .A1(wo_0[3]), .A2(subword[3]), .Z(n58) );
  MOAI22D1 U282 ( .A1(n208), .A2(n124), .B1(key[66]), .B2(n195), .ZN(N110) );
  CKXOR2D1 U284 ( .A1(wo_0[2]), .A2(subword[2]), .Z(n60) );
  MOAI22D1 U288 ( .A1(n208), .A2(n128), .B1(key[64]), .B2(n196), .ZN(N108) );
  CKXOR2D1 U290 ( .A1(wo_0[0]), .A2(subword[0]), .Z(n64) );
  DFQD4 w_reg_3__17_ ( .D(N257), .CP(clk), .Q(wo_3[17]) );
  DFQD4 w_reg_3__11_ ( .D(N251), .CP(clk), .Q(wo_3[11]) );
  DFQD1 w_reg_3__24_ ( .D(N264), .CP(clk), .Q(n209) );
  DFQD1 w_reg_3__1_ ( .D(N241), .CP(clk), .Q(wo_3[1]) );
  DFQD1 w_reg_3__16_ ( .D(N256), .CP(clk), .Q(n211) );
  DFQD1 w_reg_3__8_ ( .D(N248), .CP(clk), .Q(n212) );
  DFQD1 w_reg_3__0_ ( .D(N240), .CP(clk), .Q(n213) );
  DFQD1 w_reg_3__12_ ( .D(N252), .CP(clk), .Q(wo_3[12]) );
  DFQD1 w_reg_3__19_ ( .D(N259), .CP(clk), .Q(n210) );
  DFQD1 w_reg_3__7_ ( .D(N247), .CP(clk), .Q(wo_3[7]) );
  DFQD1 w_reg_3__15_ ( .D(N255), .CP(clk), .Q(wo_3[15]) );
  DFQD1 w_reg_3__20_ ( .D(N260), .CP(clk), .Q(wo_3[20]) );
  DFQD1 w_reg_3__6_ ( .D(N246), .CP(clk), .Q(wo_3[6]) );
  DFQD1 w_reg_3__2_ ( .D(N242), .CP(clk), .Q(wo_3[2]) );
  DFQD1 w_reg_3__4_ ( .D(N244), .CP(clk), .Q(wo_3[4]) );
  DFQD4 w_reg_3__10_ ( .D(N250), .CP(clk), .Q(wo_3[10]) );
  DFQD4 w_reg_3__18_ ( .D(N258), .CP(clk), .Q(wo_3[18]) );
  DFQD2 w_reg_3__25_ ( .D(N265), .CP(clk), .Q(wo_3[25]) );
  DFQD2 w_reg_3__27_ ( .D(N267), .CP(clk), .Q(wo_3[27]) );
  DFQD2 w_reg_3__30_ ( .D(N270), .CP(clk), .Q(wo_3[30]) );
  DFQD4 w_reg_3__5_ ( .D(N245), .CP(clk), .Q(wo_3[5]) );
  DFQD1 w_reg_3__28_ ( .D(N268), .CP(clk), .Q(wo_3[28]) );
  DFQD2 w_reg_3__26_ ( .D(N266), .CP(clk), .Q(wo_3[26]) );
  DFQD1 w_reg_3__9_ ( .D(N249), .CP(clk), .Q(wo_3[9]) );
  DFQD1 w_reg_1__20_ ( .D(N128), .CP(clk), .Q(wo_1[20]) );
  DFQD1 w_reg_3__3_ ( .D(N243), .CP(clk), .Q(wo_3[3]) );
  DFQD2 w_reg_3__22_ ( .D(N262), .CP(clk), .Q(wo_3[22]) );
  DFQD4 w_reg_3__13_ ( .D(N253), .CP(clk), .Q(wo_3[13]) );
  DFQD4 w_reg_1__17_ ( .D(N125), .CP(clk), .Q(wo_1[17]) );
  DFQD2 w_reg_3__14_ ( .D(N254), .CP(clk), .Q(wo_3[14]) );
  DFQD2 w_reg_3__29_ ( .D(N269), .CP(clk), .Q(wo_3[29]) );
  CKXOR2D1 U20 ( .A1(n122), .A2(wo_2[3]), .Z(n157) );
  MOAI22D0 U22 ( .A1(n208), .A2(n122), .B1(key[67]), .B2(n196), .ZN(N111) );
  MOAI22D1 U24 ( .A1(n65), .A2(n71), .B1(n77), .B2(n73), .ZN(N259) );
  INVD16 U26 ( .I(key[19]), .ZN(n65) );
  INVD16 U28 ( .I(n196), .ZN(n71) );
  XNR3D4 U30 ( .A1(wo_3[19]), .A2(wo_2[19]), .A3(n90), .ZN(n73) );
  MOAI22D1 U32 ( .A1(n87), .A2(n77), .B1(n77), .B2(n89), .ZN(N244) );
  INVD12 U34 ( .I(n208), .ZN(n77) );
  INVD16 U36 ( .I(key[4]), .ZN(n87) );
  XNR3D1 U38 ( .A1(wo_3[4]), .A2(wo_2[4]), .A3(n120), .ZN(n89) );
  MOAI22D1 U40 ( .A1(n103), .A2(n119), .B1(key[28]), .B2(n194), .ZN(N268) );
  INVD16 U42 ( .I(n187), .ZN(n103) );
  XOR3D1 U44 ( .A1(wo_3[28]), .A2(wo_2[28]), .A3(n72), .Z(n119) );
  XOR3D4 U46 ( .A1(wo_3[13]), .A2(wo_2[13]), .A3(n102), .Z(n101) );
  XOR3D4 U48 ( .A1(wo_3[24]), .A2(wo_2[24]), .A3(n80), .Z(n79) );
  XNR2D1 U50 ( .A1(wo_1[17]), .A2(n30), .ZN(n125) );
  CKXOR2D1 U52 ( .A1(n126), .A2(wo_2[1]), .Z(n159) );
  CKXOR2D1 U54 ( .A1(n104), .A2(wo_2[12]), .Z(n148) );
  MOAI22D2 U56 ( .A1(n179), .A2(n187), .B1(n180), .B2(n187), .ZN(N241) );
  XOR3D4 U58 ( .A1(n199), .A2(wo_2[1]), .A3(n126), .Z(n180) );
  OAI22D2 U60 ( .A1(n208), .A2(n113), .B1(n173), .B2(n174), .ZN(N247) );
  XOR3D2 U62 ( .A1(wo_3[7]), .A2(wo_2[7]), .A3(n114), .Z(n113) );
  XOR3D4 U64 ( .A1(wo_3[8]), .A2(wo_2[8]), .A3(n112), .Z(n111) );
  CKND0 U66 ( .I(wo_3[1]), .ZN(n199) );
  XNR2D2 U67 ( .A1(subword[25]), .A2(n193), .ZN(n14) );
  XOR3D4 U68 ( .A1(wo_3[12]), .A2(wo_2[12]), .A3(n104), .Z(n163) );
  XOR3D4 U70 ( .A1(wo_3[14]), .A2(wo_2[14]), .A3(n100), .Z(n99) );
  XOR3D4 U72 ( .A1(wo_3[3]), .A2(wo_2[3]), .A3(n122), .Z(n121) );
  INVD3 U73 ( .I(n207), .ZN(wo_3[24]) );
  INVD1 U74 ( .I(wo_0[1]), .ZN(n165) );
  INVD1 U75 ( .I(n196), .ZN(n181) );
  INVD1 U76 ( .I(key[9]), .ZN(n185) );
  INVD1 U78 ( .I(n196), .ZN(n186) );
  INVD1 U79 ( .I(key[25]), .ZN(n183) );
  INVD1 U80 ( .I(key[7]), .ZN(n173) );
  INVD1 U82 ( .I(n196), .ZN(n174) );
  INVD1 U83 ( .I(key[17]), .ZN(n175) );
  INVD1 U84 ( .I(wo_0[19]), .ZN(n164) );
  INVD1 U86 ( .I(wo_0[9]), .ZN(n166) );
  BUFFD2 U88 ( .I(kld), .Z(n208) );
  INVD2 U89 ( .I(n203), .ZN(wo_3[16]) );
  XOR3D1 U90 ( .A1(wo_3[30]), .A2(wo_2[30]), .A3(n68), .Z(n67) );
  INVD1 U91 ( .I(key[27]), .ZN(n170) );
  XOR3D1 U92 ( .A1(wo_3[26]), .A2(wo_2[26]), .A3(n76), .Z(n75) );
  XOR3D1 U94 ( .A1(wo_3[6]), .A2(wo_2[6]), .A3(n116), .Z(n115) );
  INVD1 U95 ( .I(key[20]), .ZN(n167) );
  INVD1 U96 ( .I(n196), .ZN(n161) );
  XOR3D1 U98 ( .A1(wo_3[29]), .A2(wo_2[29]), .A3(n70), .Z(n69) );
  XOR3D1 U100 ( .A1(wo_3[0]), .A2(wo_2[0]), .A3(n128), .Z(n127) );
  INVD1 U102 ( .I(key[1]), .ZN(n179) );
  INVD1 U104 ( .I(key[11]), .ZN(n172) );
  INVD1 U105 ( .I(key[23]), .ZN(n176) );
  MOAI22D1 U106 ( .A1(n167), .A2(n184), .B1(n161), .B2(n162), .ZN(N260) );
  XNR3D1 U107 ( .A1(wo_3[20]), .A2(wo_2[20]), .A3(n88), .ZN(n162) );
  INVD1 U108 ( .I(n208), .ZN(n169) );
  INVD1 U110 ( .I(n208), .ZN(n187) );
  CKXOR2D1 U111 ( .A1(n106), .A2(wo_2[11]), .Z(n149) );
  XNR3D1 U112 ( .A1(wo_3[27]), .A2(wo_2[27]), .A3(n74), .ZN(n171) );
  MOAI22D1 U114 ( .A1(n196), .A2(n163), .B1(key[12]), .B2(n195), .ZN(N252) );
  XNR2D1 U115 ( .A1(subword[19]), .A2(n164), .ZN(n26) );
  XNR2D1 U116 ( .A1(n165), .A2(subword[1]), .ZN(n62) );
  CKXOR2D1 U118 ( .A1(n90), .A2(wo_2[19]), .Z(n141) );
  MOAI22D0 U120 ( .A1(n208), .A2(n90), .B1(key[83]), .B2(n196), .ZN(N127) );
  XNR2D1 U121 ( .A1(n166), .A2(subword[9]), .ZN(n46) );
  CKND0 U122 ( .I(n24), .ZN(n23) );
  XNR2D4 U124 ( .A1(n62), .A2(wo_1[1]), .ZN(n126) );
  XNR2D1 U126 ( .A1(wo_1[20]), .A2(n24), .ZN(n168) );
  CKXOR2D0 U127 ( .A1(n125), .A2(wo_2[17]), .Z(n143) );
  ND2D0 U128 ( .A1(subword[28]), .A2(n192), .ZN(n190) );
  MOAI22D0 U130 ( .A1(n208), .A2(n74), .B1(key[91]), .B2(n195), .ZN(N135) );
  XNR3D4 U144 ( .A1(wo_1[27]), .A2(rcon[27]), .A3(n10), .ZN(n74) );
  MOAI22D0 U156 ( .A1(n208), .A2(n70), .B1(key[93]), .B2(n195), .ZN(N137) );
  XNR3D4 U160 ( .A1(wo_1[29]), .A2(rcon[29]), .A3(n6), .ZN(n70) );
  MOAI22D1 U170 ( .A1(n170), .A2(n181), .B1(n169), .B2(n171), .ZN(N267) );
  OAI22D2 U172 ( .A1(n105), .A2(n208), .B1(n172), .B2(n188), .ZN(N251) );
  CKND2 U188 ( .I(n187), .ZN(n196) );
  INVD1 U192 ( .I(n194), .ZN(n177) );
  INVD1 U196 ( .I(n194), .ZN(n184) );
  INVD1 U199 ( .I(n194), .ZN(n188) );
  CKND1 U201 ( .I(n169), .ZN(n194) );
  XOR3D1 U202 ( .A1(wo_3[21]), .A2(wo_2[21]), .A3(n86), .Z(n85) );
  XOR3D1 U205 ( .A1(wo_3[2]), .A2(wo_2[2]), .A3(n124), .Z(n123) );
  OAI22D2 U206 ( .A1(n208), .A2(n93), .B1(n175), .B2(n187), .ZN(N257) );
  OAI22D2 U207 ( .A1(n208), .A2(n81), .B1(n176), .B2(n177), .ZN(N263) );
  XNR3D1 U208 ( .A1(wo_3[25]), .A2(wo_2[25]), .A3(n78), .ZN(n178) );
  XNR3D4 U211 ( .A1(wo_1[25]), .A2(rcon[25]), .A3(n14), .ZN(n78) );
  MOAI22D1 U213 ( .A1(n183), .A2(n184), .B1(n187), .B2(n178), .ZN(N265) );
  CKXOR2D1 U214 ( .A1(n78), .A2(wo_2[25]), .Z(n135) );
  XOR3D4 U215 ( .A1(wo_3[23]), .A2(wo_2[23]), .A3(n82), .Z(n81) );
  XOR3D4 U217 ( .A1(wo_3[18]), .A2(wo_2[18]), .A3(n92), .Z(n91) );
  AO22D1 U220 ( .A1(n181), .A2(n182), .B1(key[31]), .B2(n194), .Z(N271) );
  XNR3D1 U223 ( .A1(wo_3[31]), .A2(wo_2[31]), .A3(n66), .ZN(n182) );
  INVD4 U226 ( .I(n205), .ZN(wo_3[19]) );
  CKND2 U228 ( .I(n210), .ZN(n205) );
  XOR3D4 U229 ( .A1(wo_3[10]), .A2(wo_2[10]), .A3(n108), .Z(n107) );
  XOR3D4 U231 ( .A1(wo_3[5]), .A2(wo_2[5]), .A3(n118), .Z(n117) );
  XNR3D4 U232 ( .A1(wo_1[28]), .A2(rcon[28]), .A3(n8), .ZN(n72) );
  ND2D2 U233 ( .A1(n190), .A2(n191), .ZN(n8) );
  OAI22D2 U235 ( .A1(n109), .A2(n208), .B1(n185), .B2(n186), .ZN(N249) );
  XOR3D4 U237 ( .A1(wo_3[16]), .A2(wo_2[16]), .A3(n96), .Z(n95) );
  XOR3D4 U238 ( .A1(wo_3[11]), .A2(wo_2[11]), .A3(n106), .Z(n105) );
  XOR3D4 U241 ( .A1(wo_3[17]), .A2(wo_2[17]), .A3(n94), .Z(n93) );
  XOR3D4 U244 ( .A1(wo_3[9]), .A2(wo_2[9]), .A3(n110), .Z(n109) );
  CKND2 U247 ( .I(n198), .ZN(wo_3[0]) );
  CKND1 U250 ( .I(subword[28]), .ZN(n189) );
  CKND0 U252 ( .I(n38), .ZN(n37) );
  IND2D1 U253 ( .A1(n192), .B1(n189), .ZN(n191) );
  CKND0 U255 ( .I(n62), .ZN(n61) );
  CKND0 U256 ( .I(n52), .ZN(n51) );
  CKND0 U259 ( .I(n34), .ZN(n33) );
  CKND0 U261 ( .I(n58), .ZN(n57) );
  CKND0 U262 ( .I(n46), .ZN(n45) );
  CKND0 U263 ( .I(n44), .ZN(n43) );
  CKND0 U265 ( .I(n50), .ZN(n49) );
  CKND0 U268 ( .I(n54), .ZN(n53) );
  CKND0 U271 ( .I(n36), .ZN(n35) );
  CKND0 U274 ( .I(n26), .ZN(n25) );
  XOR3D0 U277 ( .A1(wo_3[22]), .A2(wo_2[22]), .A3(n84), .Z(n83) );
  CKND0 U279 ( .I(n64), .ZN(n63) );
  CKND0 U280 ( .I(n20), .ZN(n19) );
  CKND0 U283 ( .I(n22), .ZN(n21) );
  MOAI22D0 U285 ( .A1(n208), .A2(n168), .B1(key[84]), .B2(n194), .ZN(N128) );
  CKND0 U286 ( .I(n32), .ZN(n31) );
  CKND0 U287 ( .I(n42), .ZN(n41) );
  CKND0 U289 ( .I(n18), .ZN(n17) );
  CKND0 U291 ( .I(n56), .ZN(n55) );
  CKND0 U292 ( .I(n60), .ZN(n59) );
  CKND0 U293 ( .I(n28), .ZN(n27) );
  CKND0 U294 ( .I(n48), .ZN(n47) );
  CKND2 U295 ( .I(n201), .ZN(wo_3[8]) );
  INVD1 U296 ( .I(n169), .ZN(n195) );
  INVD1 U297 ( .I(wo_0[25]), .ZN(n193) );
  XOR3D1 U298 ( .A1(wo_3[15]), .A2(wo_2[15]), .A3(n98), .Z(n97) );
  XNR3D1 U299 ( .A1(wo_1[26]), .A2(rcon[26]), .A3(n12), .ZN(n76) );
  XNR3D1 U300 ( .A1(wo_1[24]), .A2(rcon[24]), .A3(n16), .ZN(n80) );
  XNR3D1 U301 ( .A1(wo_1[30]), .A2(rcon[30]), .A3(n4), .ZN(n68) );
  XNR3D1 U302 ( .A1(wo_1[31]), .A2(rcon[31]), .A3(n2), .ZN(n66) );
  INVD1 U303 ( .I(n209), .ZN(n207) );
  INVD1 U304 ( .I(n212), .ZN(n201) );
  INVD1 U305 ( .I(n211), .ZN(n203) );
  INVD1 U306 ( .I(n213), .ZN(n198) );
  MOAI22D0 U307 ( .A1(n208), .A2(n78), .B1(key[89]), .B2(n195), .ZN(N133) );
  CKND0 U308 ( .I(n30), .ZN(n29) );
  MOAI22D0 U309 ( .A1(n208), .A2(n106), .B1(key[75]), .B2(n195), .ZN(N119) );
  CKND0 U310 ( .I(n40), .ZN(n39) );
  MOAI22D0 U311 ( .A1(n208), .A2(n110), .B1(key[73]), .B2(n195), .ZN(N117) );
  MOAI22D0 U312 ( .A1(n208), .A2(n126), .B1(key[65]), .B2(n195), .ZN(N109) );
  MOAI22D0 U313 ( .A1(n208), .A2(n125), .B1(key[81]), .B2(n195), .ZN(N125) );
  MOAI22D0 U314 ( .A1(n208), .A2(n104), .B1(key[76]), .B2(n196), .ZN(N120) );
  INVD1 U315 ( .I(wo_0[28]), .ZN(n192) );
  XNR2D1 U316 ( .A1(wo_1[0]), .A2(n64), .ZN(n128) );
  XNR2D1 U317 ( .A1(wo_1[2]), .A2(n60), .ZN(n124) );
  XNR2D1 U318 ( .A1(wo_1[3]), .A2(n58), .ZN(n122) );
  XNR2D1 U319 ( .A1(wo_1[4]), .A2(n56), .ZN(n120) );
  XNR2D1 U320 ( .A1(wo_1[5]), .A2(n54), .ZN(n118) );
  XNR2D1 U321 ( .A1(wo_1[6]), .A2(n52), .ZN(n116) );
  XNR2D1 U322 ( .A1(wo_1[7]), .A2(n50), .ZN(n114) );
  XNR2D1 U323 ( .A1(wo_1[8]), .A2(n48), .ZN(n112) );
  XNR2D1 U324 ( .A1(n46), .A2(wo_1[9]), .ZN(n110) );
  XNR2D1 U325 ( .A1(wo_1[10]), .A2(n44), .ZN(n108) );
  XNR2D1 U326 ( .A1(wo_1[11]), .A2(n42), .ZN(n106) );
  XNR2D1 U327 ( .A1(wo_1[12]), .A2(n40), .ZN(n104) );
  XNR2D1 U328 ( .A1(wo_1[13]), .A2(n38), .ZN(n102) );
  XNR2D1 U329 ( .A1(wo_1[14]), .A2(n36), .ZN(n100) );
  XNR2D1 U330 ( .A1(wo_1[15]), .A2(n34), .ZN(n98) );
  XNR2D1 U331 ( .A1(wo_1[16]), .A2(n32), .ZN(n96) );
  XNR2D1 U332 ( .A1(wo_1[17]), .A2(n30), .ZN(n94) );
  XNR2D1 U333 ( .A1(wo_1[18]), .A2(n28), .ZN(n92) );
  XNR2D1 U334 ( .A1(wo_1[19]), .A2(n26), .ZN(n90) );
  XNR2D1 U335 ( .A1(wo_1[20]), .A2(n24), .ZN(n88) );
  XNR2D1 U336 ( .A1(wo_1[21]), .A2(n22), .ZN(n86) );
  XNR2D1 U337 ( .A1(wo_1[22]), .A2(n20), .ZN(n84) );
  XNR2D1 U338 ( .A1(wo_1[23]), .A2(n18), .ZN(n82) );
endmodule


module aes_sbox_0 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n50, n51, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n66, n67, n69, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n117,
         n118, n119, n120, n121, n122, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n293, n297, n298, n312, n315, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n406, n407,
         n408, n409, n410, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, net7393, net7391, net7389, net7419, net7422,
         net7425, net7427, net7429, net7431, net7435, net8311, net8553,
         net8772, net9112, net12708, net12814, net12847, net12846, n52, n323,
         n322, n321, n320, n319, n318, n317, n316, n314, n313, n311, n310,
         n309, n308, n307, n306, n305, n304, n301, n300, n299, n296, n295,
         n294, n292, n291, n290, n289, n288, n20, n9, n49, n65, n68, n70, n116,
         n123, n142, n192, n287, n302, n303, n404, n405, n411, n424, n425,
         n426, n427, n428;

  AN2XD1 U28 ( .A1(n147), .A2(n148), .Z(n143) );
  OA21D1 U35 ( .A1(n163), .A2(n164), .B(n165), .Z(n158) );
  OR3D1 U88 ( .A1(n196), .A2(n53), .A3(net7393), .Z(n235) );
  OA21D1 U101 ( .A1(n182), .A2(net7422), .B(n254), .Z(n250) );
  OR4D1 U199 ( .A1(n211), .A2(n293), .A3(n349), .A4(n350), .Z(n347) );
  AN2XD1 U215 ( .A1(n348), .A2(n55), .Z(n349) );
  AO31D1 U286 ( .A1(n62), .A2(n5), .A3(n185), .B(n149), .Z(n409) );
  AO21D1 U297 ( .A1(n9), .A2(n29), .B(n132), .Z(n410) );
  AOI221D1 U1 ( .A1(n9), .A2(n184), .B1(n185), .B2(n59), .C(n186), .ZN(n183)
         );
  OAI22D0 U2 ( .A1(n401), .A2(n157), .B1(n402), .B2(n106), .ZN(n400) );
  OAI211D1 U3 ( .A1(net7427), .A2(n84), .B(n242), .C(n117), .ZN(n333) );
  OAI222D0 U4 ( .A1(n161), .A2(n135), .B1(net7435), .B2(n331), .C1(n81), .C2(
        n92), .ZN(n330) );
  ND4D2 U5 ( .A1(n389), .A2(n390), .A3(n391), .A4(n392), .ZN(d[7]) );
  INR2XD0 U6 ( .A1(n116), .B1(n199), .ZN(n188) );
  OAI222D1 U7 ( .A1(n54), .A2(n237), .B1(n315), .B2(n335), .C1(n336), .C2(n86), 
        .ZN(n329) );
  NR4D0 U8 ( .A1(n337), .A2(n338), .A3(n339), .A4(n274), .ZN(n336) );
  AOI22D1 U9 ( .A1(n34), .A2(n48), .B1(n59), .B2(n37), .ZN(n311) );
  INVD2 U10 ( .I(n226), .ZN(n48) );
  ND2D0 U11 ( .A1(n48), .A2(n45), .ZN(n265) );
  AOI221D2 U12 ( .A1(n64), .A2(n6), .B1(n55), .B2(n27), .C(n410), .ZN(n406) );
  AOI221D2 U13 ( .A1(n408), .A2(n57), .B1(n12), .B2(n47), .C(n409), .ZN(n407)
         );
  OAI221D1 U14 ( .A1(n128), .A2(n135), .B1(n162), .B2(n122), .C(n275), .ZN(
        n267) );
  INVD2 U15 ( .I(n91), .ZN(n68) );
  INVD2 U16 ( .I(n148), .ZN(n71) );
  OAI222D1 U17 ( .A1(net9112), .A2(n335), .B1(n381), .B2(n115), .C1(n382), 
        .C2(n111), .ZN(n377) );
  AOI221D1 U18 ( .A1(n67), .A2(n179), .B1(n31), .B2(net8311), .C(n180), .ZN(
        n178) );
  INVD2 U19 ( .I(n109), .ZN(n5) );
  AOI221D1 U20 ( .A1(n19), .A2(n412), .B1(n413), .B2(net7422), .C(n414), .ZN(
        n389) );
  AOI221D1 U21 ( .A1(n398), .A2(net7391), .B1(n43), .B2(n399), .C(n400), .ZN(
        n391) );
  OAI222D1 U22 ( .A1(n340), .A2(n91), .B1(net9112), .B2(n243), .C1(n341), .C2(
        n148), .ZN(n328) );
  ND2D1 U23 ( .A1(a[6]), .A2(n25), .ZN(n86) );
  INVD2 U24 ( .I(net12846), .ZN(net12847) );
  CKND1 U25 ( .I(net7389), .ZN(net12846) );
  INVD3 U26 ( .I(net7431), .ZN(n51) );
  ND2D0 U27 ( .A1(net7422), .A2(net7419), .ZN(n103) );
  CKND3 U29 ( .I(n49), .ZN(net12708) );
  CKND2D2 U30 ( .A1(net7427), .A2(n45), .ZN(n101) );
  INVD1 U31 ( .I(n94), .ZN(n53) );
  BUFFD4 U32 ( .I(a[4]), .Z(net7429) );
  CKND2D1 U33 ( .A1(net7389), .A2(a[2]), .ZN(n119) );
  INVD2 U34 ( .I(n81), .ZN(n62) );
  CKND2D1 U36 ( .A1(net7431), .A2(n45), .ZN(n117) );
  INVD1 U37 ( .I(a[1]), .ZN(net7393) );
  CKND2D1 U38 ( .A1(n51), .A2(n45), .ZN(n111) );
  INVD1 U39 ( .I(n98), .ZN(n31) );
  INVD1 U40 ( .I(n114), .ZN(n64) );
  ND2D3 U41 ( .A1(net7393), .A2(net7419), .ZN(n114) );
  ND2D2 U42 ( .A1(net7431), .A2(a[2]), .ZN(n226) );
  ND2D1 U43 ( .A1(net7389), .A2(net7435), .ZN(n148) );
  OAI221D0 U44 ( .A1(n253), .A2(n101), .B1(net12708), .B2(n106), .C(n375), 
        .ZN(n372) );
  IAO21D1 U45 ( .A1(n94), .A2(n146), .B(n302), .ZN(n287) );
  INVD1 U46 ( .I(net12847), .ZN(n303) );
  INVD2 U47 ( .I(n162), .ZN(n16) );
  INVD1 U48 ( .I(n190), .ZN(n46) );
  INVD1 U49 ( .I(n191), .ZN(n3) );
  INVD1 U50 ( .I(n101), .ZN(n32) );
  INVD1 U51 ( .I(n203), .ZN(n59) );
  ND4D1 U52 ( .A1(n150), .A2(n151), .A3(n152), .A4(n153), .ZN(d[1]) );
  AOI221D0 U53 ( .A1(n8), .A2(n71), .B1(n175), .B2(n5), .C(n176), .ZN(n151) );
  AOI221D1 U54 ( .A1(n14), .A2(n55), .B1(n174), .B2(n62), .C(n187), .ZN(n150)
         );
  AOI221D0 U55 ( .A1(n22), .A2(n214), .B1(n19), .B2(n215), .C(n216), .ZN(n207)
         );
  AOI221D0 U56 ( .A1(n52), .A2(n297), .B1(n298), .B2(n42), .C(n299), .ZN(n289)
         );
  ND4D1 U57 ( .A1(n361), .A2(n362), .A3(n363), .A4(n364), .ZN(d[6]) );
  NR3D0 U58 ( .A1(n302), .A2(n200), .A3(n192), .ZN(n116) );
  INVD1 U59 ( .I(n198), .ZN(n192) );
  INVD1 U60 ( .I(n232), .ZN(n10) );
  ND2D2 U61 ( .A1(net7425), .A2(a[6]), .ZN(n162) );
  ND2D1 U62 ( .A1(n45), .A2(n37), .ZN(n97) );
  ND2D2 U63 ( .A1(net7389), .A2(net7419), .ZN(n81) );
  ND2D1 U64 ( .A1(net7419), .A2(n51), .ZN(n182) );
  ND2D1 U65 ( .A1(n12), .A2(net7422), .ZN(n231) );
  AOI21D1 U66 ( .A1(n65), .A2(n68), .B(n70), .ZN(net8553) );
  OA222D1 U67 ( .A1(n406), .A2(n117), .B1(n181), .B2(n355), .C1(n407), .C2(
        net7422), .Z(n427) );
  INVD1 U68 ( .I(n287), .ZN(n70) );
  OAI21D1 U69 ( .A1(n142), .A2(n302), .B(n303), .ZN(n123) );
  INVD1 U70 ( .I(n136), .ZN(n12) );
  INVD1 U71 ( .I(n182), .ZN(n50) );
  OAI222D0 U72 ( .A1(n114), .A2(n262), .B1(n263), .B2(net7419), .C1(n264), 
        .C2(n191), .ZN(n261) );
  MAOI22D1 U73 ( .A1(n7), .A2(n51), .B1(n242), .B2(n93), .ZN(n356) );
  ND2D1 U74 ( .A1(n425), .A2(n426), .ZN(n204) );
  OR2D1 U75 ( .A1(n144), .A2(n114), .Z(n425) );
  OA221D1 U76 ( .A1(n182), .A2(n193), .B1(n194), .B2(n81), .C(n195), .Z(n428)
         );
  AOI211XD1 U77 ( .A1(n35), .A2(n281), .B(n282), .C(n283), .ZN(n280) );
  OAI211D0 U78 ( .A1(n164), .A2(n190), .B(n320), .C(n321), .ZN(n304) );
  INVD1 U79 ( .I(n9), .ZN(net12814) );
  CKND3 U80 ( .I(a[1]), .ZN(net7391) );
  INVD2 U81 ( .I(net7391), .ZN(net7389) );
  CKAN2D1 U82 ( .A1(net7435), .A2(net7391), .Z(n9) );
  AN2XD1 U83 ( .A1(net7429), .A2(net7431), .Z(n49) );
  ND2D2 U84 ( .A1(net12847), .A2(net7422), .ZN(n128) );
  OR2D1 U85 ( .A1(n3), .A2(n17), .Z(n65) );
  INVD0 U86 ( .I(n312), .ZN(n63) );
  OAI221D1 U87 ( .A1(n300), .A2(n157), .B1(n301), .B2(net12814), .C(n123), 
        .ZN(n299) );
  IND2D1 U89 ( .A1(n232), .B1(n53), .ZN(n404) );
  ND2D1 U90 ( .A1(n16), .A2(n32), .ZN(n232) );
  INVD1 U91 ( .I(n404), .ZN(n302) );
  ND2D3 U92 ( .A1(net7422), .A2(net7391), .ZN(n122) );
  NR2D1 U93 ( .A1(n164), .A2(n122), .ZN(n132) );
  AOI22D1 U94 ( .A1(n62), .A2(n28), .B1(n53), .B2(n45), .ZN(n95) );
  ND2D1 U95 ( .A1(a[2]), .A2(net7393), .ZN(n203) );
  AOI221D1 U96 ( .A1(n166), .A2(n6), .B1(n48), .B2(n167), .C(n168), .ZN(n152)
         );
  OAI221D0 U97 ( .A1(n419), .A2(n226), .B1(n94), .B2(n135), .C(n420), .ZN(n413) );
  INR2D1 U98 ( .A1(n48), .B1(n191), .ZN(n142) );
  OAI33D0 U99 ( .A1(n226), .A2(net7425), .A3(n97), .B1(n164), .B2(net7419), 
        .B3(net12708), .ZN(n334) );
  ND2D1 U100 ( .A1(n64), .A2(net7435), .ZN(n312) );
  BUFFD6 U102 ( .I(a[7]), .Z(net7425) );
  AO221D0 U103 ( .A1(n64), .A2(n31), .B1(n67), .B2(n68), .C(n166), .Z(n215) );
  OAI22D1 U104 ( .A1(n101), .A2(n91), .B1(net12847), .B2(n102), .ZN(n100) );
  AOI221D1 U105 ( .A1(n29), .A2(n71), .B1(n276), .B2(net7391), .C(n132), .ZN(
        n275) );
  OAI21D0 U106 ( .A1(n115), .A2(n257), .B(n146), .ZN(n276) );
  OAI222D1 U107 ( .A1(n121), .A2(n148), .B1(n97), .B2(n286), .C1(net12708), 
        .C2(n106), .ZN(n282) );
  ND2D1 U108 ( .A1(n53), .A2(net12847), .ZN(n286) );
  AOI221D2 U109 ( .A1(n63), .A2(n14), .B1(n71), .B2(n1), .C(n277), .ZN(n244)
         );
  NR4D1 U110 ( .A1(n77), .A2(n78), .A3(n79), .A4(n80), .ZN(n76) );
  INVD2 U111 ( .I(n257), .ZN(n34) );
  ND2D2 U112 ( .A1(net7429), .A2(n37), .ZN(n257) );
  AOI221D2 U113 ( .A1(n42), .A2(n69), .B1(n33), .B2(n57), .C(n310), .ZN(n309)
         );
  OAI222D2 U114 ( .A1(net8772), .A2(n98), .B1(net7435), .B2(n311), .C1(
        net12708), .C2(n312), .ZN(n310) );
  ND2D1 U115 ( .A1(a[6]), .A2(n37), .ZN(n93) );
  ND2D1 U116 ( .A1(net7425), .A2(n37), .ZN(n139) );
  AOI222D1 U117 ( .A1(n57), .A2(n34), .B1(n59), .B2(n386), .C1(n63), .C2(n31), 
        .ZN(n381) );
  ND4D2 U118 ( .A1(n244), .A2(n245), .A3(n246), .A4(n247), .ZN(d[3]) );
  AOI221D1 U119 ( .A1(n19), .A2(n259), .B1(n260), .B2(net7422), .C(n261), .ZN(
        n246) );
  NR4D1 U120 ( .A1(n327), .A2(n328), .A3(n329), .A4(n330), .ZN(n326) );
  AOI221D1 U121 ( .A1(net7435), .A2(n304), .B1(n22), .B2(n305), .C(n306), .ZN(
        n288) );
  OAI222D1 U122 ( .A1(n307), .A2(n109), .B1(n308), .B2(n182), .C1(n115), .C2(
        n309), .ZN(n306) );
  OAI222D1 U123 ( .A1(net7435), .A2(n188), .B1(n115), .B2(n189), .C1(n190), 
        .C2(n191), .ZN(n187) );
  ND3D0 U124 ( .A1(n48), .A2(n197), .A3(n19), .ZN(n107) );
  CKND2D1 U125 ( .A1(n19), .A2(n32), .ZN(n83) );
  INVD2 U126 ( .I(n115), .ZN(n19) );
  OAI221D1 U127 ( .A1(n201), .A2(n190), .B1(n202), .B2(net8772), .C(n18), .ZN(
        n199) );
  INVD0 U128 ( .I(n122), .ZN(n69) );
  OAI32D1 U129 ( .A1(n284), .A2(n122), .A3(n181), .B1(n285), .B2(n101), .ZN(
        n283) );
  AOI221D1 U130 ( .A1(n68), .A2(n267), .B1(n22), .B2(n268), .C(n269), .ZN(n245) );
  OAI222D1 U131 ( .A1(n226), .A2(n233), .B1(n278), .B2(n279), .C1(n280), .C2(
        n109), .ZN(n277) );
  IND4D1 U132 ( .A1(n424), .B1(n288), .B2(n289), .B3(n290), .ZN(d[4]) );
  ND2D2 U133 ( .A1(net7431), .A2(n37), .ZN(n120) );
  AOI221D1 U134 ( .A1(n4), .A2(net7422), .B1(n12), .B2(n57), .C(n236), .ZN(
        n205) );
  AOI211XD0 U135 ( .A1(n1), .A2(n56), .B(n388), .C(n204), .ZN(n361) );
  OAI222D0 U136 ( .A1(n226), .A2(n144), .B1(n278), .B2(n135), .C1(n232), .C2(
        net8772), .ZN(n388) );
  AOI211XD0 U137 ( .A1(n23), .A2(n56), .B(n383), .C(n384), .ZN(n382) );
  ND2D1 U138 ( .A1(net7431), .A2(net7393), .ZN(n190) );
  CKND2D2 U139 ( .A1(n37), .A2(n30), .ZN(n212) );
  OA221D1 U140 ( .A1(n120), .A2(n128), .B1(n111), .B2(net8772), .C(n428), .Z(
        n189) );
  OAI222D1 U141 ( .A1(n83), .A2(n286), .B1(n91), .B2(n231), .C1(n374), .C2(
        n103), .ZN(n373) );
  AOI211D0 U142 ( .A1(n90), .A2(n212), .B(n284), .C(net12814), .ZN(n395) );
  OAI33D0 U143 ( .A1(n111), .A2(net7419), .A3(n139), .B1(n212), .B2(net12847), 
        .B3(n213), .ZN(n209) );
  OAI221D1 U144 ( .A1(n258), .A2(n284), .B1(net7431), .B2(n92), .C(n165), .ZN(
        n342) );
  INVD6 U145 ( .I(net7427), .ZN(n37) );
  ND2D1 U146 ( .A1(n22), .A2(n197), .ZN(n135) );
  AOI221D1 U147 ( .A1(n3), .A2(net7391), .B1(n21), .B2(n148), .C(n343), .ZN(
        n340) );
  AO221D0 U148 ( .A1(n53), .A2(n20), .B1(n12), .B2(n47), .C(n323), .Z(n424) );
  CKND0 U149 ( .I(n146), .ZN(n20) );
  ND2D1 U150 ( .A1(n22), .A2(n36), .ZN(n146) );
  INVD1 U151 ( .I(n84), .ZN(n47) );
  OAI222D0 U152 ( .A1(net9112), .A2(n271), .B1(n135), .B2(n190), .C1(n232), 
        .C2(n106), .ZN(n323) );
  ND2D1 U153 ( .A1(net7435), .A2(n66), .ZN(net9112) );
  CKND2D0 U154 ( .A1(n35), .A2(n16), .ZN(n271) );
  ND2D1 U155 ( .A1(net7435), .A2(a[2]), .ZN(n106) );
  BUFFD6 U156 ( .I(a[0]), .Z(net7435) );
  ND2D1 U157 ( .A1(net7427), .A2(net7425), .ZN(n164) );
  AOI32D0 U158 ( .A1(net7429), .A2(n25), .A3(n68), .B1(n48), .B2(n322), .ZN(
        n320) );
  INVD4 U159 ( .I(net7425), .ZN(n25) );
  OAI22D0 U160 ( .A1(a[6]), .A2(net7429), .B1(net7427), .B2(n109), .ZN(n322)
         );
  BUFFD4 U161 ( .I(a[5]), .Z(net7427) );
  ND2D3 U162 ( .A1(net7425), .A2(n30), .ZN(n109) );
  AOI22D0 U163 ( .A1(n3), .A2(n62), .B1(n47), .B2(n17), .ZN(n321) );
  INVD1 U164 ( .I(n83), .ZN(n17) );
  INVD1 U165 ( .I(n86), .ZN(n22) );
  OAI211D1 U166 ( .A1(n316), .A2(n148), .B(n317), .C(n318), .ZN(n305) );
  ND2D1 U167 ( .A1(net7419), .A2(n45), .ZN(n316) );
  AOI32D0 U168 ( .A1(n64), .A2(net7422), .A3(n31), .B1(n67), .B2(n319), .ZN(
        n317) );
  BUFFD8 U169 ( .I(n72), .Z(net7422) );
  INVD1 U170 ( .I(n128), .ZN(n67) );
  CKND2D0 U171 ( .A1(net12708), .A2(n121), .ZN(n319) );
  CKND2D0 U172 ( .A1(a[2]), .A2(net7427), .ZN(n121) );
  AOI222D0 U173 ( .A1(n57), .A2(n40), .B1(n42), .B2(net8311), .C1(n33), .C2(
        n59), .ZN(n318) );
  INVD1 U174 ( .I(n119), .ZN(n57) );
  INVD1 U175 ( .I(n157), .ZN(n40) );
  INVD2 U176 ( .I(n117), .ZN(n42) );
  AN2XD1 U177 ( .A1(net7435), .A2(n66), .Z(net8311) );
  CKND1 U178 ( .I(n181), .ZN(n33) );
  AOI221D0 U179 ( .A1(n61), .A2(n31), .B1(n36), .B2(n314), .C(n166), .ZN(n307)
         );
  INVD1 U180 ( .I(n315), .ZN(n61) );
  INVD1 U181 ( .I(n97), .ZN(n36) );
  CKND2D0 U182 ( .A1(n84), .A2(n315), .ZN(n314) );
  ND2D2 U183 ( .A1(net12847), .A2(net7431), .ZN(n84) );
  ND2D2 U184 ( .A1(n62), .A2(net7422), .ZN(n315) );
  NR2D1 U185 ( .A1(n242), .A2(n148), .ZN(n166) );
  NR3D0 U186 ( .A1(n405), .A2(n411), .A3(n313), .ZN(n308) );
  CKAN2D1 U187 ( .A1(n174), .A2(n122), .Z(n405) );
  NR2D0 U188 ( .A1(n115), .A2(n97), .ZN(n174) );
  CKAN2D1 U189 ( .A1(net12847), .A2(n10), .Z(n411) );
  OAI31D0 U190 ( .A1(n162), .A2(net7427), .A3(net12847), .B(n231), .ZN(n313)
         );
  BUFFD1 U191 ( .I(n203), .Z(net8772) );
  ND2D1 U192 ( .A1(net7427), .A2(n51), .ZN(n98) );
  ND2D1 U193 ( .A1(n30), .A2(n25), .ZN(n115) );
  INVD1 U194 ( .I(n286), .ZN(n52) );
  CKND2D0 U195 ( .A1(n93), .A2(n139), .ZN(n297) );
  NR2D1 U196 ( .A1(n360), .A2(net8772), .ZN(n298) );
  AOI22D0 U197 ( .A1(n56), .A2(n6), .B1(n64), .B2(n27), .ZN(n300) );
  INVD1 U198 ( .I(n161), .ZN(n56) );
  INVD1 U200 ( .I(n139), .ZN(n6) );
  INVD1 U201 ( .I(n93), .ZN(n27) );
  ND2D2 U202 ( .A1(net7429), .A2(n51), .ZN(n157) );
  AOI21D1 U203 ( .A1(n44), .A2(n2), .B(n15), .ZN(n301) );
  INVD1 U204 ( .I(n316), .ZN(n44) );
  CKND0 U205 ( .I(n164), .ZN(n2) );
  INVD1 U206 ( .I(n262), .ZN(n15) );
  NR4D0 U207 ( .A1(n291), .A2(n292), .A3(n293), .A4(n127), .ZN(n290) );
  OAI222D0 U208 ( .A1(n294), .A2(n92), .B1(n83), .B2(n295), .C1(n296), .C2(n90), .ZN(n291) );
  NR2D1 U209 ( .A1(n61), .A2(n58), .ZN(n294) );
  INVD1 U210 ( .I(n138), .ZN(n58) );
  ND2D0 U211 ( .A1(n197), .A2(n5), .ZN(n92) );
  CKND2D0 U212 ( .A1(n148), .A2(n51), .ZN(n295) );
  AOI22D0 U213 ( .A1(n39), .A2(n69), .B1(n41), .B2(a[2]), .ZN(n296) );
  INVD1 U214 ( .I(n163), .ZN(n39) );
  INVD1 U216 ( .I(net12708), .ZN(n41) );
  CKND2D0 U217 ( .A1(net7427), .A2(a[6]), .ZN(n90) );
  NR4D0 U218 ( .A1(net7435), .A2(n30), .A3(n97), .A4(n91), .ZN(n292) );
  INVD2 U219 ( .I(a[6]), .ZN(n30) );
  ND2D0 U220 ( .A1(a[2]), .A2(n51), .ZN(n91) );
  NR3D0 U221 ( .A1(n148), .A2(n45), .A3(n137), .ZN(n293) );
  NR4D0 U222 ( .A1(n97), .A2(n109), .A3(net8772), .A4(net7431), .ZN(n127) );
  INVD6 U223 ( .I(net7429), .ZN(n45) );
  NR2D2 U224 ( .A1(n45), .A2(n37), .ZN(n197) );
  ND4D1 U225 ( .A1(n205), .A2(n206), .A3(n207), .A4(n208), .ZN(d[2]) );
  OAI31D0 U226 ( .A1(n119), .A2(n90), .A3(n117), .B(n255), .ZN(n248) );
  AOI221D1 U227 ( .A1(n42), .A2(n5), .B1(n53), .B2(n32), .C(n342), .ZN(n341)
         );
  OAI33D0 U228 ( .A1(n114), .A2(n115), .A3(net12708), .B1(n93), .B2(net7419), 
        .B3(n117), .ZN(n113) );
  AOI221D1 U229 ( .A1(n28), .A2(n40), .B1(n42), .B2(n297), .C(n13), .ZN(n374)
         );
  AOI221D1 U230 ( .A1(n17), .A2(net7422), .B1(n7), .B2(net12847), .C(n228), 
        .ZN(n227) );
  OAI22D0 U231 ( .A1(n122), .A2(n160), .B1(n229), .B2(n128), .ZN(n228) );
  AOI221D1 U232 ( .A1(n64), .A2(n40), .B1(n56), .B2(n33), .C(n100), .ZN(n85)
         );
  OAI222D1 U233 ( .A1(n85), .A2(n86), .B1(net7431), .B2(n24), .C1(n87), .C2(
        net7422), .ZN(n79) );
  NR2XD0 U234 ( .A1(n88), .A2(n89), .ZN(n87) );
  OA221D1 U235 ( .A1(net7391), .A2(net8553), .B1(n270), .B2(n212), .C(n427), 
        .Z(n390) );
  BUFFD8 U236 ( .I(a[3]), .Z(net7431) );
  OR2XD1 U237 ( .A1(net7419), .A2(n137), .Z(n426) );
  ND2D1 U238 ( .A1(n34), .A2(n22), .ZN(n144) );
  BUFFD8 U239 ( .I(n66), .Z(net7419) );
  ND2D2 U240 ( .A1(n185), .A2(n19), .ZN(n137) );
  AOI221D1 U241 ( .A1(n22), .A2(n372), .B1(n63), .B2(n359), .C(n373), .ZN(n363) );
  AOI221D1 U242 ( .A1(n5), .A2(n223), .B1(n8), .B2(n62), .C(n224), .ZN(n206)
         );
  OAI222D1 U243 ( .A1(n225), .A2(n226), .B1(n106), .B2(n104), .C1(n227), .C2(
        n94), .ZN(n224) );
  ND2D1 U244 ( .A1(n57), .A2(net7422), .ZN(n161) );
  NR2D0 U245 ( .A1(n27), .A2(n16), .ZN(n229) );
  NR2D0 U246 ( .A1(n21), .A2(n10), .ZN(n201) );
  AOI211XD0 U247 ( .A1(n5), .A2(n376), .B(n377), .C(n378), .ZN(n362) );
  ND2D0 U248 ( .A1(n37), .A2(n25), .ZN(n258) );
  NR2XD0 U249 ( .A1(n31), .A2(n35), .ZN(n194) );
  CKND0 U250 ( .I(n90), .ZN(n26) );
  ND2D0 U251 ( .A1(n29), .A2(n40), .ZN(n335) );
  NR2D0 U252 ( .A1(n243), .A2(net12814), .ZN(n99) );
  NR2D0 U253 ( .A1(n57), .A2(n71), .ZN(n254) );
  CKND2D0 U254 ( .A1(n34), .A2(net7391), .ZN(n193) );
  NR2D0 U255 ( .A1(n69), .A2(n59), .ZN(n218) );
  ND2D1 U256 ( .A1(net7425), .A2(n371), .ZN(n368) );
  ND2D0 U257 ( .A1(net7427), .A2(n25), .ZN(n160) );
  ND2D0 U258 ( .A1(net7435), .A2(n59), .ZN(n138) );
  NR2D0 U259 ( .A1(n60), .A2(n64), .ZN(n396) );
  OAI22D0 U260 ( .A1(n111), .A2(n114), .B1(n213), .B2(n128), .ZN(n351) );
  OAI31D0 U261 ( .A1(n64), .A2(n9), .A3(n53), .B(n4), .ZN(n380) );
  CKND2D0 U262 ( .A1(n2), .A2(n40), .ZN(n82) );
  ND2D0 U263 ( .A1(n34), .A2(n5), .ZN(n191) );
  ND2D0 U264 ( .A1(n42), .A2(n2), .ZN(n105) );
  CKND2D0 U265 ( .A1(n43), .A2(n19), .ZN(n198) );
  ND2D0 U266 ( .A1(n67), .A2(n5), .ZN(n355) );
  NR2D0 U267 ( .A1(n149), .A2(n7), .ZN(n141) );
  CKND0 U268 ( .I(n231), .ZN(n11) );
  AOI22D0 U269 ( .A1(n12), .A2(n345), .B1(n174), .B2(n346), .ZN(n344) );
  CKND2D0 U270 ( .A1(net9112), .A2(n114), .ZN(n345) );
  CKND2D0 U271 ( .A1(n84), .A2(n182), .ZN(n346) );
  CKND2D1 U272 ( .A1(n379), .A2(n380), .ZN(n378) );
  AOI22D0 U273 ( .A1(net7422), .A2(n47), .B1(n51), .B2(n60), .ZN(n278) );
  OAI21D0 U274 ( .A1(net12708), .A2(n258), .B(n233), .ZN(n359) );
  OAI22D0 U275 ( .A1(net12814), .A2(n111), .B1(n266), .B2(n122), .ZN(n259) );
  NR2D0 U276 ( .A1(n39), .A2(n34), .ZN(n266) );
  NR2D0 U277 ( .A1(net7422), .A2(n107), .ZN(n125) );
  NR2XD0 U278 ( .A1(net8311), .A2(n9), .ZN(n177) );
  NR2D0 U279 ( .A1(n48), .A2(n41), .ZN(n213) );
  CKND2D0 U280 ( .A1(n68), .A2(net12847), .ZN(n147) );
  CKND2D0 U281 ( .A1(n36), .A2(n16), .ZN(n233) );
  CKND2D0 U282 ( .A1(n197), .A2(n16), .ZN(n279) );
  CKND2D0 U283 ( .A1(n185), .A2(n16), .ZN(n237) );
  CKND2D0 U284 ( .A1(n69), .A2(n51), .ZN(n145) );
  CKND2D0 U285 ( .A1(n33), .A2(n16), .ZN(n104) );
  CKND2D0 U287 ( .A1(n42), .A2(n16), .ZN(n262) );
  CKND2D1 U288 ( .A1(n272), .A2(n273), .ZN(n268) );
  OAI21D0 U289 ( .A1(net7435), .A2(n181), .B(n117), .ZN(n386) );
  NR2D0 U290 ( .A1(n55), .A2(n57), .ZN(n403) );
  AOI21D0 U291 ( .A1(n42), .A2(n6), .B(n172), .ZN(n367) );
  NR2XD0 U292 ( .A1(n221), .A2(n99), .ZN(n263) );
  AOI211D0 U293 ( .A1(n46), .A2(net7435), .B(n48), .C(n55), .ZN(n264) );
  AOI21D0 U294 ( .A1(n7), .A2(n47), .B(n172), .ZN(n169) );
  CKND2D0 U295 ( .A1(n181), .A2(n117), .ZN(n179) );
  OAI22D0 U296 ( .A1(net7422), .A2(n146), .B1(net7393), .B2(n135), .ZN(n343)
         );
  AOI32D0 U298 ( .A1(net7425), .A2(n45), .A3(n64), .B1(n59), .B2(n421), .ZN(
        n420) );
  NR2D0 U299 ( .A1(n7), .A2(n174), .ZN(n419) );
  CKND1 U300 ( .I(n204), .ZN(n18) );
  AOI21D0 U301 ( .A1(n8), .A2(net12847), .B(n174), .ZN(n173) );
  ND4D0 U302 ( .A1(n9), .A2(n28), .A3(net7429), .A4(net7425), .ZN(n140) );
  NR2D0 U303 ( .A1(n53), .A2(n60), .ZN(n422) );
  CKND2D0 U304 ( .A1(n138), .A2(n128), .ZN(n281) );
  OAI22D0 U305 ( .A1(n81), .A2(n82), .B1(n83), .B2(n84), .ZN(n80) );
  AOI21D0 U306 ( .A1(n182), .A2(n284), .B(net12814), .ZN(n418) );
  OAI32D0 U307 ( .A1(n98), .A2(n396), .A3(n162), .B1(n397), .B2(n128), .ZN(
        n393) );
  AOI31D0 U308 ( .A1(net7429), .A2(n30), .A3(n53), .B(n172), .ZN(n397) );
  AOI33D0 U309 ( .A1(n256), .A2(n30), .A3(n62), .B1(n10), .B2(n51), .B3(n67), 
        .ZN(n255) );
  CKND0 U310 ( .I(n258), .ZN(n23) );
  AOI22D0 U311 ( .A1(n57), .A2(net7435), .B1(net12847), .B2(n48), .ZN(n387) );
  OAI31D0 U312 ( .A1(n128), .A2(n41), .A3(n115), .B(n129), .ZN(n124) );
  AOI22D0 U313 ( .A1(n28), .A2(n118), .B1(n26), .B2(n59), .ZN(n110) );
  CKND2D0 U314 ( .A1(n103), .A2(n106), .ZN(n118) );
  AOI22D0 U315 ( .A1(n26), .A2(n59), .B1(n56), .B2(n27), .ZN(n401) );
  CKAN2D1 U316 ( .A1(n335), .A2(n135), .Z(n402) );
  ND2D0 U317 ( .A1(net7429), .A2(net7419), .ZN(n284) );
  AOI21D0 U318 ( .A1(n17), .A2(n48), .B(n113), .ZN(n112) );
  OAI21D0 U319 ( .A1(n158), .A2(n128), .B(n159), .ZN(n154) );
  OA33D0 U320 ( .A1(n160), .A2(net12708), .A3(net12814), .B1(n161), .B2(n162), 
        .B3(n98), .Z(n159) );
  AOI21D0 U321 ( .A1(n58), .A2(n19), .B(n298), .ZN(n357) );
  NR2D0 U322 ( .A1(net7429), .A2(n30), .ZN(n408) );
  OAI22D0 U323 ( .A1(net7393), .A2(n237), .B1(n238), .B2(net12814), .ZN(n236)
         );
  CKND2D0 U324 ( .A1(net12847), .A2(a[6]), .ZN(n385) );
  INVD1 U325 ( .I(n92), .ZN(n4) );
  INVD1 U326 ( .I(n82), .ZN(n1) );
  INVD1 U327 ( .I(n279), .ZN(n7) );
  INVD1 U328 ( .I(n237), .ZN(n14) );
  INVD1 U329 ( .I(n233), .ZN(n8) );
  INVD1 U330 ( .I(n103), .ZN(n60) );
  INVD1 U331 ( .I(n144), .ZN(n21) );
  INVD1 U332 ( .I(n271), .ZN(n13) );
  ND2D1 U333 ( .A1(n44), .A2(n28), .ZN(n165) );
  AOI21D1 U334 ( .A1(n50), .A2(net12847), .B(n61), .ZN(n285) );
  OAI222D0 U335 ( .A1(n139), .A2(n270), .B1(net9112), .B2(n104), .C1(n254), 
        .C2(n271), .ZN(n269) );
  IND4D1 U336 ( .A1(n73), .B1(n74), .B2(n75), .B3(n76), .ZN(d[0]) );
  OAI222D0 U337 ( .A1(n141), .A2(net9112), .B1(n143), .B2(n144), .C1(n145), 
        .C2(n146), .ZN(n73) );
  NR4D0 U338 ( .A1(n124), .A2(n125), .A3(n126), .A4(n127), .ZN(n75) );
  AOI221D0 U339 ( .A1(n132), .A2(n68), .B1(n50), .B2(n133), .C(n134), .ZN(n74)
         );
  NR2D1 U340 ( .A1(n248), .A2(n249), .ZN(n247) );
  OAI222D0 U341 ( .A1(n114), .A2(n181), .B1(n387), .B2(n101), .C1(net12847), 
        .C2(net12708), .ZN(n376) );
  NR4D0 U342 ( .A1(n154), .A2(n131), .A3(n155), .A4(n156), .ZN(n153) );
  NR4D0 U343 ( .A1(n393), .A2(n394), .A3(n155), .A4(n395), .ZN(n392) );
  NR3D0 U344 ( .A1(n360), .A2(net12708), .A3(n81), .ZN(n394) );
  OAI221D0 U345 ( .A1(net12847), .A2(n198), .B1(n145), .B2(n191), .C(n344), 
        .ZN(n327) );
  ND3D1 U346 ( .A1(n324), .A2(n325), .A3(n326), .ZN(d[5]) );
  AOI211D1 U347 ( .A1(n2), .A2(n351), .B(n352), .C(n353), .ZN(n324) );
  INR4D0 U348 ( .A1(n107), .B1(n347), .B2(n126), .B3(n156), .ZN(n325) );
  INVD1 U349 ( .I(n120), .ZN(n35) );
  INVD1 U350 ( .I(n212), .ZN(n28) );
  INVD1 U351 ( .I(n360), .ZN(n29) );
  NR3D0 U352 ( .A1(n196), .A2(n64), .A3(n68), .ZN(n219) );
  ND2D1 U353 ( .A1(n71), .A2(n39), .ZN(n270) );
  NR2D1 U354 ( .A1(n160), .A2(n157), .ZN(n149) );
  OAI31D1 U355 ( .A1(n196), .A2(net8311), .A3(n46), .B(n197), .ZN(n195) );
  ND2D1 U356 ( .A1(n34), .A2(n16), .ZN(n136) );
  OAI222D0 U357 ( .A1(net9112), .A2(n117), .B1(n177), .B2(n181), .C1(n111), 
        .C2(n315), .ZN(n337) );
  OAI222D0 U358 ( .A1(n136), .A2(n147), .B1(n169), .B2(net7422), .C1(n170), 
        .C2(n93), .ZN(n168) );
  NR4D0 U359 ( .A1(net7389), .A2(n25), .A3(n103), .A4(n111), .ZN(n171) );
  OAI221D0 U360 ( .A1(net12708), .A2(n114), .B1(n157), .B2(n81), .C(n234), 
        .ZN(n223) );
  OAI221D0 U361 ( .A1(n128), .A2(n182), .B1(n120), .B2(n163), .C(n183), .ZN(
        n175) );
  OAI222D0 U362 ( .A1(n90), .A2(n81), .B1(n91), .B2(n92), .C1(n93), .C2(n94), 
        .ZN(n89) );
  OAI222D0 U363 ( .A1(net7425), .A2(n95), .B1(n96), .B2(n97), .C1(n86), .C2(
        n98), .ZN(n88) );
  IAO21D1 U364 ( .A1(n98), .A2(n86), .B(n13), .ZN(n202) );
  NR4D0 U365 ( .A1(n416), .A2(n417), .A3(n339), .A4(n418), .ZN(n415) );
  INVD1 U366 ( .I(n99), .ZN(n24) );
  OAI222D0 U367 ( .A1(n356), .A2(net12814), .B1(n357), .B2(net12708), .C1(n358), .C2(n103), .ZN(n352) );
  NR2D1 U368 ( .A1(n4), .A2(n359), .ZN(n358) );
  OAI222D0 U369 ( .A1(n250), .A2(n92), .B1(n251), .B2(n144), .C1(n252), .C2(
        n111), .ZN(n249) );
  OA22D0 U370 ( .A1(n90), .A2(net12814), .B1(n139), .B2(n253), .Z(n252) );
  AOI221D0 U371 ( .A1(n59), .A2(n332), .B1(n19), .B2(n333), .C(n334), .ZN(n331) );
  NR4D0 U372 ( .A1(n209), .A2(n210), .A3(n211), .A4(n125), .ZN(n208) );
  ND2D1 U373 ( .A1(net7431), .A2(net7427), .ZN(n181) );
  OAI222D0 U374 ( .A1(net12847), .A2(n90), .B1(n122), .B2(n109), .C1(n115), 
        .C2(n119), .ZN(n383) );
  NR4D0 U375 ( .A1(n365), .A2(n366), .A3(n350), .A4(n349), .ZN(n364) );
  OAI222D0 U376 ( .A1(n108), .A2(n109), .B1(n110), .B2(n111), .C1(net7435), 
        .C2(n112), .ZN(n77) );
  NR3D0 U377 ( .A1(n128), .A2(net7429), .A3(n258), .ZN(n221) );
  OAI221D0 U378 ( .A1(n128), .A2(n139), .B1(net7389), .B2(n83), .C(n140), .ZN(
        n133) );
  AOI211XD0 U379 ( .A1(n21), .A2(net7435), .B(n230), .C(n11), .ZN(n225) );
  NR3D0 U380 ( .A1(net7422), .A2(net7429), .A3(n181), .ZN(n274) );
  NR2D1 U381 ( .A1(n107), .A2(net7435), .ZN(n155) );
  OAI221D0 U382 ( .A1(net7422), .A2(n135), .B1(n162), .B2(n148), .C(n173), 
        .ZN(n167) );
  NR3D0 U383 ( .A1(n147), .A2(net7429), .A3(n25), .ZN(n210) );
  AOI21D1 U384 ( .A1(n71), .A2(n220), .B(n221), .ZN(n217) );
  OAI222D0 U385 ( .A1(n396), .A2(n160), .B1(n403), .B2(n162), .C1(n139), .C2(
        n138), .ZN(n399) );
  INVD1 U386 ( .I(net7435), .ZN(n72) );
  OAI222D0 U387 ( .A1(n367), .A2(n122), .B1(n45), .B2(n368), .C1(n369), .C2(
        n148), .ZN(n365) );
  INR2D1 U388 ( .A1(n105), .B1(n370), .ZN(n369) );
  ND2D1 U389 ( .A1(net7431), .A2(net7419), .ZN(n94) );
  OAI222D0 U390 ( .A1(n114), .A2(n105), .B1(n177), .B2(n146), .C1(n178), .C2(
        n86), .ZN(n176) );
  AOI222D0 U391 ( .A1(n62), .A2(n43), .B1(n41), .B2(n60), .C1(n58), .C2(
        net7427), .ZN(n272) );
  AOI221D0 U392 ( .A1(n71), .A2(n50), .B1(n63), .B2(n35), .C(n274), .ZN(n273)
         );
  NR4D0 U393 ( .A1(n239), .A2(n240), .A3(n15), .A4(n241), .ZN(n238) );
  INVD2 U394 ( .I(a[2]), .ZN(n66) );
  AN2XD1 U395 ( .A1(net7435), .A2(n51), .Z(n196) );
  NR2XD0 U396 ( .A1(n32), .A2(n53), .ZN(n354) );
  OAI22D0 U397 ( .A1(n101), .A2(n182), .B1(n177), .B2(n157), .ZN(n417) );
  AOI21D0 U398 ( .A1(n181), .A2(n101), .B(net9112), .ZN(n186) );
  ND2D1 U399 ( .A1(n32), .A2(n25), .ZN(n243) );
  OAI22D0 U400 ( .A1(n120), .A2(n114), .B1(n101), .B2(n81), .ZN(n180) );
  ND2D0 U401 ( .A1(net7429), .A2(a[2]), .ZN(n163) );
  CKND2D0 U402 ( .A1(a[2]), .A2(n45), .ZN(n242) );
  AOI21D0 U403 ( .A1(n136), .A2(n198), .B(a[2]), .ZN(n240) );
  OAI222D0 U404 ( .A1(a[2]), .A2(n217), .B1(n218), .B2(n82), .C1(n219), .C2(
        n83), .ZN(n216) );
  CKND2D0 U405 ( .A1(a[2]), .A2(n128), .ZN(n130) );
  OA222D0 U406 ( .A1(n119), .A2(n120), .B1(n121), .B2(n122), .C1(n117), .C2(
        net12814), .Z(n108) );
  OAI33D0 U407 ( .A1(n212), .A2(net7435), .A3(net7419), .B1(n385), .B2(n139), 
        .B3(n106), .ZN(n384) );
  OAI22D0 U408 ( .A1(n226), .A2(net12814), .B1(n122), .B2(n94), .ZN(n371) );
  OAI21D0 U409 ( .A1(n226), .A2(n136), .B(n82), .ZN(n398) );
  OAI222D0 U410 ( .A1(n120), .A2(n315), .B1(n226), .B2(n148), .C1(n119), .C2(
        n181), .ZN(n416) );
  OAI222D0 U411 ( .A1(n109), .A2(n242), .B1(net7431), .B2(n243), .C1(n115), 
        .C2(n98), .ZN(n239) );
  INVD1 U412 ( .I(n106), .ZN(n55) );
  OAI222D0 U413 ( .A1(n103), .A2(n104), .B1(n105), .B2(n106), .C1(net12847), 
        .C2(n107), .ZN(n78) );
  NR4D0 U414 ( .A1(a[6]), .A2(n51), .A3(n139), .A4(n106), .ZN(n366) );
  OAI222D0 U415 ( .A1(n106), .A2(n98), .B1(n84), .B2(n222), .C1(n117), .C2(
        n161), .ZN(n214) );
  NR3D0 U416 ( .A1(n91), .A2(net7425), .A3(net7429), .ZN(n200) );
  OAI221D0 U417 ( .A1(n422), .A2(n257), .B1(n91), .B2(n148), .C(n423), .ZN(
        n412) );
  INVD1 U418 ( .I(n130), .ZN(n54) );
  AOI31D1 U419 ( .A1(n16), .A2(n130), .A3(n41), .B(n131), .ZN(n129) );
  AOI32D0 U420 ( .A1(net7427), .A2(net7422), .A3(n47), .B1(n36), .B2(n235), 
        .ZN(n234) );
  CKND2D0 U421 ( .A1(net7427), .A2(n30), .ZN(n360) );
  OAI32D0 U422 ( .A1(n312), .A2(n109), .A3(n120), .B1(n354), .B2(n355), .ZN(
        n353) );
  AOI21D0 U423 ( .A1(n257), .A2(n212), .B(n182), .ZN(n370) );
  OAI22D0 U424 ( .A1(net7425), .A2(n212), .B1(net12708), .B2(n139), .ZN(n421)
         );
  OAI22D0 U425 ( .A1(n30), .A2(n157), .B1(n45), .B2(n212), .ZN(n220) );
  INR2D1 U426 ( .A1(n348), .B1(net8772), .ZN(n156) );
  NR2D1 U427 ( .A1(n232), .A2(n145), .ZN(n126) );
  OAI222D0 U428 ( .A1(n232), .A2(net7419), .B1(n258), .B2(n265), .C1(net7431), 
        .C2(n146), .ZN(n260) );
  OAI22D0 U429 ( .A1(net7393), .A2(n146), .B1(net12847), .B2(n232), .ZN(n230)
         );
  INVD1 U430 ( .I(n270), .ZN(n38) );
  AN4D1 U431 ( .A1(n197), .A2(n47), .A3(net7435), .A4(n19), .Z(n350) );
  AOI31D0 U432 ( .A1(a[2]), .A2(n37), .A3(n9), .B(n38), .ZN(n375) );
  NR3D0 U433 ( .A1(n162), .A2(n37), .A3(n157), .ZN(n348) );
  NR4D0 U434 ( .A1(n157), .A2(n103), .A3(n109), .A4(n37), .ZN(n131) );
  NR3D0 U435 ( .A1(n37), .A2(net7389), .A3(net9112), .ZN(n339) );
  OAI211D0 U436 ( .A1(n37), .A2(n111), .B(n94), .C(net12708), .ZN(n184) );
  AOI22D1 U437 ( .A1(n53), .A2(n32), .B1(n50), .B2(n37), .ZN(n102) );
  INVD1 U438 ( .I(n111), .ZN(n43) );
  AOI31D0 U439 ( .A1(n135), .A2(n136), .A3(n137), .B(n138), .ZN(n134) );
  OAI21D0 U440 ( .A1(n212), .A2(n117), .B(n137), .ZN(n332) );
  OAI31D0 U441 ( .A1(n51), .A2(n61), .A3(n55), .B(n174), .ZN(n379) );
  AOI211D1 U442 ( .A1(n61), .A2(n41), .B(n38), .C(n171), .ZN(n170) );
  NR2D1 U443 ( .A1(n55), .A2(net7431), .ZN(n251) );
  OAI22D0 U444 ( .A1(net7431), .A2(n257), .B1(net7422), .B2(n258), .ZN(n256)
         );
  NR3D0 U445 ( .A1(n128), .A2(net7431), .A3(n101), .ZN(n338) );
  NR2D1 U446 ( .A1(n136), .A2(net7431), .ZN(n172) );
  AOI21D0 U447 ( .A1(net7431), .A2(n5), .B(n46), .ZN(n96) );
  NR2D1 U448 ( .A1(net7431), .A2(net7427), .ZN(n185) );
  NR2XD0 U449 ( .A1(net8311), .A2(n69), .ZN(n253) );
  CKND2D0 U450 ( .A1(net8311), .A2(n32), .ZN(n222) );
  AOI22D0 U451 ( .A1(n35), .A2(n59), .B1(n62), .B2(n33), .ZN(n423) );
  OAI22D0 U452 ( .A1(n415), .A2(n86), .B1(n119), .B2(n233), .ZN(n414) );
  NR4D0 U453 ( .A1(n181), .A2(n114), .A3(n86), .A4(n45), .ZN(n211) );
  AOI21D0 U454 ( .A1(n91), .A2(n121), .B(n86), .ZN(n241) );
endmodule


module aes_sbox_19 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n65, n67, n70, n73, n74, n77, n78, n192, n277, n304, n305, n306, n404,
         n405, n408, n409, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852;

  AN2XD1 U28 ( .A1(n713), .A2(n712), .Z(n717) );
  OA21D1 U35 ( .A1(n697), .A2(n696), .B(n695), .Z(n702) );
  OR3D1 U88 ( .A1(n665), .A2(n800), .A3(n445), .Z(n626) );
  OR4D1 U199 ( .A1(n650), .A2(n569), .A3(n516), .A4(n515), .Z(n518) );
  MAOI22D1 U209 ( .A1(n846), .A2(n802), .B1(n619), .B2(n767), .ZN(n509) );
  AN2XD1 U215 ( .A1(n517), .A2(n798), .Z(n516) );
  AN4XD1 U217 ( .A1(n664), .A2(n806), .A3(n436), .A4(n834), .Z(n515) );
  AN2XD1 U271 ( .A1(n530), .A2(n725), .Z(n463) );
  AO21D1 U297 ( .A1(n787), .A2(n824), .B(n728), .Z(n459) );
  BUFFD3 U1 ( .I(a[4]), .Z(n438) );
  OAI221D1 U2 ( .A1(n784), .A2(n725), .B1(n698), .B2(n712), .C(n687), .ZN(n693) );
  INVD2 U3 ( .I(n658), .ZN(n794) );
  CKND2D2 U4 ( .A1(a[2]), .A2(n445), .ZN(n658) );
  OAI222D1 U5 ( .A1(n775), .A2(n774), .B1(n437), .B2(n829), .C1(n773), .C2(
        n784), .ZN(n781) );
  CKND2D2 U6 ( .A1(n438), .A2(n802), .ZN(n703) );
  INVD3 U7 ( .I(n437), .ZN(n802) );
  ND2D3 U8 ( .A1(n784), .A2(n444), .ZN(n738) );
  AOI211XD0 U9 ( .A1(n830), .A2(n797), .B(n482), .C(n481), .ZN(n483) );
  OAI22D1 U10 ( .A1(n454), .A2(n774), .B1(n741), .B2(n628), .ZN(n455) );
  INVD2 U11 ( .I(n759), .ZN(n821) );
  OAI222D1 U12 ( .A1(n746), .A2(n755), .B1(n683), .B2(n714), .C1(n682), .C2(
        n774), .ZN(n684) );
  CKND2D2 U13 ( .A1(n816), .A2(n823), .ZN(n649) );
  INVD6 U14 ( .I(n439), .ZN(n816) );
  OAI222D1 U15 ( .A1(n799), .A2(n624), .B1(n550), .B2(n530), .C1(n529), .C2(
        n774), .ZN(n536) );
  AN2XD1 U16 ( .A1(n804), .A2(n594), .Z(n408) );
  OA222D0 U17 ( .A1(n461), .A2(n743), .B1(n679), .B2(n510), .C1(n460), .C2(
        n784), .Z(n74) );
  ND2D1 U18 ( .A1(n811), .A2(n837), .ZN(n599) );
  OA221D1 U19 ( .A1(n740), .A2(n732), .B1(n67), .B2(n658), .C(n435), .Z(n671)
         );
  AOI21D1 U20 ( .A1(n845), .A2(n442), .B(n686), .ZN(n687) );
  ND2D1 U21 ( .A1(n837), .A2(n821), .ZN(n629) );
  AOI211XD1 U22 ( .A1(n818), .A2(n581), .B(n579), .C(n580), .ZN(n582) );
  OAI222D1 U23 ( .A1(n739), .A2(n712), .B1(n763), .B2(n576), .C1(n744), .C2(
        n754), .ZN(n580) );
  ND2D4 U24 ( .A1(n819), .A2(n837), .ZN(n724) );
  INVD2 U25 ( .I(n604), .ZN(n819) );
  ND2D2 U26 ( .A1(n841), .A2(n784), .ZN(n630) );
  INVD1 U27 ( .I(n749), .ZN(n65) );
  INVD2 U29 ( .I(n65), .ZN(n67) );
  OAI222D1 U30 ( .A1(n658), .A2(n762), .B1(n436), .B2(n554), .C1(n744), .C2(
        n553), .ZN(n555) );
  OAI221D1 U31 ( .A1(n660), .A2(n670), .B1(n659), .B2(n658), .C(n835), .ZN(
        n662) );
  INVD3 U32 ( .I(n444), .ZN(n443) );
  BUFFD2 U33 ( .I(a[5]), .Z(n439) );
  ND2D1 U34 ( .A1(n785), .A2(n814), .ZN(n591) );
  INVD1 U36 ( .I(n629), .ZN(n843) );
  INVD2 U37 ( .I(a[6]), .ZN(n823) );
  ND2D1 U38 ( .A1(n438), .A2(n816), .ZN(n604) );
  ND2D1 U39 ( .A1(n443), .A2(a[2]), .ZN(n741) );
  ND2D1 U40 ( .A1(n808), .A2(n816), .ZN(n763) );
  NR2D1 U41 ( .A1(n427), .A2(n787), .ZN(n683) );
  BUFFD4 U42 ( .I(n788), .Z(n441) );
  INVD2 U43 ( .I(a[2]), .ZN(n788) );
  ND2D0 U44 ( .A1(n802), .A2(n808), .ZN(n749) );
  CKND2D1 U45 ( .A1(n437), .A2(n808), .ZN(n743) );
  INVD4 U46 ( .I(n438), .ZN(n808) );
  CKBD4 U47 ( .I(a[0]), .Z(n436) );
  ND2D1 U48 ( .A1(n800), .A2(n442), .ZN(n576) );
  INVD1 U49 ( .I(n766), .ZN(n800) );
  AOI211D1 U50 ( .A1(n792), .A2(n812), .B(n815), .C(n689), .ZN(n690) );
  INVD1 U51 ( .I(n779), .ZN(n791) );
  ND2D1 U52 ( .A1(n791), .A2(n784), .ZN(n550) );
  ND2D1 U53 ( .A1(n436), .A2(n444), .ZN(n737) );
  INVD2 U54 ( .I(n635), .ZN(n805) );
  ND2D1 U55 ( .A1(n784), .A2(n441), .ZN(n757) );
  OA221D1 U56 ( .A1(n445), .A2(n73), .B1(n591), .B2(n649), .C(n74), .Z(n475)
         );
  AOI221D1 U57 ( .A1(n789), .A2(n847), .B1(n798), .B2(n826), .C(n459), .ZN(
        n461) );
  OAI222D0 U58 ( .A1(a[2]), .A2(n644), .B1(n643), .B2(n778), .C1(n642), .C2(
        n777), .ZN(n645) );
  OAI221D0 U59 ( .A1(n732), .A2(n725), .B1(n698), .B2(n738), .C(n586), .ZN(
        n594) );
  INVD1 U60 ( .I(n751), .ZN(n848) );
  OAI222D0 U61 ( .A1(n718), .A2(n530), .B1(n484), .B2(n745), .C1(n483), .C2(
        n67), .ZN(n488) );
  OAI222D2 U62 ( .A1(n562), .A2(n703), .B1(n561), .B2(n737), .C1(n442), .C2(
        n560), .ZN(n563) );
  INVD2 U63 ( .I(n436), .ZN(n784) );
  INVD1 U64 ( .I(n444), .ZN(n442) );
  INVD1 U65 ( .I(a[1]), .ZN(n445) );
  CKND1 U66 ( .I(n732), .ZN(n424) );
  ND2D1 U67 ( .A1(a[1]), .A2(n784), .ZN(n732) );
  INVD1 U68 ( .I(n741), .ZN(n796) );
  AN3XD1 U69 ( .A1(n709), .A2(n708), .A3(n707), .Z(n70) );
  AOI21D2 U70 ( .A1(n850), .A2(n805), .B(n844), .ZN(n560) );
  OAI22D0 U71 ( .A1(n716), .A2(n746), .B1(n441), .B2(n723), .ZN(n657) );
  CKND2D0 U72 ( .A1(n441), .A2(n808), .ZN(n549) );
  ND2D3 U73 ( .A1(n445), .A2(n441), .ZN(n746) );
  AOI21D1 U74 ( .A1(n846), .A2(n806), .B(n688), .ZN(n691) );
  ND2D1 U75 ( .A1(n810), .A2(n834), .ZN(n663) );
  OAI32D0 U76 ( .A1(n762), .A2(n469), .A3(n698), .B1(n468), .B2(n732), .ZN(
        n472) );
  ND2D0 U77 ( .A1(n821), .A2(n828), .ZN(n618) );
  ND4D2 U78 ( .A1(n617), .A2(n616), .A3(n615), .A4(n614), .ZN(d[3]) );
  OAI222D0 U79 ( .A1(n746), .A2(n599), .B1(n598), .B2(n441), .C1(n669), .C2(
        n597), .ZN(n600) );
  AOI211XD0 U80 ( .A1(n807), .A2(n436), .B(n805), .C(n798), .ZN(n597) );
  NR2D0 U81 ( .A1(n505), .A2(n658), .ZN(n564) );
  AOI31D1 U82 ( .A1(n791), .A2(n848), .A3(n675), .B(n711), .ZN(n433) );
  NR3D1 U83 ( .A1(n425), .A2(n426), .A3(n673), .ZN(n710) );
  AOI221D2 U84 ( .A1(n801), .A2(n565), .B1(n564), .B2(n811), .C(n563), .ZN(
        n573) );
  AOI221D1 U85 ( .A1(n850), .A2(n444), .B1(n832), .B2(n712), .C(n522), .ZN(
        n525) );
  OAI222D0 U86 ( .A1(n525), .A2(n769), .B1(n718), .B2(n618), .C1(n524), .C2(
        n712), .ZN(n537) );
  CKND2D2 U87 ( .A1(n437), .A2(a[2]), .ZN(n635) );
  ND2D2 U89 ( .A1(n440), .A2(n823), .ZN(n751) );
  OA221D0 U90 ( .A1(n458), .A2(n769), .B1(n714), .B2(n766), .C(n559), .Z(n73)
         );
  NR3D1 U91 ( .A1(n408), .A2(n409), .A3(n592), .ZN(n616) );
  AOI211XD0 U92 ( .A1(n852), .A2(n797), .B(n477), .C(n657), .ZN(n504) );
  CKND2D2 U93 ( .A1(n823), .A2(n828), .ZN(n745) );
  AOI211XD0 U94 ( .A1(n832), .A2(n436), .B(n631), .C(n842), .ZN(n636) );
  ND2D1 U95 ( .A1(n437), .A2(n441), .ZN(n766) );
  ND4D3 U96 ( .A1(n476), .A2(n475), .A3(n474), .A4(n473), .ZN(d[7]) );
  INVD2 U97 ( .I(n746), .ZN(n789) );
  INVD1 U98 ( .I(n553), .ZN(n790) );
  OAI22D1 U99 ( .A1(n738), .A2(n700), .B1(n632), .B2(n732), .ZN(n633) );
  OAI222D1 U100 ( .A1(n751), .A2(n619), .B1(n437), .B2(n618), .C1(n745), .C2(
        n762), .ZN(n622) );
  INVD1 U101 ( .I(n791), .ZN(n77) );
  AOI22D1 U102 ( .A1(n791), .A2(n825), .B1(n800), .B2(n808), .ZN(n765) );
  CKND3 U103 ( .I(a[1]), .ZN(n444) );
  NR2XD1 U104 ( .A1(n772), .A2(n771), .ZN(n773) );
  NR2XD0 U105 ( .A1(n808), .A2(n816), .ZN(n664) );
  OAI22D1 U106 ( .A1(n759), .A2(n769), .B1(n442), .B2(n758), .ZN(n760) );
  AOI32D1 U107 ( .A1(n439), .A2(n784), .A3(n806), .B1(n817), .B2(n626), .ZN(
        n627) );
  OAI33D0 U108 ( .A1(n649), .A2(n436), .A3(n441), .B1(n480), .B2(n721), .B3(
        n754), .ZN(n481) );
  CKND2D1 U109 ( .A1(n440), .A2(n816), .ZN(n721) );
  OAI22D0 U110 ( .A1(n440), .A2(n649), .B1(n744), .B2(n721), .ZN(n448) );
  INVD1 U111 ( .I(n721), .ZN(n847) );
  AOI221D1 U112 ( .A1(n834), .A2(n602), .B1(n601), .B2(n784), .C(n600), .ZN(
        n615) );
  IAO21D2 U113 ( .A1(n678), .A2(n445), .B(n792), .ZN(n577) );
  ND2D1 U114 ( .A1(n437), .A2(n816), .ZN(n740) );
  OAI33D0 U115 ( .A1(n67), .A2(n441), .A3(n721), .B1(n649), .B2(n442), .B3(
        n648), .ZN(n652) );
  OA221D1 U116 ( .A1(n553), .A2(n624), .B1(n712), .B2(n778), .C(n78), .Z(n617)
         );
  OA222D1 U117 ( .A1(n635), .A2(n628), .B1(n584), .B2(n583), .C1(n751), .C2(
        n582), .Z(n78) );
  CKND1 U118 ( .I(n712), .ZN(n785) );
  OA221D1 U119 ( .A1(n432), .A2(n741), .B1(n724), .B2(n776), .C(n433), .Z(n460) );
  OAI222D1 U120 ( .A1(n440), .A2(n765), .B1(n764), .B2(n763), .C1(n774), .C2(
        n762), .ZN(n772) );
  AOI22D1 U121 ( .A1(n800), .A2(n821), .B1(n803), .B2(n816), .ZN(n758) );
  AOI221D1 U122 ( .A1(n831), .A2(n647), .B1(n834), .B2(n646), .C(n645), .ZN(
        n654) );
  OAI22D1 U123 ( .A1(n445), .A2(n624), .B1(n623), .B2(n737), .ZN(n625) );
  OAI222D1 U124 ( .A1(n636), .A2(n635), .B1(n754), .B2(n756), .C1(n766), .C2(
        n634), .ZN(n637) );
  OAI221D1 U125 ( .A1(n603), .A2(n578), .B1(n437), .B2(n768), .C(n695), .ZN(
        n523) );
  AOI221D1 U126 ( .A1(n811), .A2(n848), .B1(n800), .B2(n821), .C(n523), .ZN(
        n524) );
  NR3D1 U127 ( .A1(n637), .A2(n305), .A3(n306), .ZN(n655) );
  AOI22D1 U128 ( .A1(n819), .A2(n805), .B1(n794), .B2(n816), .ZN(n554) );
  AOI221D1 U129 ( .A1(n787), .A2(n676), .B1(n675), .B2(n794), .C(n674), .ZN(
        n677) );
  CKND2D1 U130 ( .A1(n436), .A2(n441), .ZN(n718) );
  OAI222D1 U131 ( .A1(n718), .A2(n743), .B1(n683), .B2(n679), .C1(n67), .C2(
        n550), .ZN(n528) );
  ND2D1 U132 ( .A1(n789), .A2(n436), .ZN(n553) );
  OAI222D1 U133 ( .A1(n777), .A2(n576), .B1(n769), .B2(n630), .C1(n491), .C2(
        n757), .ZN(n492) );
  ND2D1 U134 ( .A1(n438), .A2(n437), .ZN(n744) );
  INVD0 U135 ( .I(n744), .ZN(n812) );
  AOI221D1 U136 ( .A1(n794), .A2(n533), .B1(n834), .B2(n532), .C(n531), .ZN(
        n534) );
  OAI21D1 U137 ( .A1(n744), .A2(n603), .B(n628), .ZN(n506) );
  OA221D1 U138 ( .A1(n784), .A2(n192), .B1(n774), .B2(n277), .C(n304), .Z(n574) );
  OA211D0 U139 ( .A1(n696), .A2(n670), .B(n545), .C(n544), .Z(n192) );
  OA211D0 U140 ( .A1(n549), .A2(n712), .B(n548), .C(n547), .Z(n277) );
  OA222D1 U141 ( .A1(n558), .A2(n751), .B1(n678), .B2(n557), .C1(n745), .C2(
        n556), .Z(n304) );
  ND2D1 U142 ( .A1(a[6]), .A2(n828), .ZN(n774) );
  INVD4 U143 ( .I(n440), .ZN(n828) );
  OAI222D1 U144 ( .A1(n436), .A2(n672), .B1(n671), .B2(n745), .C1(n670), .C2(
        n669), .ZN(n673) );
  NR4D1 U145 ( .A1(n528), .A2(n527), .A3(n526), .A4(n587), .ZN(n529) );
  AOI221D1 U146 ( .A1(n424), .A2(n681), .B1(n822), .B2(n427), .C(n680), .ZN(
        n682) );
  AOI221D1 U147 ( .A1(n825), .A2(n813), .B1(n811), .B2(n565), .C(n840), .ZN(
        n491) );
  OA222D0 U148 ( .A1(n719), .A2(n718), .B1(n717), .B2(n716), .C1(n715), .C2(
        n714), .Z(n430) );
  OAI33D0 U149 ( .A1(n746), .A2(n745), .A3(n744), .B1(n767), .B2(n441), .B3(
        n743), .ZN(n747) );
  ND2D2 U150 ( .A1(n443), .A2(n436), .ZN(n712) );
  ND2D2 U151 ( .A1(n440), .A2(a[6]), .ZN(n698) );
  CKBD4 U152 ( .I(a[7]), .Z(n440) );
  AOI221D1 U153 ( .A1(n686), .A2(n738), .B1(n442), .B2(n843), .C(n552), .ZN(
        n557) );
  OAI31D0 U154 ( .A1(n698), .A2(n439), .A3(n442), .B(n630), .ZN(n552) );
  ND2D1 U155 ( .A1(n831), .A2(n664), .ZN(n725) );
  NR4D1 U156 ( .A1(n622), .A2(n621), .A3(n838), .A4(n620), .ZN(n623) );
  AOI221D1 U157 ( .A1(n824), .A2(n785), .B1(n585), .B2(n444), .C(n434), .ZN(
        n586) );
  AOI221D1 U158 ( .A1(n834), .A2(n457), .B1(n456), .B2(n784), .C(n455), .ZN(
        n476) );
  AOI221D1 U159 ( .A1(n467), .A2(n444), .B1(n810), .B2(n466), .C(n465), .ZN(
        n474) );
  OAI22D0 U160 ( .A1(n464), .A2(n703), .B1(n463), .B2(n754), .ZN(n465) );
  ND4D2 U161 ( .A1(n656), .A2(n655), .A3(n654), .A4(n653), .ZN(d[2]) );
  AOI221D4 U162 ( .A1(n849), .A2(n784), .B1(n841), .B2(n796), .C(n625), .ZN(
        n656) );
  AOI211XD0 U163 ( .A1(n848), .A2(n489), .B(n488), .C(n487), .ZN(n503) );
  ND4D2 U164 ( .A1(n574), .A2(n575), .A3(n573), .A4(n572), .ZN(d[4]) );
  CKAN2D1 U165 ( .A1(n848), .A2(n638), .Z(n305) );
  CKAN2D1 U166 ( .A1(n845), .A2(n791), .Z(n306) );
  CKAN2D1 U167 ( .A1(n789), .A2(n813), .Z(n404) );
  CKAN2D1 U168 ( .A1(n797), .A2(n820), .Z(n405) );
  NR3D0 U169 ( .A1(n404), .A2(n405), .A3(n760), .ZN(n775) );
  INVD1 U170 ( .I(n703), .ZN(n813) );
  INVD0 U171 ( .I(n679), .ZN(n820) );
  CKAN2D1 U172 ( .A1(n831), .A2(n593), .Z(n409) );
  INVD2 U173 ( .I(n774), .ZN(n831) );
  NR4D1 U174 ( .A1(n428), .A2(n429), .A3(n781), .A4(n780), .ZN(n782) );
  AOI221D1 U175 ( .A1(n831), .A2(n493), .B1(n790), .B2(n506), .C(n492), .ZN(
        n502) );
  NR4D1 U176 ( .A1(n537), .A2(n538), .A3(n536), .A4(n535), .ZN(n539) );
  AOI222D1 U177 ( .A1(n796), .A2(n819), .B1(n794), .B2(n479), .C1(n790), .C2(
        n822), .ZN(n484) );
  NR2D1 U178 ( .A1(n784), .A2(n437), .ZN(n665) );
  OA21D0 U179 ( .A1(n678), .A2(n784), .B(n607), .Z(n611) );
  CKND1 U180 ( .I(n754), .ZN(n798) );
  ND2D0 U181 ( .A1(n436), .A2(n794), .ZN(n722) );
  NR2D0 U182 ( .A1(n745), .A2(n763), .ZN(n686) );
  OAI31D0 U183 ( .A1(n741), .A2(n770), .A3(n743), .B(n606), .ZN(n613) );
  ND2D0 U184 ( .A1(n439), .A2(n828), .ZN(n700) );
  CKAN2D1 U185 ( .A1(n839), .A2(n798), .Z(n425) );
  CKAN2D1 U186 ( .A1(n686), .A2(n791), .Z(n426) );
  CKND2D2 U187 ( .A1(n710), .A2(n70), .ZN(d[1]) );
  CKAN2D1 U188 ( .A1(n436), .A2(n441), .Z(n427) );
  CKND2D0 U189 ( .A1(n804), .A2(n442), .ZN(n713) );
  NR2D0 U190 ( .A1(n805), .A2(n812), .ZN(n648) );
  INVD1 U191 ( .I(n724), .ZN(n841) );
  NR2D0 U192 ( .A1(n826), .A2(n837), .ZN(n632) );
  CKND2D0 U193 ( .A1(n664), .A2(n837), .ZN(n583) );
  CKND2D0 U194 ( .A1(n817), .A2(n837), .ZN(n628) );
  CKND2D0 U195 ( .A1(n675), .A2(n837), .ZN(n624) );
  ND2D0 U196 ( .A1(a[2]), .A2(n802), .ZN(n769) );
  ND2D1 U197 ( .A1(n442), .A2(n437), .ZN(n776) );
  ND2D0 U198 ( .A1(n440), .A2(n494), .ZN(n497) );
  NR2XD0 U200 ( .A1(n849), .A2(n506), .ZN(n507) );
  OAI211D0 U201 ( .A1(n439), .A2(n776), .B(n619), .C(n743), .ZN(n532) );
  AOI221D1 U202 ( .A1(n811), .A2(n786), .B1(n820), .B2(n796), .C(n555), .ZN(
        n556) );
  ND2D0 U203 ( .A1(a[2]), .A2(n808), .ZN(n619) );
  CKND0 U204 ( .I(n730), .ZN(n799) );
  CKND2D1 U205 ( .A1(n767), .A2(n721), .ZN(n565) );
  CKND2D0 U206 ( .A1(n438), .A2(a[2]), .ZN(n697) );
  BUFFD4 U207 ( .I(a[3]), .Z(n437) );
  NR2D0 U208 ( .A1(n793), .A2(n789), .ZN(n469) );
  CKND0 U210 ( .I(n768), .ZN(n849) );
  CKND0 U211 ( .I(n576), .ZN(n801) );
  ND3D0 U212 ( .A1(n805), .A2(n664), .A3(n834), .ZN(n753) );
  AOI22D0 U213 ( .A1(n850), .A2(n791), .B1(n806), .B2(n836), .ZN(n544) );
  NR2D0 U214 ( .A1(n796), .A2(n785), .ZN(n607) );
  ND2D0 U216 ( .A1(n819), .A2(n848), .ZN(n669) );
  ND2D0 U218 ( .A1(n811), .A2(n851), .ZN(n755) );
  ND2D0 U219 ( .A1(n800), .A2(n843), .ZN(n559) );
  NR2D0 U220 ( .A1(n711), .A2(n846), .ZN(n719) );
  ND2D0 U221 ( .A1(n824), .A2(n813), .ZN(n530) );
  ND2D0 U222 ( .A1(n424), .A2(n848), .ZN(n510) );
  NR2D0 U223 ( .A1(n850), .A2(n836), .ZN(n458) );
  AOI21D0 U224 ( .A1(n809), .A2(n851), .B(n838), .ZN(n561) );
  AOI22D0 U225 ( .A1(n797), .A2(n847), .B1(n789), .B2(n826), .ZN(n562) );
  ND2D0 U226 ( .A1(n427), .A2(n821), .ZN(n639) );
  ND2D0 U227 ( .A1(n679), .A2(n743), .ZN(n681) );
  ND2D0 U228 ( .A1(n441), .A2(n802), .ZN(n678) );
  CKND2D0 U229 ( .A1(n776), .A2(n678), .ZN(n519) );
  CKND2D0 U230 ( .A1(n718), .A2(n746), .ZN(n520) );
  NR2D0 U231 ( .A1(n800), .A2(n793), .ZN(n447) );
  AOI22D0 U232 ( .A1(n818), .A2(n794), .B1(n791), .B2(n820), .ZN(n446) );
  OAI32D0 U233 ( .A1(n553), .A2(n751), .A3(n740), .B1(n511), .B2(n510), .ZN(
        n512) );
  NR2D0 U234 ( .A1(n821), .A2(n800), .ZN(n511) );
  CKND2D0 U235 ( .A1(n722), .A2(n732), .ZN(n581) );
  OAI31D0 U236 ( .A1(n732), .A2(n812), .A3(n745), .B(n731), .ZN(n736) );
  ND2D0 U237 ( .A1(n816), .A2(n828), .ZN(n603) );
  AOI22D0 U238 ( .A1(n784), .A2(n806), .B1(n802), .B2(n793), .ZN(n584) );
  AOI32D0 U239 ( .A1(n789), .A2(n784), .A3(n822), .B1(n424), .B2(n546), .ZN(
        n548) );
  CKND2D0 U240 ( .A1(n744), .A2(n739), .ZN(n546) );
  NR2D0 U241 ( .A1(n814), .A2(n819), .ZN(n595) );
  NR2D0 U242 ( .A1(n784), .A2(n753), .ZN(n735) );
  AOI22D0 U243 ( .A1(n827), .A2(n794), .B1(n797), .B2(n826), .ZN(n464) );
  CKND2D0 U244 ( .A1(n796), .A2(n784), .ZN(n699) );
  OAI211D0 U245 ( .A1(n816), .A2(n67), .B(n766), .C(n744), .ZN(n676) );
  ND2D0 U246 ( .A1(n819), .A2(n831), .ZN(n716) );
  AOI21D0 U247 ( .A1(n604), .A2(n649), .B(n678), .ZN(n495) );
  AOI31D0 U248 ( .A1(n725), .A2(n724), .A3(n723), .B(n722), .ZN(n726) );
  AOI22D0 U249 ( .A1(n825), .A2(n742), .B1(n827), .B2(n794), .ZN(n750) );
  CKND2D0 U250 ( .A1(n757), .A2(n754), .ZN(n742) );
  AOI21D0 U251 ( .A1(n679), .A2(n759), .B(n718), .ZN(n674) );
  OAI21D0 U252 ( .A1(n649), .A2(n743), .B(n723), .ZN(n533) );
  CKND2D0 U253 ( .A1(n786), .A2(n802), .ZN(n715) );
  OAI21D0 U254 ( .A1(n635), .A2(n724), .B(n778), .ZN(n467) );
  CKND0 U255 ( .I(n696), .ZN(n851) );
  CKND2D0 U256 ( .A1(n819), .A2(n444), .ZN(n668) );
  OAI31D0 U257 ( .A1(n789), .A2(n787), .A3(n800), .B(n849), .ZN(n485) );
  OAI31D0 U258 ( .A1(n802), .A2(n792), .A3(n798), .B(n686), .ZN(n486) );
  OAI21D0 U259 ( .A1(n436), .A2(n679), .B(n743), .ZN(n479) );
  AOI31D0 U260 ( .A1(a[2]), .A2(n816), .A3(n787), .B(n815), .ZN(n490) );
  AOI22D0 U261 ( .A1(n796), .A2(n436), .B1(n442), .B2(n805), .ZN(n478) );
  AOI21D0 U262 ( .A1(n795), .A2(n834), .B(n564), .ZN(n508) );
  AOI21D0 U263 ( .A1(n437), .A2(n848), .B(n807), .ZN(n764) );
  NR2D0 U264 ( .A1(n798), .A2(n437), .ZN(n610) );
  NR2D0 U265 ( .A1(n798), .A2(n796), .ZN(n462) );
  AOI21D0 U266 ( .A1(n678), .A2(n578), .B(n737), .ZN(n451) );
  AOI21D0 U267 ( .A1(n811), .A2(n847), .B(n688), .ZN(n498) );
  CKND2D0 U268 ( .A1(n712), .A2(n802), .ZN(n567) );
  NR2D0 U269 ( .A1(n792), .A2(n795), .ZN(n568) );
  AOI22D0 U270 ( .A1(n814), .A2(n786), .B1(n812), .B2(a[2]), .ZN(n566) );
  OAI33D0 U272 ( .A1(n635), .A2(n440), .A3(n763), .B1(n696), .B2(n441), .B3(
        n744), .ZN(n531) );
  CKND2D0 U273 ( .A1(n805), .A2(n808), .ZN(n596) );
  NR2XD0 U274 ( .A1(n640), .A2(n761), .ZN(n598) );
  NR2XD0 U275 ( .A1(n786), .A2(n794), .ZN(n643) );
  ND4D0 U276 ( .A1(n787), .A2(n825), .A3(n438), .A4(n440), .ZN(n720) );
  AOI32D0 U277 ( .A1(n440), .A2(n808), .A3(n789), .B1(n794), .B2(n448), .ZN(
        n449) );
  NR2D0 U278 ( .A1(n846), .A2(n686), .ZN(n450) );
  INVD2 U279 ( .I(n698), .ZN(n837) );
  AOI31D0 U280 ( .A1(n438), .A2(n823), .A3(n800), .B(n688), .ZN(n468) );
  OAI21D0 U281 ( .A1(n702), .A2(n732), .B(n701), .ZN(n706) );
  AOI211D0 U282 ( .A1(n770), .A2(n649), .B(n578), .C(n737), .ZN(n470) );
  AOI33D0 U283 ( .A1(n605), .A2(n823), .A3(n791), .B1(n843), .B2(n802), .B3(
        n424), .ZN(n606) );
  OAI22D0 U284 ( .A1(n437), .A2(n604), .B1(n784), .B2(n603), .ZN(n605) );
  NR2D0 U285 ( .A1(n724), .A2(n437), .ZN(n688) );
  ND2D0 U286 ( .A1(n439), .A2(n802), .ZN(n762) );
  OAI22D0 U287 ( .A1(n823), .A2(n703), .B1(n808), .B2(n649), .ZN(n641) );
  AOI21D0 U288 ( .A1(n724), .A2(n663), .B(a[2]), .ZN(n621) );
  CKND2D0 U289 ( .A1(n438), .A2(n441), .ZN(n578) );
  CKND2D0 U290 ( .A1(a[2]), .A2(n732), .ZN(n730) );
  CKND2D0 U291 ( .A1(n437), .A2(n445), .ZN(n670) );
  CKND2D1 U292 ( .A1(n589), .A2(n588), .ZN(n593) );
  AOI21D0 U293 ( .A1(n836), .A2(n805), .B(n747), .ZN(n748) );
  INVD1 U294 ( .I(n777), .ZN(n836) );
  INVD1 U295 ( .I(n669), .ZN(n850) );
  INVD1 U296 ( .I(n778), .ZN(n852) );
  INVD1 U298 ( .I(n591), .ZN(n815) );
  INVD1 U299 ( .I(n559), .ZN(n844) );
  AOI222D0 U300 ( .A1(n796), .A2(n813), .B1(n811), .B2(n427), .C1(n820), .C2(
        n794), .ZN(n547) );
  ND2D1 U301 ( .A1(n664), .A2(n848), .ZN(n768) );
  ND2D1 U302 ( .A1(n834), .A2(n821), .ZN(n777) );
  NR2D1 U303 ( .A1(n629), .A2(n715), .ZN(n734) );
  INVD1 U304 ( .I(n699), .ZN(n797) );
  INVD1 U305 ( .I(n583), .ZN(n846) );
  ND2D1 U306 ( .A1(n851), .A2(n813), .ZN(n778) );
  INVD1 U307 ( .I(n757), .ZN(n793) );
  INVD1 U308 ( .I(n678), .ZN(n803) );
  INVD1 U309 ( .I(n763), .ZN(n817) );
  INVD1 U310 ( .I(n624), .ZN(n839) );
  INVD1 U311 ( .I(n716), .ZN(n832) );
  AO221D0 U312 ( .A1(n789), .A2(n822), .B1(n424), .B2(n804), .C(n694), .Z(n646) );
  INVD1 U313 ( .I(n628), .ZN(n845) );
  ND2D1 U314 ( .A1(n809), .A2(n825), .ZN(n695) );
  INVD1 U315 ( .I(n550), .ZN(n792) );
  INVD1 U316 ( .I(n603), .ZN(n830) );
  INVD1 U317 ( .I(n549), .ZN(n809) );
  INVD1 U318 ( .I(n599), .ZN(n838) );
  INVD1 U319 ( .I(n590), .ZN(n840) );
  ND2D1 U320 ( .A1(n776), .A2(n550), .ZN(n551) );
  OAI221D0 U321 ( .A1(n744), .A2(n746), .B1(n703), .B2(n77), .C(n627), .ZN(
        n638) );
  AOI221D0 U322 ( .A1(n836), .A2(n784), .B1(n846), .B2(n442), .C(n633), .ZN(
        n634) );
  OAI222D0 U323 ( .A1(n754), .A2(n762), .B1(n776), .B2(n639), .C1(n743), .C2(
        n699), .ZN(n647) );
  NR4D0 U324 ( .A1(n703), .A2(n757), .A3(n751), .A4(n816), .ZN(n729) );
  OAI222D0 U325 ( .A1(n721), .A2(n591), .B1(n718), .B2(n756), .C1(n607), .C2(
        n590), .ZN(n592) );
  OAI222D0 U326 ( .A1(n718), .A2(n590), .B1(n725), .B2(n670), .C1(n629), .C2(
        n754), .ZN(n542) );
  NR2D1 U327 ( .A1(n696), .A2(n738), .ZN(n728) );
  NR2D1 U328 ( .A1(n832), .A2(n843), .ZN(n660) );
  INVD1 U329 ( .I(n657), .ZN(n835) );
  NR4D0 U330 ( .A1(n571), .A2(n570), .A3(n569), .A4(n733), .ZN(n572) );
  AOI221D0 U331 ( .A1(n800), .A2(n833), .B1(n841), .B2(n806), .C(n542), .ZN(
        n575) );
  INVD1 U332 ( .I(n743), .ZN(n811) );
  NR4D0 U333 ( .A1(n472), .A2(n471), .A3(n705), .A4(n470), .ZN(n473) );
  NR2D1 U334 ( .A1(n613), .A2(n612), .ZN(n614) );
  ND2D1 U335 ( .A1(n486), .A2(n485), .ZN(n487) );
  OAI221D0 U336 ( .A1(n442), .A2(n663), .B1(n715), .B2(n669), .C(n521), .ZN(
        n538) );
  NR4D0 U337 ( .A1(n652), .A2(n651), .A3(n650), .A4(n735), .ZN(n653) );
  ND4D1 U338 ( .A1(n430), .A2(n431), .A3(n783), .A4(n782), .ZN(d[0]) );
  NR4D0 U339 ( .A1(n736), .A2(n735), .A3(n734), .A4(n733), .ZN(n783) );
  AOI221D0 U340 ( .A1(n434), .A2(n804), .B1(n803), .B2(n727), .C(n726), .ZN(
        n431) );
  NR3D0 U341 ( .A1(n816), .A2(n443), .A3(n718), .ZN(n526) );
  ND2D1 U342 ( .A1(n675), .A2(n834), .ZN(n723) );
  OAI221D0 U343 ( .A1(n447), .A2(n604), .B1(n769), .B2(n712), .C(n446), .ZN(
        n457) );
  NR3D0 U344 ( .A1(n712), .A2(n808), .A3(n723), .ZN(n569) );
  OAI22D1 U345 ( .A1(n759), .A2(n678), .B1(n683), .B2(n703), .ZN(n452) );
  AOI31D1 U346 ( .A1(n837), .A2(n730), .A3(n812), .B(n729), .ZN(n731) );
  INVD1 U347 ( .I(n649), .ZN(n825) );
  INVD1 U348 ( .I(n737), .ZN(n787) );
  INVD1 U349 ( .I(n740), .ZN(n818) );
  ND3D1 U350 ( .A1(n541), .A2(n540), .A3(n539), .ZN(d[5]) );
  AOI211D1 U351 ( .A1(n851), .A2(n514), .B(n513), .C(n512), .ZN(n541) );
  INR4D0 U352 ( .A1(n753), .B1(n518), .B2(n734), .B3(n704), .ZN(n540) );
  ND2D1 U353 ( .A1(n831), .A2(n817), .ZN(n714) );
  INVD1 U354 ( .I(n762), .ZN(n822) );
  ND2D1 U355 ( .A1(n443), .A2(n441), .ZN(n779) );
  NR2D1 U356 ( .A1(n618), .A2(n737), .ZN(n761) );
  ND2D1 U357 ( .A1(n818), .A2(n837), .ZN(n590) );
  INVD1 U358 ( .I(n769), .ZN(n804) );
  NR2D1 U359 ( .A1(n619), .A2(n712), .ZN(n694) );
  ND2D1 U360 ( .A1(n820), .A2(n837), .ZN(n756) );
  INVD1 U361 ( .I(n722), .ZN(n795) );
  INVD1 U362 ( .I(n670), .ZN(n807) );
  INVD1 U363 ( .I(n745), .ZN(n834) );
  INVD1 U364 ( .I(n697), .ZN(n814) );
  OA221D0 U365 ( .A1(n678), .A2(n668), .B1(n667), .B2(n77), .C(n666), .Z(n435)
         );
  OAI31D1 U366 ( .A1(n665), .A2(n427), .A3(n807), .B(n664), .ZN(n666) );
  INVD1 U367 ( .I(n505), .ZN(n824) );
  OAI222D0 U368 ( .A1(n469), .A2(n700), .B1(n462), .B2(n698), .C1(n721), .C2(
        n722), .ZN(n466) );
  INVD1 U369 ( .I(n761), .ZN(n829) );
  OAI221D0 U370 ( .A1(n608), .A2(n759), .B1(n744), .B2(n754), .C(n490), .ZN(
        n493) );
  INR4D0 U371 ( .A1(n663), .B1(n844), .B2(n661), .B3(n662), .ZN(n672) );
  NR3D0 U372 ( .A1(n769), .A2(n440), .A3(n438), .ZN(n661) );
  OAI222D0 U373 ( .A1(n746), .A2(n679), .B1(n478), .B2(n759), .C1(n442), .C2(
        n744), .ZN(n489) );
  OAI222D0 U374 ( .A1(n498), .A2(n738), .B1(n808), .B2(n497), .C1(n496), .C2(
        n712), .ZN(n500) );
  INR2D1 U375 ( .A1(n755), .B1(n495), .ZN(n496) );
  OAI222D0 U376 ( .A1(n699), .A2(n725), .B1(n436), .B2(n534), .C1(n77), .C2(
        n768), .ZN(n535) );
  OAI221D0 U377 ( .A1(n732), .A2(n678), .B1(n740), .B2(n697), .C(n677), .ZN(
        n685) );
  OAI222D0 U378 ( .A1(n724), .A2(n713), .B1(n691), .B2(n784), .C1(n690), .C2(
        n767), .ZN(n692) );
  OAI222D0 U379 ( .A1(n509), .A2(n737), .B1(n508), .B2(n744), .C1(n507), .C2(
        n757), .ZN(n513) );
  OAI222D0 U380 ( .A1(n611), .A2(n768), .B1(n610), .B2(n716), .C1(n609), .C2(
        n67), .ZN(n612) );
  OA22D0 U381 ( .A1(n770), .A2(n737), .B1(n721), .B2(n608), .Z(n609) );
  NR3D0 U382 ( .A1(n784), .A2(n438), .A3(n679), .ZN(n587) );
  NR3D0 U383 ( .A1(n665), .A2(n789), .A3(n804), .ZN(n642) );
  AOI21D1 U384 ( .A1(n785), .A2(n641), .B(n640), .ZN(n644) );
  OAI222D0 U385 ( .A1(n752), .A2(n751), .B1(n750), .B2(n67), .C1(n436), .C2(
        n748), .ZN(n428) );
  OAI222D0 U386 ( .A1(n757), .A2(n756), .B1(n755), .B2(n754), .C1(n442), .C2(
        n753), .ZN(n429) );
  ND4D1 U387 ( .A1(n504), .A2(n503), .A3(n502), .A4(n501), .ZN(d[6]) );
  NR4D0 U388 ( .A1(n500), .A2(n499), .A3(n515), .A4(n516), .ZN(n501) );
  NR3D0 U389 ( .A1(n732), .A2(n438), .A3(n603), .ZN(n640) );
  NR4D0 U390 ( .A1(n436), .A2(n823), .A3(n763), .A4(n769), .ZN(n570) );
  OAI221D0 U391 ( .A1(n732), .A2(n721), .B1(n443), .B2(n777), .C(n720), .ZN(
        n727) );
  ND2D1 U392 ( .A1(n439), .A2(n808), .ZN(n759) );
  NR3D0 U393 ( .A1(n732), .A2(n437), .A3(n759), .ZN(n527) );
  OAI222D0 U394 ( .A1(n568), .A2(n768), .B1(n777), .B2(n567), .C1(n566), .C2(
        n770), .ZN(n571) );
  NR4D0 U395 ( .A1(n453), .A2(n452), .A3(n526), .A4(n451), .ZN(n454) );
  OAI222D0 U396 ( .A1(n740), .A2(n550), .B1(n635), .B2(n712), .C1(n741), .C2(
        n679), .ZN(n453) );
  INVD1 U397 ( .I(n767), .ZN(n826) );
  ND2D1 U398 ( .A1(n439), .A2(n440), .ZN(n696) );
  INVD1 U399 ( .I(n770), .ZN(n827) );
  ND2D1 U400 ( .A1(n436), .A2(a[2]), .ZN(n754) );
  NR2D1 U401 ( .A1(n753), .A2(n436), .ZN(n705) );
  ND2D1 U402 ( .A1(a[2]), .A2(n439), .ZN(n739) );
  ND2D1 U403 ( .A1(n437), .A2(n439), .ZN(n679) );
  OAI221D0 U404 ( .A1(n450), .A2(n635), .B1(n766), .B2(n725), .C(n449), .ZN(
        n456) );
  AOI221D0 U405 ( .A1(n785), .A2(n803), .B1(n790), .B2(n818), .C(n587), .ZN(
        n588) );
  AOI222D0 U406 ( .A1(n791), .A2(n810), .B1(n812), .B2(n793), .C1(n795), .C2(
        n439), .ZN(n589) );
  ND2D1 U407 ( .A1(n439), .A2(n823), .ZN(n505) );
  OAI222D0 U408 ( .A1(n629), .A2(n441), .B1(n603), .B2(n596), .C1(n437), .C2(
        n714), .ZN(n601) );
  OAI222D0 U409 ( .A1(n770), .A2(n77), .B1(n769), .B2(n768), .C1(n767), .C2(
        n766), .ZN(n771) );
  INVD1 U410 ( .I(n630), .ZN(n842) );
  OAI222D0 U411 ( .A1(n635), .A2(n716), .B1(n584), .B2(n725), .C1(n629), .C2(
        n658), .ZN(n477) );
  INR2D0 U412 ( .A1(n517), .B1(n658), .ZN(n704) );
  NR4D0 U413 ( .A1(n763), .A2(n751), .A3(n658), .A4(n437), .ZN(n733) );
  NR2D1 U414 ( .A1(n700), .A2(n703), .ZN(n711) );
  OAI22D0 U415 ( .A1(n67), .A2(n746), .B1(n648), .B2(n732), .ZN(n514) );
  NR2XD0 U416 ( .A1(n437), .A2(n439), .ZN(n675) );
  INVD1 U417 ( .I(n738), .ZN(n786) );
  OA222D0 U418 ( .A1(n741), .A2(n740), .B1(n739), .B2(n738), .C1(n743), .C2(
        n737), .Z(n752) );
  OAI22D1 U419 ( .A1(n737), .A2(n67), .B1(n595), .B2(n738), .ZN(n602) );
  OAI32D1 U420 ( .A1(n578), .A2(n738), .A3(n679), .B1(n577), .B2(n759), .ZN(
        n579) );
  OAI222D0 U421 ( .A1(n442), .A2(n770), .B1(n738), .B2(n751), .C1(n745), .C2(
        n741), .ZN(n482) );
  OAI22D0 U422 ( .A1(n635), .A2(n737), .B1(n738), .B2(n766), .ZN(n494) );
  OR2D1 U423 ( .A1(n438), .A2(n823), .Z(n432) );
  INVD1 U424 ( .I(n776), .ZN(n806) );
  NR2D0 U425 ( .A1(n696), .A2(n738), .ZN(n434) );
  AOI221D0 U426 ( .A1(n792), .A2(n822), .B1(n817), .B2(n551), .C(n694), .ZN(
        n558) );
  AOI22D0 U427 ( .A1(n841), .A2(n520), .B1(n686), .B2(n519), .ZN(n521) );
  AOI221D1 U428 ( .A1(n845), .A2(n785), .B1(n848), .B2(n685), .C(n684), .ZN(
        n709) );
  AOI221D1 U429 ( .A1(n694), .A2(n847), .B1(n805), .B2(n693), .C(n692), .ZN(
        n708) );
  NR4D0 U430 ( .A1(n706), .A2(n729), .A3(n705), .A4(n704), .ZN(n707) );
  NR2D1 U431 ( .A1(n427), .A2(n786), .ZN(n608) );
  INVD1 U432 ( .I(n67), .ZN(n810) );
  NR2XD0 U433 ( .A1(n822), .A2(n818), .ZN(n667) );
  ND2D1 U434 ( .A1(n442), .A2(a[6]), .ZN(n480) );
  ND2D1 U435 ( .A1(n439), .A2(a[6]), .ZN(n770) );
  ND2D1 U436 ( .A1(a[6]), .A2(n816), .ZN(n767) );
  INVD1 U437 ( .I(n714), .ZN(n833) );
  NR3D0 U438 ( .A1(n713), .A2(n438), .A3(n828), .ZN(n651) );
  AOI32D1 U439 ( .A1(n438), .A2(n828), .A3(n804), .B1(n805), .B2(n543), .ZN(
        n545) );
  OAI22D0 U440 ( .A1(n784), .A2(n714), .B1(n445), .B2(n725), .ZN(n522) );
  OAI22D0 U441 ( .A1(n445), .A2(n714), .B1(n442), .B2(n629), .ZN(n631) );
  NR4D0 U442 ( .A1(n443), .A2(n828), .A3(n757), .A4(n67), .ZN(n689) );
  OAI21D0 U443 ( .A1(n745), .A2(n604), .B(n714), .ZN(n585) );
  NR4D0 U444 ( .A1(a[6]), .A2(n802), .A3(n721), .A4(n754), .ZN(n499) );
  OA33D0 U445 ( .A1(n700), .A2(n744), .A3(n737), .B1(n699), .B2(n698), .B3(
        n762), .Z(n701) );
  NR3D0 U446 ( .A1(n698), .A2(n816), .A3(n703), .ZN(n517) );
  OAI22D0 U447 ( .A1(a[6]), .A2(n438), .B1(n439), .B2(n751), .ZN(n543) );
  NR4D0 U448 ( .A1(n679), .A2(n746), .A3(n774), .A4(n808), .ZN(n650) );
  AOI21D0 U449 ( .A1(n769), .A2(n739), .B(n774), .ZN(n620) );
  AOI21D1 U450 ( .A1(n822), .A2(n831), .B(n840), .ZN(n659) );
  OAI22D0 U451 ( .A1(n77), .A2(n778), .B1(n777), .B2(n776), .ZN(n780) );
  NR3D0 U452 ( .A1(n505), .A2(n744), .A3(n77), .ZN(n471) );
  OAI22D0 U453 ( .A1(n740), .A2(n746), .B1(n759), .B2(n779), .ZN(n680) );
endmodule


module aes_sbox_18 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n22, n48, n59, n68, n70, n123, n148, n192, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874;

  OA222D1 U19 ( .A1(n761), .A2(n760), .B1(n759), .B2(n758), .C1(n763), .C2(
        n434), .Z(n772) );
  AN2XD1 U28 ( .A1(n734), .A2(n445), .Z(n738) );
  OA21D1 U35 ( .A1(n719), .A2(n718), .B(n717), .Z(n724) );
  OR3D1 U88 ( .A1(n687), .A2(n824), .A3(n459), .Z(n648) );
  OR4D1 U199 ( .A1(n672), .A2(n590), .A3(n534), .A4(n533), .Z(n536) );
  AN2XD1 U215 ( .A1(n535), .A2(n822), .Z(n534) );
  AN2XD1 U271 ( .A1(n548), .A2(n746), .Z(n481) );
  OAI221D1 U1 ( .A1(n59), .A2(n746), .B1(n720), .B2(n758), .C(n608), .ZN(n616)
         );
  ND2D1 U2 ( .A1(n844), .A2(n851), .ZN(n640) );
  AOI211D1 U3 ( .A1(n854), .A2(n451), .B(n653), .C(n864), .ZN(n658) );
  ND2D1 U4 ( .A1(n826), .A2(n831), .ZN(n769) );
  INVD3 U5 ( .I(n454), .ZN(n831) );
  AOI221D2 U6 ( .A1(n861), .A2(n822), .B1(n708), .B2(n816), .C(n695), .ZN(n732) );
  AOI211XD0 U7 ( .A1(n817), .A2(n835), .B(n838), .C(n711), .ZN(n712) );
  CKND2D2 U8 ( .A1(n455), .A2(n846), .ZN(n771) );
  INVD4 U9 ( .I(a[6]), .ZN(n846) );
  ND4D2 U10 ( .A1(n494), .A2(n493), .A3(n492), .A4(n491), .ZN(d[7]) );
  AOI221D2 U11 ( .A1(n475), .A2(n820), .B1(n863), .B2(n829), .C(n474), .ZN(
        n476) );
  OAI221D1 U12 ( .A1(n625), .A2(n599), .B1(n453), .B2(n788), .C(n717), .ZN(
        n541) );
  INVD2 U13 ( .I(a[5]), .ZN(n839) );
  BUFFD4 U14 ( .I(n812), .Z(n457) );
  AN2XD1 U15 ( .A1(a[6]), .A2(n851), .Z(n441) );
  BUFFD4 U16 ( .I(a[7]), .Z(n455) );
  OAI31D2 U17 ( .A1(n687), .A2(n813), .A3(n830), .B(n686), .ZN(n688) );
  AOI21D1 U18 ( .A1(n845), .A2(n441), .B(n862), .ZN(n681) );
  INVD1 U20 ( .I(n766), .ZN(n814) );
  CKND2 U21 ( .I(n455), .ZN(n851) );
  ND2D1 U22 ( .A1(n453), .A2(n839), .ZN(n760) );
  INVD1 U23 ( .I(n774), .ZN(n822) );
  NR3D1 U24 ( .A1(n438), .A2(n439), .A3(n606), .ZN(n639) );
  INVD1 U25 ( .I(n739), .ZN(n813) );
  AOI221D1 U26 ( .A1(n848), .A2(n836), .B1(n834), .B2(n586), .C(n862), .ZN(
        n509) );
  NR2D1 U27 ( .A1(n813), .A2(n70), .ZN(n705) );
  INVD1 U29 ( .I(n782), .ZN(n845) );
  ND2D1 U30 ( .A1(n820), .A2(n456), .ZN(n721) );
  NR2D1 U31 ( .A1(n831), .A2(n839), .ZN(n686) );
  NR3D0 U32 ( .A1(n442), .A2(n443), .A3(n473), .ZN(n477) );
  ND2D1 U33 ( .A1(n453), .A2(a[5]), .ZN(n701) );
  ND2D1 U34 ( .A1(n455), .A2(n839), .ZN(n742) );
  ND2D1 U36 ( .A1(a[5]), .A2(n826), .ZN(n782) );
  ND2D1 U37 ( .A1(n839), .A2(n846), .ZN(n671) );
  ND2D1 U38 ( .A1(n453), .A2(n457), .ZN(n786) );
  CKBD1 U39 ( .I(n657), .Z(n447) );
  ND2D1 U40 ( .A1(a[1]), .A2(n452), .ZN(n761) );
  INVD1 U41 ( .I(n786), .ZN(n824) );
  ND2D1 U42 ( .A1(n432), .A2(n433), .ZN(n679) );
  INVD1 U43 ( .I(n444), .ZN(n809) );
  INR4D1 U44 ( .A1(n685), .B1(n866), .B2(n683), .B3(n684), .ZN(n694) );
  BUFFD4 U45 ( .I(n808), .Z(n456) );
  INVD1 U46 ( .I(n765), .ZN(n856) );
  OAI222D0 U47 ( .A1(n766), .A2(n621), .B1(n620), .B2(n457), .C1(n619), .C2(
        n691), .ZN(n622) );
  AOI21D1 U48 ( .A1(n453), .A2(n870), .B(n830), .ZN(n784) );
  INVD1 U49 ( .I(n753), .ZN(n22) );
  INVD1 U50 ( .I(n22), .ZN(n48) );
  INVD2 U51 ( .I(n22), .ZN(n59) );
  CKND2 U52 ( .I(a[1]), .ZN(n458) );
  INVD1 U53 ( .I(n70), .ZN(n434) );
  CKAN2D1 U54 ( .A1(n451), .A2(n458), .Z(n70) );
  CKAN2D1 U55 ( .A1(a[1]), .A2(n451), .Z(n68) );
  INVD1 U56 ( .I(n68), .ZN(n444) );
  ND2D1 U57 ( .A1(a[1]), .A2(n456), .ZN(n753) );
  AN3XD1 U58 ( .A1(n676), .A2(n678), .A3(n675), .Z(n123) );
  OAI222D1 U59 ( .A1(n680), .A2(n782), .B1(n451), .B2(n572), .C1(n764), .C2(
        n571), .ZN(n573) );
  OAI22D1 U60 ( .A1(n455), .A2(n671), .B1(n764), .B2(n742), .ZN(n462) );
  NR2D1 U61 ( .A1(n476), .A2(n456), .ZN(n426) );
  AN2D1 U62 ( .A1(n451), .A2(n826), .Z(n687) );
  AOI22D1 U63 ( .A1(n842), .A2(n446), .B1(n440), .B2(n839), .ZN(n572) );
  CKND2D1 U64 ( .A1(n451), .A2(n452), .ZN(n774) );
  OAI222D1 U65 ( .A1(n658), .A2(n447), .B1(n774), .B2(n776), .C1(n656), .C2(
        n786), .ZN(n659) );
  AOI222D1 U66 ( .A1(n816), .A2(n833), .B1(n835), .B2(n818), .C1(n819), .C2(
        a[5]), .ZN(n611) );
  AOI221D1 U67 ( .A1(n828), .A2(n616), .B1(n441), .B2(n615), .C(n614), .ZN(
        n638) );
  OAI222D1 U68 ( .A1(n721), .A2(n746), .B1(n451), .B2(n552), .C1(n799), .C2(
        n788), .ZN(n553) );
  ND4D2 U69 ( .A1(n596), .A2(n595), .A3(n594), .A4(n593), .ZN(d[4]) );
  OAI222D1 U70 ( .A1(n797), .A2(n597), .B1(n789), .B2(n652), .C1(n777), .C2(
        n509), .ZN(n510) );
  ND2D0 U71 ( .A1(n456), .A2(n457), .ZN(n777) );
  ND2D3 U72 ( .A1(n456), .A2(n458), .ZN(n758) );
  BUFFD8 U73 ( .I(a[3]), .Z(n453) );
  AOI221D1 U74 ( .A1(n441), .A2(n669), .B1(n856), .B2(n668), .C(n667), .ZN(
        n676) );
  OAI222D0 U75 ( .A1(n452), .A2(n666), .B1(n665), .B2(n798), .C1(n664), .C2(
        n797), .ZN(n667) );
  NR4D1 U76 ( .A1(n644), .A2(n643), .A3(n860), .A4(n642), .ZN(n645) );
  OAI22D1 U77 ( .A1(n459), .A2(n646), .B1(n645), .B2(n434), .ZN(n647) );
  AOI221D1 U78 ( .A1(n858), .A2(n456), .B1(n868), .B2(a[1]), .C(n655), .ZN(
        n656) );
  AOI221D1 U79 ( .A1(n440), .A2(n551), .B1(n856), .B2(n550), .C(n549), .ZN(
        n552) );
  OAI222D1 U80 ( .A1(n583), .A2(n725), .B1(n582), .B2(n434), .C1(a[1]), .C2(
        n581), .ZN(n584) );
  INVD1 U81 ( .I(n679), .ZN(n857) );
  OAI221D1 U82 ( .A1(n59), .A2(n700), .B1(n760), .B2(n719), .C(n699), .ZN(n707) );
  CKND2D2 U83 ( .A1(n457), .A2(n826), .ZN(n700) );
  AOI221D1 U84 ( .A1(n708), .A2(n758), .B1(a[1]), .B2(n865), .C(n570), .ZN(
        n575) );
  ND2D2 U85 ( .A1(a[1]), .A2(n457), .ZN(n799) );
  ND2D2 U86 ( .A1(n459), .A2(n457), .ZN(n766) );
  CKND2D0 U87 ( .A1(n448), .A2(n766), .ZN(n538) );
  OAI222D1 U89 ( .A1(n766), .A2(n775), .B1(n705), .B2(n735), .C1(n704), .C2(
        n794), .ZN(n706) );
  AOI221D1 U90 ( .A1(n485), .A2(n458), .B1(n833), .B2(n484), .C(n483), .ZN(
        n492) );
  AOI221D0 U91 ( .A1(n872), .A2(n458), .B1(n854), .B2(n445), .C(n540), .ZN(
        n543) );
  OAI222D1 U92 ( .A1(n543), .A2(n789), .B1(n448), .B2(n640), .C1(n542), .C2(
        n444), .ZN(n555) );
  AO31D1 U93 ( .A1(n816), .A2(n870), .A3(n697), .B(n733), .Z(n474) );
  ND4D2 U94 ( .A1(n639), .A2(n638), .A3(n637), .A4(n636), .ZN(d[3]) );
  OAI222D1 U95 ( .A1(n448), .A2(n548), .B1(n502), .B2(n765), .C1(n501), .C2(
        n769), .ZN(n506) );
  NR4D1 U96 ( .A1(n467), .A2(n466), .A3(n544), .A4(n465), .ZN(n468) );
  AOI221D1 U97 ( .A1(n834), .A2(n870), .B1(n824), .B2(n844), .C(n541), .ZN(
        n542) );
  ND2D4 U98 ( .A1(n846), .A2(n851), .ZN(n765) );
  CKND2D1 U99 ( .A1(n452), .A2(n826), .ZN(n789) );
  AO221D1 U100 ( .A1(n814), .A2(n845), .B1(n811), .B2(n828), .C(n716), .Z(n668) );
  OA21D0 U101 ( .A1(n700), .A2(n456), .B(n629), .Z(n633) );
  INVD2 U102 ( .I(n700), .ZN(n827) );
  ND2D1 U103 ( .A1(n856), .A2(n844), .ZN(n797) );
  OAI22D1 U104 ( .A1(n468), .A2(n794), .B1(n761), .B2(n650), .ZN(n469) );
  AOI221D1 U105 ( .A1(n856), .A2(n624), .B1(n623), .B2(n456), .C(n622), .ZN(
        n637) );
  NR4D1 U106 ( .A1(n555), .A2(n556), .A3(n554), .A4(n553), .ZN(n557) );
  AOI221D1 U107 ( .A1(n811), .A2(n703), .B1(n845), .B2(n449), .C(n702), .ZN(
        n704) );
  NR3D1 U108 ( .A1(n577), .A2(n428), .A3(n427), .ZN(n595) );
  OAI222D1 U109 ( .A1(n576), .A2(n771), .B1(n575), .B2(n700), .C1(n574), .C2(
        n765), .ZN(n577) );
  AOI221D2 U110 ( .A1(n814), .A2(n836), .B1(n821), .B2(n843), .C(n780), .ZN(
        n795) );
  INVD6 U111 ( .I(n453), .ZN(n826) );
  OAI221D2 U112 ( .A1(n682), .A2(n692), .B1(n681), .B2(n680), .C(n857), .ZN(
        n684) );
  ND2D1 U113 ( .A1(n831), .A2(n839), .ZN(n783) );
  ND2D4 U114 ( .A1(a[5]), .A2(n831), .ZN(n779) );
  AOI222D1 U115 ( .A1(n820), .A2(n842), .B1(n440), .B2(n497), .C1(n815), .C2(
        n845), .ZN(n502) );
  INVD1 U116 ( .I(n571), .ZN(n815) );
  ND2D2 U117 ( .A1(n451), .A2(n457), .ZN(n739) );
  OAI222D1 U118 ( .A1(n823), .A2(n646), .B1(n568), .B2(n548), .C1(n547), .C2(
        n794), .ZN(n554) );
  AOI221D1 U119 ( .A1(n825), .A2(n586), .B1(n585), .B2(n834), .C(n584), .ZN(
        n594) );
  ND2D2 U120 ( .A1(n816), .A2(n456), .ZN(n568) );
  ND2D1 U121 ( .A1(n863), .A2(n456), .ZN(n652) );
  AOI221D1 U122 ( .A1(n441), .A2(n511), .B1(n815), .B2(n524), .C(n510), .ZN(
        n520) );
  AOI221D1 U123 ( .A1(n70), .A2(n698), .B1(n697), .B2(n440), .C(n696), .ZN(
        n699) );
  AOI32D0 U124 ( .A1(a[5]), .A2(n456), .A3(n829), .B1(n840), .B2(n648), .ZN(
        n649) );
  ND2D0 U125 ( .A1(n452), .A2(a[5]), .ZN(n759) );
  CKND2D1 U126 ( .A1(a[5]), .A2(n455), .ZN(n718) );
  CKND2D0 U127 ( .A1(a[5]), .A2(n846), .ZN(n523) );
  ND2D0 U128 ( .A1(a[5]), .A2(a[6]), .ZN(n790) );
  CKND2D1 U129 ( .A1(a[5]), .A2(n851), .ZN(n722) );
  NR2XD0 U130 ( .A1(n453), .A2(a[5]), .ZN(n697) );
  CKND1 U131 ( .I(n739), .ZN(n449) );
  OA221D1 U132 ( .A1(n700), .A2(n690), .B1(n689), .B2(n799), .C(n688), .Z(n450) );
  AOI221D1 U133 ( .A1(n871), .A2(n456), .B1(n863), .B2(n820), .C(n647), .ZN(
        n678) );
  OAI22D1 U134 ( .A1(n779), .A2(n789), .B1(a[1]), .B2(n778), .ZN(n780) );
  AOI221D1 U135 ( .A1(n847), .A2(n809), .B1(n607), .B2(n458), .C(n749), .ZN(
        n608) );
  AOI221D1 U136 ( .A1(n870), .A2(n660), .B1(n867), .B2(n816), .C(n659), .ZN(
        n677) );
  CKAN2D1 U137 ( .A1(a[1]), .A2(n479), .Z(n148) );
  CKAN2D1 U138 ( .A1(n838), .A2(n848), .Z(n192) );
  NR3D1 U139 ( .A1(n148), .A2(n192), .A3(n478), .ZN(n493) );
  NR2D0 U140 ( .A1(n477), .A2(n763), .ZN(n424) );
  NR2D0 U141 ( .A1(n701), .A2(n528), .ZN(n425) );
  OR3D1 U142 ( .A1(n424), .A2(n425), .A3(n426), .Z(n478) );
  ND2D1 U143 ( .A1(n453), .A2(n831), .ZN(n763) );
  CKND2D0 U144 ( .A1(n811), .A2(n870), .ZN(n528) );
  AOI211XD0 U145 ( .A1(n870), .A2(n507), .B(n506), .C(n505), .ZN(n521) );
  OAI222D1 U146 ( .A1(n795), .A2(n794), .B1(n453), .B2(n852), .C1(n793), .C2(
        n456), .ZN(n801) );
  INVD2 U147 ( .I(n799), .ZN(n816) );
  ND2D1 U148 ( .A1(n453), .A2(n459), .ZN(n692) );
  INVD1 U149 ( .I(a[1]), .ZN(n459) );
  OA221D1 U150 ( .A1(n760), .A2(n59), .B1(n769), .B2(n680), .C(n450), .Z(n693)
         );
  CKAN2D1 U151 ( .A1(n451), .A2(n579), .Z(n427) );
  CKAN2D1 U152 ( .A1(n441), .A2(n578), .Z(n428) );
  OR2D0 U153 ( .A1(a[1]), .A2(n790), .Z(n429) );
  OR2D0 U154 ( .A1(n758), .A2(n771), .Z(n430) );
  OR2D0 U155 ( .A1(n765), .A2(n761), .Z(n431) );
  ND3D1 U156 ( .A1(n429), .A2(n430), .A3(n431), .ZN(n500) );
  AOI211XD0 U157 ( .A1(n853), .A2(n821), .B(n500), .C(n499), .ZN(n501) );
  OR2D0 U158 ( .A1(n737), .A2(n766), .Z(n432) );
  OR2XD1 U159 ( .A1(n457), .A2(n744), .Z(n433) );
  ND2D1 U160 ( .A1(n842), .A2(n441), .ZN(n737) );
  AOI211XD0 U161 ( .A1(n874), .A2(n821), .B(n495), .C(n679), .ZN(n522) );
  AOI221D1 U162 ( .A1(n856), .A2(n471), .B1(n470), .B2(n456), .C(n469), .ZN(
        n494) );
  NR4D1 U163 ( .A1(n801), .A2(n802), .A3(n803), .A4(n800), .ZN(n804) );
  OAI33D0 U164 ( .A1(n769), .A2(n457), .A3(n742), .B1(n671), .B2(a[1]), .B3(
        n670), .ZN(n674) );
  CKND0 U165 ( .I(n742), .ZN(n869) );
  AOI221D1 U166 ( .A1(n834), .A2(n810), .B1(n843), .B2(n820), .C(n573), .ZN(
        n574) );
  AOI22D1 U167 ( .A1(n816), .A2(n848), .B1(n824), .B2(n831), .ZN(n785) );
  ND4D2 U168 ( .A1(n732), .A2(n730), .A3(n731), .A4(n729), .ZN(d[1]) );
  OAI222D1 U169 ( .A1(n451), .A2(n694), .B1(n693), .B2(n765), .C1(n692), .C2(
        n691), .ZN(n695) );
  NR2D0 U170 ( .A1(n447), .A2(n650), .ZN(n435) );
  NR2D0 U171 ( .A1(n605), .A2(n604), .ZN(n436) );
  NR2D0 U172 ( .A1(n771), .A2(n603), .ZN(n437) );
  OR3D1 U173 ( .A1(n435), .A2(n436), .A3(n437), .Z(n606) );
  CKAN2D1 U174 ( .A1(n815), .A2(n861), .Z(n438) );
  CKAN2D1 U175 ( .A1(n809), .A2(n874), .Z(n439) );
  ND2D1 U176 ( .A1(n840), .A2(n859), .ZN(n650) );
  ND2D0 U177 ( .A1(n686), .A2(n859), .ZN(n604) );
  CKND0 U178 ( .I(n798), .ZN(n874) );
  CKAN2D1 U179 ( .A1(n452), .A2(n459), .Z(n440) );
  BUFFD6 U180 ( .I(a[2]), .Z(n452) );
  CKAN2D1 U181 ( .A1(n814), .A2(n869), .Z(n442) );
  CKAN2D1 U182 ( .A1(n822), .A2(n849), .Z(n443) );
  AO21D0 U183 ( .A1(n70), .A2(n847), .B(n749), .Z(n473) );
  CKND1 U184 ( .I(n68), .ZN(n445) );
  ND2D2 U185 ( .A1(n455), .A2(a[6]), .ZN(n720) );
  ND2D0 U186 ( .A1(a[6]), .A2(n851), .ZN(n794) );
  CKND2D1 U187 ( .A1(n677), .A2(n123), .ZN(d[2]) );
  AOI21D0 U188 ( .A1(n832), .A2(n873), .B(n860), .ZN(n582) );
  AOI21D1 U189 ( .A1(n872), .A2(n446), .B(n866), .ZN(n581) );
  CKND2D0 U190 ( .A1(n453), .A2(n452), .ZN(n657) );
  OAI22D0 U191 ( .A1(n758), .A2(n722), .B1(n654), .B2(n48), .ZN(n655) );
  CKND2D0 U192 ( .A1(n452), .A2(n59), .ZN(n751) );
  AOI221D1 U193 ( .A1(n867), .A2(n809), .B1(n870), .B2(n707), .C(n706), .ZN(
        n731) );
  NR2D0 U194 ( .A1(n641), .A2(n445), .ZN(n716) );
  ND2D0 U195 ( .A1(n455), .A2(n512), .ZN(n515) );
  CKND2D1 U196 ( .A1(n787), .A2(n742), .ZN(n586) );
  ND2D1 U197 ( .A1(n824), .A2(a[1]), .ZN(n597) );
  ND2D0 U198 ( .A1(n834), .A2(n873), .ZN(n775) );
  NR2D0 U200 ( .A1(n820), .A2(n809), .ZN(n629) );
  NR2D0 U201 ( .A1(n449), .A2(n810), .ZN(n630) );
  AOI221D1 U202 ( .A1(n716), .A2(n869), .B1(n446), .B2(n715), .C(n714), .ZN(
        n730) );
  CKND2D0 U203 ( .A1(n796), .A2(n700), .ZN(n537) );
  CKND2D0 U204 ( .A1(n764), .A2(n759), .ZN(n564) );
  CKND2D0 U205 ( .A1(n841), .A2(n859), .ZN(n612) );
  ND2D0 U206 ( .A1(n457), .A2(n831), .ZN(n567) );
  ND2D0 U207 ( .A1(n451), .A2(n440), .ZN(n743) );
  BUFFD4 U208 ( .I(a[4]), .Z(n454) );
  CKND0 U209 ( .I(n788), .ZN(n871) );
  AOI22D0 U210 ( .A1(n872), .A2(n816), .B1(n829), .B2(n858), .ZN(n562) );
  ND2D0 U211 ( .A1(n828), .A2(a[1]), .ZN(n734) );
  NR2D0 U212 ( .A1(n651), .A2(n736), .ZN(n755) );
  CKND2D0 U213 ( .A1(n873), .A2(n836), .ZN(n798) );
  ND2D0 U214 ( .A1(n842), .A2(n870), .ZN(n691) );
  ND2D0 U216 ( .A1(n824), .A2(n865), .ZN(n580) );
  ND2D0 U217 ( .A1(n847), .A2(n836), .ZN(n548) );
  CKND2D0 U218 ( .A1(n833), .A2(n856), .ZN(n685) );
  NR2D0 U219 ( .A1(n733), .A2(n868), .ZN(n740) );
  NR2D0 U220 ( .A1(n872), .A2(n858), .ZN(n472) );
  CKND2D0 U221 ( .A1(n449), .A2(n844), .ZN(n661) );
  CKND2D0 U222 ( .A1(n796), .A2(n568), .ZN(n569) );
  NR2D0 U223 ( .A1(n765), .A2(n783), .ZN(n708) );
  NR2XD0 U224 ( .A1(n854), .A2(n865), .ZN(n682) );
  AOI22D0 U225 ( .A1(n863), .A2(n538), .B1(n708), .B2(n537), .ZN(n539) );
  NR2D0 U226 ( .A1(n824), .A2(n818), .ZN(n461) );
  AOI22D0 U227 ( .A1(n841), .A2(n440), .B1(n816), .B2(n843), .ZN(n460) );
  CKND2D0 U228 ( .A1(n743), .A2(n59), .ZN(n602) );
  OAI32D0 U229 ( .A1(n571), .A2(n771), .A3(n760), .B1(n529), .B2(n528), .ZN(
        n530) );
  NR2D0 U230 ( .A1(n844), .A2(n824), .ZN(n529) );
  NR2D0 U231 ( .A1(n837), .A2(n842), .ZN(n617) );
  CKND2D1 U232 ( .A1(n504), .A2(n503), .ZN(n505) );
  OAI31D0 U233 ( .A1(n59), .A2(n835), .A3(n765), .B(n752), .ZN(n757) );
  AOI31D0 U234 ( .A1(n859), .A2(n751), .A3(n835), .B(n750), .ZN(n752) );
  OAI31D0 U235 ( .A1(n826), .A2(n817), .A3(n822), .B(n708), .ZN(n504) );
  AOI22D0 U236 ( .A1(n456), .A2(n829), .B1(n826), .B2(n818), .ZN(n605) );
  NR2D0 U237 ( .A1(n849), .A2(n859), .ZN(n654) );
  OAI21D0 U238 ( .A1(n764), .A2(n625), .B(n650), .ZN(n524) );
  CKND0 U239 ( .I(n764), .ZN(n835) );
  NR2D0 U240 ( .A1(n456), .A2(n773), .ZN(n756) );
  CKND0 U241 ( .I(n701), .ZN(n843) );
  AOI22D0 U242 ( .A1(n850), .A2(n440), .B1(n821), .B2(n849), .ZN(n482) );
  OAI22D0 U243 ( .A1(n482), .A2(n725), .B1(n481), .B2(n774), .ZN(n483) );
  AOI31D0 U244 ( .A1(n746), .A2(n745), .A3(n744), .B(n743), .ZN(n747) );
  AOI22D0 U245 ( .A1(n848), .A2(n762), .B1(n850), .B2(n440), .ZN(n770) );
  CKND2D0 U246 ( .A1(n777), .A2(n774), .ZN(n762) );
  CKND2D0 U247 ( .A1(n697), .A2(n859), .ZN(n646) );
  CKND2D0 U248 ( .A1(n810), .A2(n826), .ZN(n736) );
  CKND0 U249 ( .I(n718), .ZN(n873) );
  CKND2D0 U250 ( .A1(n843), .A2(n859), .ZN(n776) );
  CKND2D0 U251 ( .A1(n842), .A2(n458), .ZN(n690) );
  CKND2D0 U252 ( .A1(n834), .A2(n859), .ZN(n621) );
  OAI21D0 U253 ( .A1(n451), .A2(n701), .B(n763), .ZN(n497) );
  AOI21D0 U254 ( .A1(n819), .A2(n856), .B(n585), .ZN(n526) );
  MAOI22D0 U255 ( .A1(n868), .A2(n826), .B1(n641), .B2(n787), .ZN(n527) );
  CKND0 U256 ( .I(n781), .ZN(n852) );
  NR2XD0 U257 ( .A1(n792), .A2(n791), .ZN(n793) );
  NR2D0 U258 ( .A1(n822), .A2(n820), .ZN(n480) );
  AOI21D0 U259 ( .A1(n834), .A2(n869), .B(n710), .ZN(n516) );
  CKND0 U260 ( .I(n751), .ZN(n823) );
  AOI31D0 U261 ( .A1(n454), .A2(n846), .A3(n824), .B(n710), .ZN(n486) );
  CKND2D0 U262 ( .A1(n446), .A2(n831), .ZN(n618) );
  NR2XD0 U263 ( .A1(n810), .A2(n440), .ZN(n665) );
  AOI21D0 U264 ( .A1(n868), .A2(n829), .B(n710), .ZN(n713) );
  AOI21D0 U265 ( .A1(n867), .A2(a[1]), .B(n708), .ZN(n709) );
  ND4D0 U266 ( .A1(n70), .A2(n848), .A3(n454), .A4(n455), .ZN(n741) );
  OAI211D0 U267 ( .A1(n718), .A2(n692), .B(n563), .C(n562), .ZN(n579) );
  OAI211D0 U268 ( .A1(n567), .A2(n445), .B(n566), .C(n565), .ZN(n578) );
  NR2D0 U269 ( .A1(n868), .A2(n708), .ZN(n464) );
  CKND2D0 U270 ( .A1(n701), .A2(n763), .ZN(n703) );
  OAI22D0 U272 ( .A1(n799), .A2(n798), .B1(n797), .B2(n796), .ZN(n800) );
  AOI21D0 U273 ( .A1(n700), .A2(n599), .B(n434), .ZN(n465) );
  AOI33D0 U274 ( .A1(n627), .A2(n846), .A3(n816), .B1(n865), .B2(n826), .B3(
        n811), .ZN(n628) );
  OAI31D0 U275 ( .A1(n761), .A2(n790), .A3(n763), .B(n628), .ZN(n635) );
  OAI33D0 U276 ( .A1(n671), .A2(n451), .A3(n457), .B1(n498), .B2(n742), .B3(
        n774), .ZN(n499) );
  CKND0 U277 ( .I(n625), .ZN(n853) );
  ND2D0 U278 ( .A1(n452), .A2(n459), .ZN(n680) );
  NR2D0 U279 ( .A1(n817), .A2(n819), .ZN(n589) );
  CKND2D0 U280 ( .A1(n445), .A2(n826), .ZN(n588) );
  NR2D0 U281 ( .A1(n745), .A2(n453), .ZN(n710) );
  NR2D0 U282 ( .A1(n773), .A2(n451), .ZN(n727) );
  AOI22D0 U283 ( .A1(n820), .A2(n451), .B1(a[1]), .B2(n446), .ZN(n496) );
  OAI21D0 U284 ( .A1(n724), .A2(n59), .B(n723), .ZN(n728) );
  CKND2D0 U285 ( .A1(n454), .A2(n457), .ZN(n599) );
  AOI21D0 U286 ( .A1(n858), .A2(n446), .B(n767), .ZN(n768) );
  CKND2D1 U287 ( .A1(n611), .A2(n610), .ZN(n615) );
  NR2D0 U288 ( .A1(n822), .A2(n453), .ZN(n632) );
  NR2D0 U289 ( .A1(n454), .A2(n846), .ZN(n475) );
  CKBD4 U290 ( .I(a[0]), .Z(n451) );
  INVD1 U291 ( .I(n691), .ZN(n872) );
  INVD1 U292 ( .I(n797), .ZN(n858) );
  INVD1 U293 ( .I(n613), .ZN(n838) );
  INVD1 U294 ( .I(n580), .ZN(n866) );
  INVD1 U295 ( .I(n597), .ZN(n825) );
  AOI222D0 U296 ( .A1(n820), .A2(n836), .B1(n834), .B2(n449), .C1(n843), .C2(
        n440), .ZN(n565) );
  INVD1 U297 ( .I(n59), .ZN(n811) );
  INVD1 U298 ( .I(n604), .ZN(n868) );
  NR2D1 U299 ( .A1(n446), .A2(n835), .ZN(n670) );
  INVD1 U300 ( .I(n650), .ZN(n867) );
  INVD1 U301 ( .I(n777), .ZN(n818) );
  INVD1 U302 ( .I(n651), .ZN(n865) );
  INVD1 U303 ( .I(n737), .ZN(n854) );
  INVD1 U304 ( .I(n783), .ZN(n840) );
  INVD1 U305 ( .I(n646), .ZN(n861) );
  ND2D1 U306 ( .A1(n809), .A2(n837), .ZN(n613) );
  INVD1 U307 ( .I(n568), .ZN(n817) );
  INVD1 U308 ( .I(n721), .ZN(n821) );
  INVD1 U309 ( .I(n745), .ZN(n863) );
  ND2D1 U310 ( .A1(n832), .A2(n848), .ZN(n717) );
  INVD1 U311 ( .I(n612), .ZN(n862) );
  INVD1 U312 ( .I(n567), .ZN(n832) );
  INVD1 U313 ( .I(n621), .ZN(n860) );
  INVD1 U314 ( .I(n652), .ZN(n864) );
  OAI222D0 U315 ( .A1(n766), .A2(n701), .B1(n496), .B2(n779), .C1(a[1]), .C2(
        n764), .ZN(n507) );
  AOI21D1 U316 ( .A1(n827), .A2(a[1]), .B(n817), .ZN(n598) );
  OAI222D0 U317 ( .A1(n448), .A2(n763), .B1(n705), .B2(n701), .C1(n769), .C2(
        n568), .ZN(n546) );
  AOI221D0 U318 ( .A1(n817), .A2(n845), .B1(n840), .B2(n569), .C(n716), .ZN(
        n576) );
  OAI222D0 U319 ( .A1(n759), .A2(n445), .B1(n783), .B2(n597), .C1(n764), .C2(
        n774), .ZN(n601) );
  OAI221D0 U320 ( .A1(n472), .A2(n789), .B1(n735), .B2(n786), .C(n580), .ZN(
        n479) );
  INVD1 U321 ( .I(n763), .ZN(n834) );
  NR2D1 U322 ( .A1(n635), .A2(n634), .ZN(n636) );
  IND4D1 U323 ( .A1(n807), .B1(n806), .B2(n805), .B3(n804), .ZN(d[0]) );
  AOI221D0 U324 ( .A1(n749), .A2(n828), .B1(n827), .B2(n748), .C(n747), .ZN(
        n806) );
  OAI222D0 U325 ( .A1(n740), .A2(n448), .B1(n738), .B2(n737), .C1(n736), .C2(
        n735), .ZN(n807) );
  NR4D0 U326 ( .A1(n757), .A2(n756), .A3(n755), .A4(n754), .ZN(n805) );
  NR4D0 U327 ( .A1(n674), .A2(n673), .A3(n672), .A4(n756), .ZN(n675) );
  AOI221D0 U328 ( .A1(n824), .A2(n855), .B1(n863), .B2(n829), .C(n560), .ZN(
        n596) );
  NR4D0 U329 ( .A1(n592), .A2(n591), .A3(n590), .A4(n754), .ZN(n593) );
  INVD1 U330 ( .I(n779), .ZN(n844) );
  ND2D1 U331 ( .A1(n697), .A2(n856), .ZN(n744) );
  INVD1 U332 ( .I(n796), .ZN(n829) );
  NR4D0 U333 ( .A1(n490), .A2(n489), .A3(n727), .A4(n488), .ZN(n491) );
  NR4D0 U334 ( .A1(n728), .A2(n750), .A3(n727), .A4(n726), .ZN(n729) );
  NR3D0 U335 ( .A1(n445), .A2(n831), .A3(n744), .ZN(n590) );
  AOI211XD0 U336 ( .A1(n841), .A2(n602), .B(n600), .C(n601), .ZN(n603) );
  ND2D1 U337 ( .A1(n441), .A2(n840), .ZN(n735) );
  AOI22D1 U338 ( .A1(n824), .A2(n844), .B1(n827), .B2(n839), .ZN(n778) );
  INVD1 U339 ( .I(n761), .ZN(n820) );
  ND3D1 U340 ( .A1(n559), .A2(n558), .A3(n557), .ZN(d[5]) );
  INR4D0 U341 ( .A1(n773), .B1(n536), .B2(n755), .B3(n726), .ZN(n558) );
  AOI211D1 U342 ( .A1(n873), .A2(n532), .B(n531), .C(n530), .ZN(n559) );
  INVD1 U343 ( .I(n671), .ZN(n848) );
  NR3D0 U344 ( .A1(n523), .A2(n764), .A3(n799), .ZN(n489) );
  INVD1 U345 ( .I(n789), .ZN(n828) );
  ND2D1 U346 ( .A1(n859), .A2(n844), .ZN(n651) );
  NR2D1 U347 ( .A1(n722), .A2(n725), .ZN(n733) );
  NR2D1 U348 ( .A1(n640), .A2(n434), .ZN(n781) );
  NR2D1 U349 ( .A1(n718), .A2(n758), .ZN(n749) );
  OAI221D0 U350 ( .A1(a[1]), .A2(n685), .B1(n736), .B2(n691), .C(n539), .ZN(
        n556) );
  INVD1 U351 ( .I(n692), .ZN(n830) );
  INVD1 U352 ( .I(n760), .ZN(n841) );
  INVD1 U353 ( .I(n719), .ZN(n837) );
  INVD1 U354 ( .I(n771), .ZN(n870) );
  ND2D1 U355 ( .A1(n842), .A2(n859), .ZN(n745) );
  INVD1 U356 ( .I(n743), .ZN(n819) );
  INVD1 U357 ( .I(n523), .ZN(n847) );
  INVD1 U358 ( .I(n626), .ZN(n842) );
  OAI222D0 U359 ( .A1(n448), .A2(n612), .B1(n746), .B2(n692), .C1(n651), .C2(
        n774), .ZN(n560) );
  OAI221D0 U360 ( .A1(n461), .A2(n626), .B1(n789), .B2(n445), .C(n460), .ZN(
        n471) );
  OAI222D0 U361 ( .A1(n742), .A2(n613), .B1(n448), .B2(n776), .C1(n629), .C2(
        n612), .ZN(n614) );
  NR4D0 U362 ( .A1(n546), .A2(n545), .A3(n544), .A4(n609), .ZN(n547) );
  NR3D0 U363 ( .A1(n59), .A2(n453), .A3(n779), .ZN(n545) );
  NR2D1 U364 ( .A1(n662), .A2(n781), .ZN(n620) );
  AOI211D1 U365 ( .A1(n830), .A2(n451), .B(n446), .C(n822), .ZN(n619) );
  OAI222D0 U366 ( .A1(n487), .A2(n722), .B1(n480), .B2(n720), .C1(n742), .C2(
        n743), .ZN(n484) );
  AOI221D0 U367 ( .A1(n809), .A2(n827), .B1(n815), .B2(n841), .C(n609), .ZN(
        n610) );
  OAI221D0 U368 ( .A1(n630), .A2(n779), .B1(n764), .B2(n774), .C(n508), .ZN(
        n511) );
  OAI222D0 U369 ( .A1(n589), .A2(n788), .B1(n797), .B2(n588), .C1(n587), .C2(
        n790), .ZN(n592) );
  AOI21D1 U370 ( .A1(n809), .A2(n663), .B(n662), .ZN(n666) );
  OAI222D0 U371 ( .A1(n633), .A2(n788), .B1(n632), .B2(n737), .C1(n631), .C2(
        n769), .ZN(n634) );
  NR3D0 U372 ( .A1(n456), .A2(n454), .A3(n701), .ZN(n609) );
  OAI221D0 U373 ( .A1(n59), .A2(n742), .B1(a[1]), .B2(n797), .C(n741), .ZN(
        n748) );
  ND4D1 U374 ( .A1(n522), .A2(n521), .A3(n520), .A4(n519), .ZN(d[6]) );
  NR4D0 U375 ( .A1(n518), .A2(n517), .A3(n533), .A4(n534), .ZN(n519) );
  NR3D0 U376 ( .A1(n59), .A2(n454), .A3(n625), .ZN(n662) );
  OAI222D0 U377 ( .A1(n777), .A2(n776), .B1(n775), .B2(n774), .C1(a[1]), .C2(
        n773), .ZN(n802) );
  OAI222D0 U378 ( .A1(n772), .A2(n771), .B1(n770), .B2(n769), .C1(n451), .C2(
        n768), .ZN(n803) );
  NR3D0 U379 ( .A1(n789), .A2(n455), .A3(n454), .ZN(n683) );
  NR4D0 U380 ( .A1(n451), .A2(n846), .A3(n783), .A4(n789), .ZN(n591) );
  ND2D1 U381 ( .A1(a[1]), .A2(n453), .ZN(n796) );
  OAI222D0 U382 ( .A1(n745), .A2(n734), .B1(n713), .B2(n456), .C1(n712), .C2(
        n787), .ZN(n714) );
  INVD1 U383 ( .I(n720), .ZN(n859) );
  INVD1 U384 ( .I(n787), .ZN(n849) );
  ND2D1 U385 ( .A1(n454), .A2(n453), .ZN(n764) );
  ND2D1 U386 ( .A1(n454), .A2(n839), .ZN(n626) );
  ND2D1 U387 ( .A1(n454), .A2(n826), .ZN(n725) );
  INVD1 U388 ( .I(n451), .ZN(n808) );
  INVD1 U389 ( .I(n452), .ZN(n812) );
  OAI222D0 U390 ( .A1(n516), .A2(n758), .B1(n831), .B2(n515), .C1(n514), .C2(
        n445), .ZN(n518) );
  INR2D1 U391 ( .A1(n775), .B1(n513), .ZN(n514) );
  ND2D1 U392 ( .A1(n814), .A2(n451), .ZN(n571) );
  OAI222D0 U393 ( .A1(n527), .A2(n434), .B1(n526), .B2(n764), .C1(n525), .C2(
        n777), .ZN(n531) );
  NR2D1 U394 ( .A1(n871), .A2(n524), .ZN(n525) );
  OAI222D0 U395 ( .A1(n651), .A2(n457), .B1(n625), .B2(n618), .C1(n453), .C2(
        n735), .ZN(n623) );
  OAI221D0 U396 ( .A1(n456), .A2(n746), .B1(n720), .B2(n445), .C(n709), .ZN(
        n715) );
  OAI22D0 U397 ( .A1(n434), .A2(n769), .B1(n617), .B2(n758), .ZN(n624) );
  OAI32D1 U398 ( .A1(n599), .A2(n758), .A3(n701), .B1(n598), .B2(n779), .ZN(
        n600) );
  INVD1 U399 ( .I(n758), .ZN(n810) );
  INVD1 U400 ( .I(n657), .ZN(n446) );
  OAI31D0 U401 ( .A1(n814), .A2(n70), .A3(n824), .B(n871), .ZN(n503) );
  AOI32D0 U402 ( .A1(n814), .A2(n456), .A3(n845), .B1(n811), .B2(n564), .ZN(
        n566) );
  AOI22D0 U403 ( .A1(n821), .A2(n869), .B1(n814), .B2(n849), .ZN(n583) );
  NR2XD0 U404 ( .A1(n818), .A2(n814), .ZN(n487) );
  AOI32D0 U405 ( .A1(n455), .A2(n831), .A3(n814), .B1(n440), .B2(n462), .ZN(
        n463) );
  INVD1 U406 ( .I(n449), .ZN(n448) );
  NR4D0 U407 ( .A1(n725), .A2(n777), .A3(n771), .A4(n839), .ZN(n750) );
  OAI33D0 U408 ( .A1(n766), .A2(n765), .A3(n764), .B1(n787), .B2(n457), .B3(
        n763), .ZN(n767) );
  OAI211D0 U409 ( .A1(n839), .A2(n769), .B(n786), .C(n764), .ZN(n698) );
  OAI211D0 U410 ( .A1(a[5]), .A2(n796), .B(n641), .C(n763), .ZN(n550) );
  OAI222D0 U411 ( .A1(n790), .A2(n799), .B1(n789), .B2(n788), .C1(n787), .C2(
        n786), .ZN(n791) );
  ND2D1 U412 ( .A1(n839), .A2(n851), .ZN(n625) );
  OAI32D0 U413 ( .A1(n782), .A2(n487), .A3(n720), .B1(n486), .B2(n59), .ZN(
        n490) );
  OAI222D0 U414 ( .A1(n774), .A2(n782), .B1(n796), .B2(n661), .C1(n763), .C2(
        n721), .ZN(n669) );
  OAI222D0 U415 ( .A1(n771), .A2(n641), .B1(n453), .B2(n640), .C1(n765), .C2(
        n782), .ZN(n644) );
  AOI21D0 U416 ( .A1(n701), .A2(n779), .B(n448), .ZN(n696) );
  NR3D0 U417 ( .A1(n839), .A2(a[1]), .A3(n739), .ZN(n544) );
  AN4D1 U418 ( .A1(n686), .A2(n829), .A3(n451), .A4(n856), .Z(n533) );
  ND2D1 U419 ( .A1(n686), .A2(n870), .ZN(n788) );
  ND3D0 U420 ( .A1(n446), .A2(n686), .A3(n856), .ZN(n773) );
  ND2D1 U421 ( .A1(n441), .A2(n686), .ZN(n746) );
  INVD1 U422 ( .I(n790), .ZN(n850) );
  OA22D0 U423 ( .A1(n790), .A2(n434), .B1(n742), .B2(n630), .Z(n631) );
  OAI221D0 U424 ( .A1(n764), .A2(n766), .B1(n725), .B2(n799), .C(n649), .ZN(
        n660) );
  INR2D1 U425 ( .A1(n535), .B1(n680), .ZN(n726) );
  NR2D1 U426 ( .A1(n523), .A2(n680), .ZN(n585) );
  NR4D0 U427 ( .A1(n783), .A2(n771), .A3(n680), .A4(n453), .ZN(n754) );
  ND2D1 U428 ( .A1(n452), .A2(n831), .ZN(n641) );
  ND2D1 U429 ( .A1(n454), .A2(n452), .ZN(n719) );
  OAI21D0 U430 ( .A1(n765), .A2(n626), .B(n735), .ZN(n607) );
  INVD0 U431 ( .I(n725), .ZN(n836) );
  OAI22D0 U432 ( .A1(n779), .A2(n700), .B1(n705), .B2(n725), .ZN(n466) );
  OAI33D0 U433 ( .A1(n447), .A2(n455), .A3(n783), .B1(n718), .B2(n457), .B3(
        n764), .ZN(n549) );
  OAI22D0 U434 ( .A1(n447), .A2(n434), .B1(n758), .B2(n786), .ZN(n512) );
  OAI222D0 U435 ( .A1(n447), .A2(n737), .B1(n605), .B2(n746), .C1(n651), .C2(
        n680), .ZN(n495) );
  OAI21D0 U436 ( .A1(n447), .A2(n745), .B(n798), .ZN(n485) );
  OAI222D0 U437 ( .A1(n760), .A2(n568), .B1(n447), .B2(n444), .C1(n761), .C2(
        n701), .ZN(n467) );
  OAI221D0 U438 ( .A1(n464), .A2(n447), .B1(n786), .B2(n746), .C(n463), .ZN(
        n470) );
  NR3D0 U439 ( .A1(n687), .A2(n814), .A3(n828), .ZN(n664) );
  OAI22D0 U440 ( .A1(n769), .A2(n766), .B1(n670), .B2(n59), .ZN(n532) );
  OAI22D0 U441 ( .A1(n760), .A2(n766), .B1(n779), .B2(n799), .ZN(n702) );
  OAI22D0 U442 ( .A1(n453), .A2(n626), .B1(n456), .B2(n625), .ZN(n627) );
  CKND2D0 U443 ( .A1(a[1]), .A2(a[6]), .ZN(n498) );
  AOI22D0 U444 ( .A1(n837), .A2(n810), .B1(n835), .B2(n452), .ZN(n587) );
  AOI31D0 U445 ( .A1(n452), .A2(n839), .A3(n70), .B(n838), .ZN(n508) );
  AOI21D0 U446 ( .A1(n745), .A2(n685), .B(n452), .ZN(n643) );
  INVD1 U447 ( .I(n735), .ZN(n855) );
  NR3D0 U448 ( .A1(n734), .A2(n454), .A3(n851), .ZN(n673) );
  AOI32D1 U449 ( .A1(n454), .A2(n851), .A3(n828), .B1(n446), .B2(n561), .ZN(
        n563) );
  OAI22D0 U450 ( .A1(n456), .A2(n735), .B1(n459), .B2(n746), .ZN(n540) );
  OAI22D0 U451 ( .A1(n459), .A2(n735), .B1(a[1]), .B2(n651), .ZN(n653) );
  NR4D0 U452 ( .A1(a[1]), .A2(n851), .A3(n777), .A4(n769), .ZN(n711) );
  OAI222D0 U453 ( .A1(n455), .A2(n785), .B1(n784), .B2(n783), .C1(n794), .C2(
        n782), .ZN(n792) );
  INVD1 U454 ( .I(n769), .ZN(n833) );
  AOI211D1 U455 ( .A1(n790), .A2(n671), .B(n599), .C(n434), .ZN(n488) );
  AOI21D0 U456 ( .A1(n626), .A2(n671), .B(n700), .ZN(n513) );
  OAI21D0 U457 ( .A1(n671), .A2(n763), .B(n744), .ZN(n551) );
  OAI22D0 U458 ( .A1(n846), .A2(n725), .B1(n831), .B2(n671), .ZN(n663) );
  ND2D1 U459 ( .A1(a[6]), .A2(n839), .ZN(n787) );
  OAI31D0 U460 ( .A1(n720), .A2(a[5]), .A3(a[1]), .B(n652), .ZN(n570) );
  NR2D0 U461 ( .A1(n845), .A2(n841), .ZN(n689) );
  NR4D0 U462 ( .A1(a[6]), .A2(n826), .A3(n742), .A4(n774), .ZN(n517) );
  OA33D0 U463 ( .A1(n722), .A2(n764), .A3(n434), .B1(n721), .B2(n720), .B3(
        n782), .Z(n723) );
  NR3D0 U464 ( .A1(n720), .A2(n839), .A3(n725), .ZN(n535) );
  OAI22D0 U465 ( .A1(a[6]), .A2(n454), .B1(a[5]), .B2(n771), .ZN(n561) );
  NR4D0 U466 ( .A1(n701), .A2(n766), .A3(n794), .A4(n831), .ZN(n672) );
  AOI21D0 U467 ( .A1(n789), .A2(n759), .B(n794), .ZN(n642) );
endmodule


module aes_sbox_17 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n64, n70, n287, n304, n305, n306, n342, n404, n405, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860;

  AN2XD1 U28 ( .A1(n716), .A2(n715), .Z(n720) );
  OA21D1 U35 ( .A1(n700), .A2(n699), .B(n698), .Z(n705) );
  OR3D1 U88 ( .A1(n667), .A2(n808), .A3(n446), .Z(n628) );
  OA21D1 U101 ( .A1(n681), .A2(n441), .B(n609), .Z(n613) );
  OR4D1 U199 ( .A1(n652), .A2(n571), .A3(n519), .A4(n518), .Z(n521) );
  AN2XD1 U215 ( .A1(n520), .A2(n806), .Z(n519) );
  AO31D1 U286 ( .A1(n799), .A2(n856), .A3(n678), .B(n714), .Z(n461) );
  ND4D2 U1 ( .A1(n507), .A2(n506), .A3(n505), .A4(n504), .ZN(d[6]) );
  NR4D1 U2 ( .A1(n786), .A2(n785), .A3(n784), .A4(n783), .ZN(n787) );
  OAI22D2 U3 ( .A1(n719), .A2(n749), .B1(n796), .B2(n726), .ZN(n659) );
  INVD2 U4 ( .I(n743), .ZN(n826) );
  NR2D2 U5 ( .A1(n830), .A2(n826), .ZN(n669) );
  CKND2D1 U6 ( .A1(n428), .A2(n436), .ZN(n555) );
  OAI222D1 U7 ( .A1(n807), .A2(n626), .B1(n552), .B2(n532), .C1(n531), .C2(
        n777), .ZN(n538) );
  NR4D0 U8 ( .A1(n530), .A2(n529), .A3(n528), .A4(n589), .ZN(n531) );
  ND2D0 U9 ( .A1(n436), .A2(n796), .ZN(n721) );
  ND4D3 U10 ( .A1(n478), .A2(n479), .A3(n477), .A4(n476), .ZN(d[7]) );
  AOI221D4 U11 ( .A1(n842), .A2(n458), .B1(n457), .B2(n441), .C(n456), .ZN(
        n479) );
  ND3D3 U12 ( .A1(n431), .A2(n432), .A3(n433), .ZN(n586) );
  NR2D1 U13 ( .A1(n699), .A2(n741), .ZN(n731) );
  OAI22D1 U14 ( .A1(n446), .A2(n626), .B1(n625), .B2(n740), .ZN(n627) );
  ND2D2 U15 ( .A1(n678), .A2(n842), .ZN(n726) );
  CKND2D1 U16 ( .A1(n441), .A2(n796), .ZN(n760) );
  OAI222D1 U17 ( .A1(n749), .A2(n601), .B1(n600), .B2(n796), .C1(n599), .C2(
        n672), .ZN(n602) );
  INR4D1 U18 ( .A1(n665), .B1(n664), .B2(n663), .B3(n852), .ZN(n675) );
  CKND2D2 U19 ( .A1(n427), .A2(n441), .ZN(n735) );
  INVD0 U20 ( .I(n735), .ZN(n795) );
  OAI221D1 U21 ( .A1(n735), .A2(n681), .B1(n743), .B2(n700), .C(n680), .ZN(
        n688) );
  ND2D2 U22 ( .A1(n445), .A2(n796), .ZN(n782) );
  INVD1 U23 ( .I(n443), .ZN(n445) );
  INVD6 U24 ( .I(a[2]), .ZN(n796) );
  OAI31D2 U25 ( .A1(n667), .A2(n797), .A3(n815), .B(n666), .ZN(n668) );
  AOI221D1 U26 ( .A1(n470), .A2(n446), .B1(n818), .B2(n469), .C(n468), .ZN(
        n477) );
  ND4D3 U27 ( .A1(n619), .A2(n618), .A3(n617), .A4(n616), .ZN(d[3]) );
  AOI221XD4 U29 ( .A1(n798), .A2(n847), .B1(n792), .B2(n860), .C(n586), .ZN(
        n619) );
  INVD2 U30 ( .I(a[6]), .ZN(n64) );
  CKND2 U31 ( .I(n64), .ZN(n70) );
  INVD1 U32 ( .I(n64), .ZN(n287) );
  CKND0 U33 ( .I(n64), .ZN(n304) );
  AOI21D2 U34 ( .A1(n811), .A2(n427), .B(n800), .ZN(n578) );
  AOI221D2 U36 ( .A1(n428), .A2(n855), .B1(n806), .B2(n834), .C(n460), .ZN(
        n464) );
  AO21D1 U37 ( .A1(n794), .A2(n832), .B(n731), .Z(n460) );
  ND2D1 U38 ( .A1(n438), .A2(n810), .ZN(n706) );
  INVD1 U39 ( .I(n701), .ZN(n845) );
  ND2D1 U40 ( .A1(n437), .A2(n796), .ZN(n769) );
  CKND3 U41 ( .I(n442), .ZN(n446) );
  INVD1 U42 ( .I(n436), .ZN(n791) );
  CKND2D0 U43 ( .A1(n445), .A2(a[2]), .ZN(n744) );
  BUFFD4 U44 ( .I(a[3]), .Z(n437) );
  CKND2D1 U45 ( .A1(n437), .A2(n816), .ZN(n746) );
  ND2D2 U46 ( .A1(n831), .A2(n836), .ZN(n748) );
  BUFFD4 U47 ( .I(a[0]), .Z(n436) );
  IND2D2 U48 ( .A1(n446), .B1(n436), .ZN(n715) );
  INVD3 U49 ( .I(n437), .ZN(n810) );
  ND2D1 U50 ( .A1(n436), .A2(a[2]), .ZN(n757) );
  INVD1 U51 ( .I(n770), .ZN(n834) );
  BUFFD1 U52 ( .I(n721), .Z(n429) );
  AOI221D0 U53 ( .A1(n857), .A2(n441), .B1(n849), .B2(n804), .C(n627), .ZN(
        n658) );
  INVD1 U54 ( .I(n659), .ZN(n843) );
  INVD1 U55 ( .I(n721), .ZN(n797) );
  OAI222D0 U56 ( .A1(n754), .A2(n621), .B1(n437), .B2(n620), .C1(n748), .C2(
        n765), .ZN(n624) );
  OAI222D0 U57 ( .A1(n778), .A2(n777), .B1(n437), .B2(n837), .C1(n776), .C2(
        n441), .ZN(n784) );
  ND2D1 U58 ( .A1(n799), .A2(n441), .ZN(n552) );
  AOI221D1 U59 ( .A1(n462), .A2(n804), .B1(n849), .B2(n814), .C(n461), .ZN(
        n463) );
  INVD3 U60 ( .I(n782), .ZN(n799) );
  INVD1 U61 ( .I(n715), .ZN(n792) );
  ND2D2 U62 ( .A1(n437), .A2(a[2]), .ZN(n637) );
  AN2XD1 U63 ( .A1(n446), .A2(n796), .Z(n428) );
  INVD1 U64 ( .I(n746), .ZN(n819) );
  AOI221D0 U65 ( .A1(n858), .A2(n446), .B1(n840), .B2(n715), .C(n525), .ZN(
        n527) );
  OA221D0 U66 ( .A1(n746), .A2(n754), .B1(n769), .B2(n762), .C(n404), .Z(n526)
         );
  MAOI22D1 U67 ( .A1(n854), .A2(n810), .B1(n621), .B2(n770), .ZN(n512) );
  BUFFD4 U68 ( .I(n791), .Z(n441) );
  INVD1 U69 ( .I(n748), .ZN(n842) );
  OAI222D0 U70 ( .A1(n429), .A2(n532), .B1(n487), .B2(n748), .C1(n486), .C2(
        n752), .ZN(n491) );
  INVD1 U71 ( .I(n754), .ZN(n856) );
  OAI222D0 U72 ( .A1(n660), .A2(n765), .B1(n436), .B2(n556), .C1(n747), .C2(
        n555), .ZN(n557) );
  ND2D2 U73 ( .A1(a[2]), .A2(n446), .ZN(n660) );
  ND2D3 U74 ( .A1(n441), .A2(n446), .ZN(n741) );
  INVD1 U75 ( .I(n741), .ZN(n793) );
  AOI211XD0 U76 ( .A1(n859), .A2(n517), .B(n516), .C(n515), .ZN(n543) );
  AOI211XD0 U77 ( .A1(n860), .A2(n805), .B(n480), .C(n659), .ZN(n507) );
  INVD1 U78 ( .I(n673), .ZN(n815) );
  ND2D1 U79 ( .A1(n437), .A2(n446), .ZN(n673) );
  OA211D0 U80 ( .A1(n699), .A2(n673), .B(n547), .C(n546), .Z(n305) );
  ND2D2 U81 ( .A1(n849), .A2(n441), .ZN(n632) );
  CKND2D2 U82 ( .A1(n439), .A2(n816), .ZN(n762) );
  INVD4 U83 ( .I(n438), .ZN(n816) );
  AOI221D2 U84 ( .A1(n812), .A2(n596), .B1(n839), .B2(n595), .C(n594), .ZN(
        n618) );
  OAI222D1 U85 ( .A1(n749), .A2(n758), .B1(n686), .B2(n717), .C1(n685), .C2(
        n777), .ZN(n687) );
  AOI221D1 U86 ( .A1(n802), .A2(n535), .B1(n842), .B2(n534), .C(n533), .ZN(
        n536) );
  OAI222D0 U87 ( .A1(n702), .A2(n728), .B1(n436), .B2(n536), .C1(n782), .C2(
        n771), .ZN(n537) );
  AOI211XD1 U89 ( .A1(n826), .A2(n582), .B(n580), .C(n581), .ZN(n583) );
  OA221D1 U90 ( .A1(n446), .A2(n434), .B1(n593), .B2(n651), .C(n435), .Z(n478)
         );
  ND2D2 U91 ( .A1(n440), .A2(n831), .ZN(n754) );
  AOI22D1 U92 ( .A1(n808), .A2(n829), .B1(n811), .B2(n824), .ZN(n761) );
  NR2XD0 U93 ( .A1(n775), .A2(n774), .ZN(n776) );
  ND2D1 U94 ( .A1(n438), .A2(n437), .ZN(n747) );
  ND2D1 U95 ( .A1(n437), .A2(n824), .ZN(n743) );
  ND2D1 U96 ( .A1(n437), .A2(n439), .ZN(n682) );
  NR2D1 U97 ( .A1(n791), .A2(n437), .ZN(n667) );
  NR2D0 U98 ( .A1(n437), .A2(n439), .ZN(n678) );
  AOI211XD0 U99 ( .A1(n800), .A2(n820), .B(n823), .C(n692), .ZN(n693) );
  OA221D1 U100 ( .A1(n441), .A2(n305), .B1(n777), .B2(n306), .C(n342), .Z(n576) );
  OA211D0 U102 ( .A1(n551), .A2(n715), .B(n550), .C(n549), .Z(n306) );
  OA222D1 U103 ( .A1(n560), .A2(n754), .B1(n559), .B2(n681), .C1(n748), .C2(
        n558), .Z(n342) );
  INVD2 U104 ( .I(n777), .ZN(n839) );
  OAI32D0 U105 ( .A1(n765), .A2(n472), .A3(n701), .B1(n471), .B2(n735), .ZN(
        n475) );
  CKND2D1 U106 ( .A1(n816), .A2(n824), .ZN(n766) );
  OAI221D1 U107 ( .A1(n735), .A2(n728), .B1(n701), .B2(n741), .C(n588), .ZN(
        n596) );
  OA221D0 U108 ( .A1(n605), .A2(n579), .B1(n437), .B2(n771), .C(n698), .Z(n404) );
  INVD2 U109 ( .I(n769), .ZN(n808) );
  INVD2 U110 ( .I(n762), .ZN(n829) );
  INVD2 U111 ( .I(n440), .ZN(n836) );
  AOI222D1 U112 ( .A1(n804), .A2(n827), .B1(n802), .B2(n482), .C1(n798), .C2(
        n830), .ZN(n487) );
  INVD2 U113 ( .I(n765), .ZN(n830) );
  ND2D1 U114 ( .A1(n810), .A2(n816), .ZN(n752) );
  OAI222D1 U115 ( .A1(n780), .A2(n577), .B1(n772), .B2(n632), .C1(n494), .C2(
        n760), .ZN(n495) );
  OAI222D1 U116 ( .A1(n638), .A2(n637), .B1(n757), .B2(n759), .C1(n636), .C2(
        n769), .ZN(n639) );
  AOI221D1 U117 ( .A1(n809), .A2(n567), .B1(n566), .B2(n819), .C(n565), .ZN(
        n575) );
  OAI222D0 U118 ( .A1(n564), .A2(n706), .B1(n563), .B2(n740), .C1(n427), .C2(
        n562), .ZN(n565) );
  CKND2D1 U119 ( .A1(n440), .A2(n824), .ZN(n724) );
  AOI211XD0 U120 ( .A1(n840), .A2(n436), .B(n633), .C(n850), .ZN(n638) );
  CKND2D1 U121 ( .A1(a[2]), .A2(n810), .ZN(n772) );
  OA222D1 U122 ( .A1(n464), .A2(n746), .B1(n682), .B2(n513), .C1(n441), .C2(
        n463), .Z(n435) );
  ND2D1 U123 ( .A1(n446), .A2(n796), .ZN(n749) );
  AOI221D1 U124 ( .A1(n689), .A2(n741), .B1(n427), .B2(n851), .C(n554), .ZN(
        n559) );
  AOI22D1 U125 ( .A1(n827), .A2(n813), .B1(n802), .B2(n824), .ZN(n556) );
  AOI221D1 U126 ( .A1(n842), .A2(n604), .B1(n603), .B2(n441), .C(n602), .ZN(
        n617) );
  OAI221D1 U127 ( .A1(n681), .A2(n670), .B1(n669), .B2(n782), .C(n668), .ZN(
        n671) );
  CKND1 U128 ( .I(n555), .ZN(n798) );
  OAI221D1 U129 ( .A1(n662), .A2(n673), .B1(n661), .B2(n660), .C(n843), .ZN(
        n664) );
  CKND2D1 U130 ( .A1(n287), .A2(n824), .ZN(n770) );
  OAI222D1 U131 ( .A1(n527), .A2(n772), .B1(n429), .B2(n620), .C1(n526), .C2(
        n715), .ZN(n539) );
  AOI221D1 U132 ( .A1(n833), .A2(n821), .B1(n819), .B2(n567), .C(n848), .ZN(
        n494) );
  AOI221D1 U133 ( .A1(n428), .A2(n821), .B1(n805), .B2(n828), .C(n763), .ZN(
        n778) );
  AOI221D1 U134 ( .A1(n853), .A2(n792), .B1(n856), .B2(n688), .C(n687), .ZN(
        n712) );
  OAI222D1 U135 ( .A1(n675), .A2(n436), .B1(n674), .B2(n748), .C1(n673), .C2(
        n672), .ZN(n676) );
  NR2XD0 U136 ( .A1(n806), .A2(n437), .ZN(n612) );
  NR2XD0 U137 ( .A1(n727), .A2(n437), .ZN(n691) );
  CKND2D0 U138 ( .A1(n427), .A2(n437), .ZN(n779) );
  ND2D2 U139 ( .A1(n796), .A2(n810), .ZN(n681) );
  INVD2 U140 ( .I(n660), .ZN(n802) );
  AOI221D1 U141 ( .A1(n819), .A2(n793), .B1(n828), .B2(n804), .C(n557), .ZN(
        n558) );
  ND2D3 U142 ( .A1(n824), .A2(n831), .ZN(n651) );
  INVD6 U143 ( .I(n439), .ZN(n824) );
  OAI33D0 U144 ( .A1(n752), .A2(n796), .A3(n724), .B1(n651), .B2(n427), .B3(
        n650), .ZN(n654) );
  CKND2D1 U145 ( .A1(n439), .A2(n810), .ZN(n765) );
  AOI221D1 U146 ( .A1(n839), .A2(n496), .B1(n798), .B2(n509), .C(n495), .ZN(
        n505) );
  ND2D2 U147 ( .A1(n827), .A2(n845), .ZN(n727) );
  INVD2 U148 ( .I(n606), .ZN(n827) );
  ND2D2 U149 ( .A1(n440), .A2(n287), .ZN(n701) );
  BUFFD6 U150 ( .I(a[7]), .Z(n440) );
  OAI31D0 U151 ( .A1(n701), .A2(n439), .A3(n427), .B(n632), .ZN(n554) );
  NR4D1 U152 ( .A1(n539), .A2(n540), .A3(n538), .A4(n537), .ZN(n541) );
  AOI221D1 U153 ( .A1(n697), .A2(n855), .B1(n813), .B2(n696), .C(n695), .ZN(
        n711) );
  ND2D2 U154 ( .A1(n839), .A2(n825), .ZN(n717) );
  ND2D2 U155 ( .A1(n304), .A2(n836), .ZN(n777) );
  CKND1 U156 ( .I(n724), .ZN(n855) );
  ND2D2 U157 ( .A1(n436), .A2(n446), .ZN(n740) );
  AOI221D1 U158 ( .A1(n844), .A2(n441), .B1(n854), .B2(n427), .C(n635), .ZN(
        n636) );
  OAI22D0 U159 ( .A1(n741), .A2(n703), .B1(n634), .B2(n735), .ZN(n635) );
  CKND1 U160 ( .I(n780), .ZN(n844) );
  AOI221D1 U161 ( .A1(n856), .A2(n640), .B1(n853), .B2(n799), .C(n639), .ZN(
        n657) );
  OA222D0 U162 ( .A1(n744), .A2(n743), .B1(n742), .B2(n741), .C1(n746), .C2(
        n740), .Z(n755) );
  OAI33D0 U163 ( .A1(n749), .A2(n748), .A3(n747), .B1(n770), .B2(n796), .B3(
        n746), .ZN(n750) );
  AOI221D1 U164 ( .A1(n847), .A2(n806), .B1(n689), .B2(n799), .C(n676), .ZN(
        n713) );
  CKND2D0 U165 ( .A1(n832), .A2(n792), .ZN(n405) );
  ND2D0 U166 ( .A1(n587), .A2(n446), .ZN(n424) );
  CKND0 U167 ( .I(n731), .ZN(n425) );
  AN3XD1 U168 ( .A1(n405), .A2(n424), .A3(n425), .Z(n588) );
  CKND2 U169 ( .I(n444), .ZN(n426) );
  INVD4 U170 ( .I(n426), .ZN(n427) );
  IND4D2 U171 ( .A1(n430), .B1(n576), .B2(n575), .B3(n574), .ZN(d[4]) );
  CKND2 U172 ( .I(n443), .ZN(n442) );
  ND2D1 U173 ( .A1(n827), .A2(n839), .ZN(n719) );
  CKND2 U174 ( .I(a[1]), .ZN(n443) );
  ND2D0 U175 ( .A1(n440), .A2(n497), .ZN(n500) );
  INVD2 U176 ( .I(n70), .ZN(n831) );
  INVD0 U177 ( .I(n443), .ZN(n444) );
  ND2D0 U178 ( .A1(n819), .A2(n845), .ZN(n601) );
  NR2D0 U179 ( .A1(n804), .A2(n792), .ZN(n609) );
  INVD1 U180 ( .I(n630), .ZN(n853) );
  AOI21D1 U181 ( .A1(n817), .A2(n859), .B(n846), .ZN(n563) );
  INVD1 U182 ( .I(n757), .ZN(n806) );
  CKND2D0 U183 ( .A1(n747), .A2(n742), .ZN(n548) );
  NR2D0 U184 ( .A1(n620), .A2(n740), .ZN(n764) );
  OAI21D0 U185 ( .A1(n747), .A2(n605), .B(n630), .ZN(n509) );
  CKND2D0 U186 ( .A1(n678), .A2(n845), .ZN(n626) );
  OAI211D0 U187 ( .A1(n439), .A2(n779), .B(n621), .C(n746), .ZN(n534) );
  AOI221D1 U188 ( .A1(n826), .A2(n795), .B1(n818), .B2(n802), .C(n671), .ZN(
        n674) );
  ND2D0 U189 ( .A1(a[2]), .A2(n816), .ZN(n621) );
  ND2D0 U190 ( .A1(n436), .A2(n802), .ZN(n725) );
  CKND2D0 U191 ( .A1(n770), .A2(n724), .ZN(n567) );
  BUFFD4 U192 ( .I(a[4]), .Z(n438) );
  BUFFD4 U193 ( .I(a[5]), .Z(n439) );
  NR2D0 U194 ( .A1(n801), .A2(n428), .ZN(n472) );
  CKND0 U195 ( .I(n771), .ZN(n857) );
  CKND0 U196 ( .I(n577), .ZN(n809) );
  OAI22D0 U197 ( .A1(n752), .A2(n749), .B1(n650), .B2(n735), .ZN(n517) );
  OAI31D0 U198 ( .A1(n428), .A2(n794), .A3(n808), .B(n857), .ZN(n488) );
  ND2D0 U200 ( .A1(n842), .A2(n829), .ZN(n780) );
  NR2XD0 U201 ( .A1(n797), .A2(n794), .ZN(n686) );
  AOI22D0 U202 ( .A1(n858), .A2(n799), .B1(n814), .B2(n844), .ZN(n546) );
  NR2D0 U203 ( .A1(n631), .A2(n718), .ZN(n737) );
  CKND2D0 U204 ( .A1(n859), .A2(n821), .ZN(n781) );
  ND2D0 U205 ( .A1(n827), .A2(n856), .ZN(n672) );
  ND2D0 U206 ( .A1(n819), .A2(n859), .ZN(n758) );
  NR2D0 U207 ( .A1(n797), .A2(n793), .ZN(n610) );
  ND2D0 U208 ( .A1(n808), .A2(n851), .ZN(n561) );
  ND2D0 U209 ( .A1(n795), .A2(n856), .ZN(n513) );
  CKND2D0 U210 ( .A1(n818), .A2(n842), .ZN(n665) );
  CKND2D0 U211 ( .A1(n832), .A2(n821), .ZN(n532) );
  NR2D0 U212 ( .A1(n714), .A2(n854), .ZN(n722) );
  CKND2D0 U213 ( .A1(n797), .A2(n829), .ZN(n641) );
  AOI211XD0 U214 ( .A1(n856), .A2(n492), .B(n491), .C(n490), .ZN(n506) );
  AOI22D0 U216 ( .A1(n805), .A2(n855), .B1(n428), .B2(n834), .ZN(n564) );
  NR2XD0 U217 ( .A1(n834), .A2(n845), .ZN(n634) );
  OAI22D0 U218 ( .A1(n441), .A2(n717), .B1(n446), .B2(n728), .ZN(n525) );
  CKND2D0 U219 ( .A1(n779), .A2(n552), .ZN(n553) );
  NR2D0 U220 ( .A1(n748), .A2(n766), .ZN(n689) );
  AOI221D0 U221 ( .A1(n839), .A2(n649), .B1(n842), .B2(n648), .C(n647), .ZN(
        n656) );
  AOI22D0 U222 ( .A1(n826), .A2(n802), .B1(n799), .B2(n828), .ZN(n447) );
  NR2D0 U223 ( .A1(n808), .A2(n801), .ZN(n448) );
  AOI22D0 U224 ( .A1(n835), .A2(n802), .B1(n805), .B2(n834), .ZN(n467) );
  CKAN2D1 U225 ( .A1(n532), .A2(n728), .Z(n466) );
  CKND2D0 U226 ( .A1(n779), .A2(n681), .ZN(n522) );
  AOI22D0 U227 ( .A1(n849), .A2(n523), .B1(n689), .B2(n522), .ZN(n524) );
  NR2XD0 U228 ( .A1(n840), .A2(n851), .ZN(n662) );
  OAI32D0 U229 ( .A1(n555), .A2(n754), .A3(n743), .B1(n514), .B2(n513), .ZN(
        n515) );
  NR2D0 U230 ( .A1(n829), .A2(n808), .ZN(n514) );
  OAI31D0 U231 ( .A1(n735), .A2(n820), .A3(n748), .B(n734), .ZN(n739) );
  OAI31D0 U232 ( .A1(n810), .A2(n800), .A3(n806), .B(n689), .ZN(n489) );
  ND2D0 U233 ( .A1(n824), .A2(n836), .ZN(n605) );
  AOI32D0 U234 ( .A1(n428), .A2(n441), .A3(n830), .B1(n795), .B2(n548), .ZN(
        n550) );
  OAI22D0 U235 ( .A1(n740), .A2(n752), .B1(n597), .B2(n741), .ZN(n604) );
  NR2D0 U236 ( .A1(n822), .A2(n827), .ZN(n597) );
  CKND2D0 U237 ( .A1(n827), .A2(n446), .ZN(n670) );
  CKND0 U238 ( .I(n747), .ZN(n820) );
  OAI22D0 U239 ( .A1(n762), .A2(n772), .B1(n427), .B2(n761), .ZN(n763) );
  CKND0 U240 ( .I(n682), .ZN(n828) );
  AOI21D0 U241 ( .A1(n606), .A2(n651), .B(n681), .ZN(n498) );
  AOI31D0 U242 ( .A1(n728), .A2(n727), .A3(n726), .B(n725), .ZN(n729) );
  AOI22D0 U243 ( .A1(n833), .A2(n745), .B1(n835), .B2(n802), .ZN(n753) );
  CKND2D0 U244 ( .A1(n760), .A2(n757), .ZN(n745) );
  ND2D0 U245 ( .A1(n796), .A2(n816), .ZN(n551) );
  OAI21D0 U246 ( .A1(n637), .A2(n727), .B(n781), .ZN(n470) );
  CKND2D0 U247 ( .A1(n793), .A2(n810), .ZN(n718) );
  CKND0 U248 ( .I(n699), .ZN(n859) );
  CKND2D0 U249 ( .A1(n829), .A2(n836), .ZN(n620) );
  NR2D0 U250 ( .A1(n858), .A2(n844), .ZN(n459) );
  CKND2D0 U251 ( .A1(n725), .A2(n735), .ZN(n582) );
  OAI21D0 U252 ( .A1(n436), .A2(n682), .B(n746), .ZN(n482) );
  NR2D0 U253 ( .A1(n806), .A2(n804), .ZN(n465) );
  AOI21D0 U254 ( .A1(n792), .A2(n643), .B(n642), .ZN(n646) );
  NR2D0 U255 ( .A1(n793), .A2(n802), .ZN(n645) );
  AOI21D0 U256 ( .A1(n819), .A2(n855), .B(n691), .ZN(n501) );
  OAI21D0 U257 ( .A1(n651), .A2(n746), .B(n726), .ZN(n535) );
  CKND2D0 U258 ( .A1(n813), .A2(n816), .ZN(n598) );
  AOI211D0 U259 ( .A1(n815), .A2(n436), .B(n813), .C(n806), .ZN(n599) );
  NR2XD0 U260 ( .A1(n642), .A2(n764), .ZN(n600) );
  AOI21D0 U261 ( .A1(n854), .A2(n814), .B(n691), .ZN(n694) );
  OAI22D0 U262 ( .A1(n743), .A2(n749), .B1(n762), .B2(n782), .ZN(n683) );
  CKND2D0 U263 ( .A1(n682), .A2(n746), .ZN(n684) );
  AOI21D0 U264 ( .A1(n853), .A2(n427), .B(n689), .ZN(n690) );
  AOI32D0 U265 ( .A1(n439), .A2(n441), .A3(n814), .B1(n825), .B2(n628), .ZN(
        n629) );
  OAI22D0 U266 ( .A1(n782), .A2(n781), .B1(n780), .B2(n779), .ZN(n783) );
  AOI31D0 U267 ( .A1(n438), .A2(n831), .A3(n808), .B(n691), .ZN(n471) );
  AOI33D0 U268 ( .A1(n607), .A2(n831), .A3(n799), .B1(n851), .B2(n810), .B3(
        n795), .ZN(n608) );
  OAI31D0 U269 ( .A1(n744), .A2(n773), .A3(n746), .B(n608), .ZN(n615) );
  AOI211D0 U270 ( .A1(n773), .A2(n651), .B(n579), .C(n740), .ZN(n473) );
  AOI211XD0 U271 ( .A1(n838), .A2(n805), .B(n485), .C(n484), .ZN(n486) );
  CKND0 U272 ( .I(n605), .ZN(n838) );
  AOI21D0 U273 ( .A1(n681), .A2(n579), .B(n740), .ZN(n452) );
  OAI21D0 U274 ( .A1(n748), .A2(n606), .B(n717), .ZN(n587) );
  NR2D0 U275 ( .A1(n800), .A2(n803), .ZN(n570) );
  CKND2D0 U276 ( .A1(n715), .A2(n810), .ZN(n569) );
  CKND0 U277 ( .I(n632), .ZN(n850) );
  OAI22D0 U278 ( .A1(n446), .A2(n717), .B1(n427), .B2(n631), .ZN(n633) );
  NR2D0 U279 ( .A1(n854), .A2(n689), .ZN(n451) );
  AOI22D0 U280 ( .A1(n804), .A2(n436), .B1(n427), .B2(n813), .ZN(n481) );
  CKND2D0 U281 ( .A1(n438), .A2(n796), .ZN(n579) );
  OAI21D0 U282 ( .A1(n705), .A2(n735), .B(n704), .ZN(n709) );
  CKND2D0 U283 ( .A1(a[2]), .A2(n735), .ZN(n733) );
  AOI22D0 U284 ( .A1(n799), .A2(n833), .B1(n808), .B2(n816), .ZN(n768) );
  CKND2D1 U285 ( .A1(n591), .A2(n590), .ZN(n595) );
  CKND2D0 U287 ( .A1(n439), .A2(n836), .ZN(n703) );
  AOI21D0 U288 ( .A1(n844), .A2(n813), .B(n750), .ZN(n751) );
  NR2XD0 U289 ( .A1(n857), .A2(n509), .ZN(n510) );
  AOI21D0 U290 ( .A1(n803), .A2(n842), .B(n566), .ZN(n511) );
  CKND2D0 U291 ( .A1(n439), .A2(n287), .ZN(n773) );
  ND2D0 U292 ( .A1(n427), .A2(n304), .ZN(n483) );
  INVD1 U293 ( .I(n672), .ZN(n858) );
  INVD1 U294 ( .I(n702), .ZN(n805) );
  INVD1 U295 ( .I(n781), .ZN(n860) );
  INVD1 U296 ( .I(n552), .ZN(n800) );
  INVD1 U297 ( .I(n561), .ZN(n852) );
  NR2D1 U298 ( .A1(n441), .A2(n756), .ZN(n738) );
  INVD1 U299 ( .I(n681), .ZN(n811) );
  INVD1 U300 ( .I(n584), .ZN(n854) );
  AO221D0 U301 ( .A1(n428), .A2(n830), .B1(n795), .B2(n812), .C(n697), .Z(n648) );
  INVD1 U302 ( .I(n631), .ZN(n851) );
  INVD1 U303 ( .I(n752), .ZN(n818) );
  INVD1 U304 ( .I(n766), .ZN(n825) );
  ND2D1 U305 ( .A1(n804), .A2(n441), .ZN(n702) );
  INVD1 U306 ( .I(n626), .ZN(n847) );
  ND2D1 U307 ( .A1(n808), .A2(n427), .ZN(n577) );
  NR2D1 U308 ( .A1(n813), .A2(n820), .ZN(n650) );
  ND2D1 U309 ( .A1(n792), .A2(n822), .ZN(n593) );
  INVD1 U310 ( .I(n760), .ZN(n801) );
  INVD1 U311 ( .I(n719), .ZN(n840) );
  ND2D1 U312 ( .A1(n812), .A2(n427), .ZN(n716) );
  INVD1 U313 ( .I(n727), .ZN(n849) );
  INVD1 U314 ( .I(n592), .ZN(n848) );
  ND2D1 U315 ( .A1(n817), .A2(n833), .ZN(n698) );
  INVD1 U316 ( .I(n551), .ZN(n817) );
  INVD1 U317 ( .I(n601), .ZN(n846) );
  INVD1 U318 ( .I(n717), .ZN(n841) );
  AOI21D1 U319 ( .A1(n858), .A2(n813), .B(n852), .ZN(n562) );
  OAI222D0 U320 ( .A1(n757), .A2(n765), .B1(n779), .B2(n641), .C1(n746), .C2(
        n702), .ZN(n649) );
  AOI221D0 U321 ( .A1(n800), .A2(n830), .B1(n825), .B2(n553), .C(n697), .ZN(
        n560) );
  AOI221D0 U322 ( .A1(n731), .A2(n812), .B1(n811), .B2(n730), .C(n729), .ZN(
        n789) );
  NR4D0 U323 ( .A1(n739), .A2(n738), .A3(n737), .A4(n736), .ZN(n788) );
  OAI221D0 U324 ( .A1(n448), .A2(n606), .B1(n772), .B2(n715), .C(n447), .ZN(
        n458) );
  AOI221D0 U325 ( .A1(n794), .A2(n679), .B1(n678), .B2(n802), .C(n677), .ZN(
        n680) );
  NR2D1 U326 ( .A1(n621), .A2(n715), .ZN(n697) );
  AOI21D1 U327 ( .A1(n830), .A2(n839), .B(n848), .ZN(n661) );
  ND4D1 U328 ( .A1(n713), .A2(n712), .A3(n711), .A4(n710), .ZN(d[1]) );
  NR4D0 U329 ( .A1(n709), .A2(n732), .A3(n708), .A4(n707), .ZN(n710) );
  NR4D0 U330 ( .A1(n475), .A2(n474), .A3(n708), .A4(n473), .ZN(n476) );
  NR2D1 U331 ( .A1(n615), .A2(n614), .ZN(n616) );
  OAI222D0 U332 ( .A1(n749), .A2(n682), .B1(n481), .B2(n762), .C1(n427), .C2(
        n747), .ZN(n492) );
  ND2D1 U333 ( .A1(n489), .A2(n488), .ZN(n490) );
  AOI31D1 U334 ( .A1(n845), .A2(n733), .A3(n820), .B(n732), .ZN(n734) );
  OAI221D0 U335 ( .A1(n427), .A2(n665), .B1(n718), .B2(n672), .C(n524), .ZN(
        n540) );
  ND4D1 U336 ( .A1(n658), .A2(n657), .A3(n656), .A4(n655), .ZN(d[2]) );
  NR4D0 U337 ( .A1(n654), .A2(n653), .A3(n652), .A4(n738), .ZN(n655) );
  NR3D0 U338 ( .A1(n715), .A2(n816), .A3(n726), .ZN(n571) );
  NR4D0 U339 ( .A1(n573), .A2(n572), .A3(n571), .A4(n736), .ZN(n574) );
  INVD1 U340 ( .I(n772), .ZN(n812) );
  OAI222D0 U341 ( .A1(n742), .A2(n715), .B1(n766), .B2(n577), .C1(n747), .C2(
        n757), .ZN(n581) );
  ND3D1 U342 ( .A1(n543), .A2(n542), .A3(n541), .ZN(d[5]) );
  INR4D0 U343 ( .A1(n756), .B1(n521), .B2(n737), .B3(n707), .ZN(n542) );
  INVD1 U344 ( .I(n651), .ZN(n833) );
  INVD1 U345 ( .I(n779), .ZN(n814) );
  NR3D0 U346 ( .A1(n508), .A2(n747), .A3(n782), .ZN(n474) );
  ND2D1 U347 ( .A1(n845), .A2(n829), .ZN(n631) );
  INVD1 U348 ( .I(n740), .ZN(n794) );
  INVD1 U349 ( .I(n744), .ZN(n804) );
  NR2D1 U350 ( .A1(n703), .A2(n706), .ZN(n714) );
  ND2D1 U351 ( .A1(n828), .A2(n845), .ZN(n759) );
  INVD1 U352 ( .I(n637), .ZN(n813) );
  INVD1 U353 ( .I(n508), .ZN(n832) );
  INVD1 U354 ( .I(n725), .ZN(n803) );
  ND2D1 U355 ( .A1(n826), .A2(n845), .ZN(n592) );
  INVD1 U356 ( .I(n700), .ZN(n822) );
  NR4D0 U357 ( .A1(n454), .A2(n453), .A3(n528), .A4(n452), .ZN(n455) );
  OAI222D0 U358 ( .A1(n743), .A2(n552), .B1(n637), .B2(n715), .C1(n744), .C2(
        n682), .ZN(n454) );
  INVD1 U359 ( .I(n733), .ZN(n807) );
  OAI222D0 U360 ( .A1(a[2]), .A2(n646), .B1(n645), .B2(n781), .C1(n644), .C2(
        n780), .ZN(n647) );
  OAI222D0 U361 ( .A1(n472), .A2(n703), .B1(n465), .B2(n701), .C1(n724), .C2(
        n725), .ZN(n469) );
  OAI222D0 U362 ( .A1(n570), .A2(n771), .B1(n780), .B2(n569), .C1(n568), .C2(
        n773), .ZN(n573) );
  OAI221D0 U363 ( .A1(n610), .A2(n762), .B1(n747), .B2(n757), .C(n493), .ZN(
        n496) );
  OAI222D0 U364 ( .A1(n727), .A2(n716), .B1(n694), .B2(n441), .C1(n693), .C2(
        n770), .ZN(n695) );
  INVD1 U365 ( .I(n764), .ZN(n837) );
  OAI222D0 U366 ( .A1(n440), .A2(n768), .B1(n767), .B2(n766), .C1(n777), .C2(
        n765), .ZN(n775) );
  OAI222D0 U367 ( .A1(n773), .A2(n782), .B1(n772), .B2(n771), .C1(n770), .C2(
        n769), .ZN(n774) );
  OAI222D0 U368 ( .A1(n512), .A2(n740), .B1(n511), .B2(n747), .C1(n510), .C2(
        n760), .ZN(n516) );
  OAI222D0 U369 ( .A1(n613), .A2(n771), .B1(n612), .B2(n719), .C1(n611), .C2(
        n752), .ZN(n614) );
  OA22D0 U370 ( .A1(n773), .A2(n740), .B1(n724), .B2(n610), .Z(n611) );
  OAI222D0 U371 ( .A1(n501), .A2(n741), .B1(n816), .B2(n500), .C1(n499), .C2(
        n715), .ZN(n503) );
  INR2D1 U372 ( .A1(n758), .B1(n498), .ZN(n499) );
  OAI221D0 U373 ( .A1(n747), .A2(n749), .B1(n706), .B2(n782), .C(n629), .ZN(
        n640) );
  NR3D0 U374 ( .A1(n441), .A2(n438), .A3(n682), .ZN(n589) );
  NR2D1 U375 ( .A1(n438), .A2(n831), .ZN(n462) );
  OAI221D0 U376 ( .A1(n735), .A2(n724), .B1(n445), .B2(n780), .C(n723), .ZN(
        n730) );
  ND2D1 U377 ( .A1(n439), .A2(n440), .ZN(n699) );
  NR4D0 U378 ( .A1(n503), .A2(n502), .A3(n518), .A4(n519), .ZN(n504) );
  NR4D0 U379 ( .A1(n624), .A2(n623), .A3(n846), .A4(n622), .ZN(n625) );
  NR2D1 U380 ( .A1(n756), .A2(n436), .ZN(n708) );
  NR3D0 U381 ( .A1(n735), .A2(n438), .A3(n605), .ZN(n642) );
  NR4D0 U382 ( .A1(n436), .A2(n831), .A3(n766), .A4(n772), .ZN(n572) );
  OAI222D0 U383 ( .A1(n755), .A2(n754), .B1(n753), .B2(n752), .C1(n436), .C2(
        n751), .ZN(n786) );
  OAI222D0 U384 ( .A1(n760), .A2(n759), .B1(n758), .B2(n757), .C1(n427), .C2(
        n756), .ZN(n785) );
  OAI222D0 U385 ( .A1(n427), .A2(n773), .B1(n741), .B2(n754), .C1(n748), .C2(
        n744), .ZN(n485) );
  ND2D1 U386 ( .A1(a[2]), .A2(n439), .ZN(n742) );
  AOI222D0 U387 ( .A1(n799), .A2(n818), .B1(n820), .B2(n801), .C1(n803), .C2(
        n439), .ZN(n591) );
  AOI221D0 U388 ( .A1(n792), .A2(n811), .B1(n798), .B2(n826), .C(n589), .ZN(
        n590) );
  ND2D1 U389 ( .A1(n438), .A2(a[2]), .ZN(n700) );
  ND2D1 U390 ( .A1(n439), .A2(n831), .ZN(n508) );
  INVD1 U391 ( .I(n773), .ZN(n835) );
  ND2D1 U392 ( .A1(n438), .A2(n824), .ZN(n606) );
  OAI222D0 U393 ( .A1(n631), .A2(n796), .B1(n605), .B2(n598), .C1(n437), .C2(
        n717), .ZN(n603) );
  OAI221D0 U394 ( .A1(n451), .A2(n637), .B1(n769), .B2(n728), .C(n450), .ZN(
        n457) );
  OAI221D0 U395 ( .A1(n441), .A2(n728), .B1(n701), .B2(n715), .C(n690), .ZN(
        n696) );
  IND4D1 U396 ( .A1(n790), .B1(n789), .B2(n788), .B3(n787), .ZN(d[0]) );
  ND2D1 U397 ( .A1(n666), .A2(n856), .ZN(n771) );
  ND2D1 U398 ( .A1(n839), .A2(n666), .ZN(n728) );
  AN4D1 U399 ( .A1(n666), .A2(n814), .A3(n436), .A4(n842), .Z(n518) );
  ND3D0 U400 ( .A1(n813), .A2(n666), .A3(n842), .ZN(n756) );
  NR2D1 U401 ( .A1(n816), .A2(n824), .ZN(n666) );
  OAI22D0 U402 ( .A1(n637), .A2(n740), .B1(n741), .B2(n769), .ZN(n497) );
  OAI211D0 U403 ( .A1(n824), .A2(n752), .B(n769), .C(n747), .ZN(n679) );
  OAI33D1 U404 ( .A1(n651), .A2(n436), .A3(n796), .B1(n483), .B2(n724), .B3(
        n757), .ZN(n484) );
  OAI33D0 U405 ( .A1(n637), .A2(n440), .A3(n766), .B1(n699), .B2(n796), .B3(
        n747), .ZN(n533) );
  OAI222D0 U406 ( .A1(n637), .A2(n719), .B1(n585), .B2(n728), .C1(n631), .C2(
        n660), .ZN(n480) );
  NR2D0 U407 ( .A1(n508), .A2(n660), .ZN(n566) );
  OAI22D0 U408 ( .A1(n437), .A2(n606), .B1(n441), .B2(n605), .ZN(n607) );
  OAI22D0 U409 ( .A1(n467), .A2(n706), .B1(n466), .B2(n757), .ZN(n468) );
  NR4D0 U410 ( .A1(n706), .A2(n760), .A3(n754), .A4(n824), .ZN(n732) );
  OAI22D0 U411 ( .A1(n831), .A2(n706), .B1(n816), .B2(n651), .ZN(n643) );
  OAI22D0 U412 ( .A1(n762), .A2(n681), .B1(n686), .B2(n706), .ZN(n453) );
  NR3D0 U413 ( .A1(n735), .A2(n437), .A3(n762), .ZN(n529) );
  AOI21D0 U414 ( .A1(n437), .A2(n856), .B(n815), .ZN(n767) );
  INVD1 U415 ( .I(n706), .ZN(n821) );
  OAI222D0 U416 ( .A1(n722), .A2(n429), .B1(n720), .B2(n719), .C1(n718), .C2(
        n717), .ZN(n790) );
  CKND2D0 U417 ( .A1(n429), .A2(n749), .ZN(n523) );
  OAI222D0 U418 ( .A1(n724), .A2(n593), .B1(n429), .B2(n759), .C1(n609), .C2(
        n592), .ZN(n594) );
  OAI222D0 U419 ( .A1(n429), .A2(n592), .B1(n728), .B2(n673), .C1(n631), .C2(
        n757), .ZN(n544) );
  AOI21D0 U420 ( .A1(n682), .A2(n762), .B(n429), .ZN(n677) );
  OAI222D0 U421 ( .A1(n429), .A2(n746), .B1(n686), .B2(n682), .C1(n752), .C2(
        n552), .ZN(n530) );
  NR3D0 U422 ( .A1(n824), .A2(n445), .A3(n429), .ZN(n528) );
  AO221D0 U423 ( .A1(n808), .A2(n841), .B1(n849), .B2(n814), .C(n544), .Z(n430) );
  AOI221D0 U424 ( .A1(n795), .A2(n684), .B1(n830), .B2(n797), .C(n683), .ZN(
        n685) );
  AOI222D0 U425 ( .A1(n804), .A2(n821), .B1(n819), .B2(n797), .C1(n828), .C2(
        n802), .ZN(n549) );
  NR3D0 U426 ( .A1(n667), .A2(n428), .A3(n812), .ZN(n644) );
  AOI22D0 U427 ( .A1(n822), .A2(n793), .B1(n820), .B2(a[2]), .ZN(n568) );
  AOI31D0 U428 ( .A1(a[2]), .A2(n824), .A3(n794), .B(n823), .ZN(n493) );
  AOI21D0 U429 ( .A1(n727), .A2(n665), .B(a[2]), .ZN(n623) );
  ND4D1 U430 ( .A1(n794), .A2(n833), .A3(n438), .A4(n440), .ZN(n723) );
  NR3D0 U431 ( .A1(n772), .A2(n440), .A3(n438), .ZN(n663) );
  AOI32D1 U432 ( .A1(n440), .A2(n816), .A3(n428), .B1(n802), .B2(n449), .ZN(
        n450) );
  OAI22D0 U433 ( .A1(n440), .A2(n651), .B1(n747), .B2(n724), .ZN(n449) );
  OR2D0 U434 ( .A1(n637), .A2(n630), .Z(n431) );
  OR2D0 U435 ( .A1(n585), .A2(n584), .Z(n432) );
  OR2XD1 U436 ( .A1(n583), .A2(n754), .Z(n433) );
  CKND2D0 U437 ( .A1(n825), .A2(n845), .ZN(n630) );
  AOI22D0 U438 ( .A1(n441), .A2(n814), .B1(n810), .B2(n801), .ZN(n585) );
  ND2D1 U439 ( .A1(n666), .A2(n845), .ZN(n584) );
  OAI32D1 U440 ( .A1(n579), .A2(n741), .A3(n682), .B1(n578), .B2(n762), .ZN(
        n580) );
  OA221D0 U441 ( .A1(n459), .A2(n772), .B1(n717), .B2(n769), .C(n561), .Z(n434) );
  INVD1 U442 ( .I(n593), .ZN(n823) );
  NR3D0 U443 ( .A1(n716), .A2(n438), .A3(n836), .ZN(n653) );
  OAI22D0 U444 ( .A1(n455), .A2(n777), .B1(n744), .B2(n630), .ZN(n456) );
  AOI32D1 U445 ( .A1(n438), .A2(n836), .A3(n812), .B1(n813), .B2(n545), .ZN(
        n547) );
  NR4D0 U446 ( .A1(n682), .A2(n749), .A3(n777), .A4(n816), .ZN(n652) );
  AOI21D0 U447 ( .A1(n772), .A2(n742), .B(n777), .ZN(n622) );
  NR4D0 U448 ( .A1(n445), .A2(n836), .A3(n760), .A4(n752), .ZN(n692) );
  INR2D1 U449 ( .A1(n520), .B1(n660), .ZN(n707) );
  NR4D0 U450 ( .A1(n766), .A2(n754), .A3(n660), .A4(n437), .ZN(n736) );
  NR4D0 U451 ( .A1(n287), .A2(n810), .A3(n724), .A4(n757), .ZN(n502) );
  OA33D0 U452 ( .A1(n703), .A2(n747), .A3(n740), .B1(n702), .B2(n701), .B3(
        n765), .Z(n704) );
  NR3D0 U453 ( .A1(n701), .A2(n824), .A3(n706), .ZN(n520) );
  OAI22D0 U454 ( .A1(n304), .A2(n438), .B1(n439), .B2(n754), .ZN(n545) );
endmodule


module aes_sbox_16 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n40, n59, n64, n65, n70, n74, n192, n203, n398, n399, n400, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868;

  AN2XD1 U28 ( .A1(n728), .A2(n727), .Z(n732) );
  OA21D1 U35 ( .A1(n712), .A2(n711), .B(n710), .Z(n717) );
  OR3D1 U88 ( .A1(n680), .A2(n817), .A3(n456), .Z(n642) );
  OR4D1 U199 ( .A1(n666), .A2(n584), .A3(n528), .A4(n527), .Z(n530) );
  AN2XD1 U215 ( .A1(n529), .A2(n815), .Z(n528) );
  AN2XD1 U271 ( .A1(n542), .A2(n740), .Z(n478) );
  AO21D1 U297 ( .A1(n805), .A2(n840), .B(n743), .Z(n470) );
  AOI21D1 U1 ( .A1(n447), .A2(n864), .B(n824), .ZN(n779) );
  OAI31D2 U2 ( .A1(n680), .A2(n441), .A3(n824), .B(n679), .ZN(n681) );
  NR2D1 U3 ( .A1(n825), .A2(n832), .ZN(n679) );
  ND2D1 U4 ( .A1(n813), .A2(n451), .ZN(n714) );
  AOI211XD2 U5 ( .A1(n834), .A2(n596), .B(n594), .C(n595), .ZN(n597) );
  OAI32D2 U6 ( .A1(n593), .A2(n753), .A3(n694), .B1(n592), .B2(n774), .ZN(n594) );
  AOI221XD4 U7 ( .A1(n808), .A2(n855), .B1(n803), .B2(n868), .C(n600), .ZN(
        n633) );
  OAI222D1 U8 ( .A1(n577), .A2(n440), .B1(n576), .B2(n752), .C1(n433), .C2(
        n575), .ZN(n578) );
  OAI221D1 U9 ( .A1(n675), .A2(n685), .B1(n674), .B2(n429), .C(n851), .ZN(n677) );
  ND2D0 U10 ( .A1(n447), .A2(n456), .ZN(n685) );
  NR2D1 U11 ( .A1(n711), .A2(n753), .ZN(n743) );
  CKND2D2 U12 ( .A1(n451), .A2(n455), .ZN(n753) );
  MAOI22D0 U13 ( .A1(n862), .A2(n819), .B1(n635), .B2(n782), .ZN(n521) );
  ND2D0 U14 ( .A1(a[6]), .A2(n832), .ZN(n782) );
  ND4D2 U15 ( .A1(n589), .A2(n590), .A3(n588), .A4(n587), .ZN(d[4]) );
  NR2XD0 U16 ( .A1(n804), .A2(n40), .ZN(n659) );
  ND2D0 U17 ( .A1(a[0]), .A2(n40), .ZN(n737) );
  NR3D1 U18 ( .A1(n74), .A2(n192), .A3(n504), .ZN(n514) );
  AOI21D2 U19 ( .A1(n820), .A2(n453), .B(n810), .ZN(n592) );
  NR4D1 U20 ( .A1(n638), .A2(n637), .A3(n854), .A4(n636), .ZN(n639) );
  AOI221D1 U21 ( .A1(n865), .A2(n451), .B1(n857), .B2(n813), .C(n641), .ZN(
        n672) );
  AOI211XD0 U22 ( .A1(n868), .A2(n814), .B(n489), .C(n673), .ZN(n516) );
  OAI22D0 U23 ( .A1(n753), .A2(n715), .B1(n648), .B2(n747), .ZN(n649) );
  CKND2D2 U24 ( .A1(n857), .A2(n451), .ZN(n646) );
  ND3D2 U25 ( .A1(n553), .A2(n552), .A3(n551), .ZN(d[5]) );
  OAI222D0 U26 ( .A1(n714), .A2(n740), .B1(a[0]), .B2(n546), .C1(n794), .C2(
        n783), .ZN(n547) );
  AOI211XD1 U27 ( .A1(n846), .A2(n814), .B(n494), .C(n493), .ZN(n495) );
  ND2D2 U29 ( .A1(n452), .A2(n819), .ZN(n693) );
  CKBD4 U30 ( .I(n807), .Z(n452) );
  OAI222D2 U31 ( .A1(n432), .A2(n644), .B1(n599), .B2(n598), .C1(n766), .C2(
        n597), .ZN(n600) );
  NR4D1 U32 ( .A1(n540), .A2(n539), .A3(n538), .A4(n603), .ZN(n541) );
  AOI221D1 U33 ( .A1(n709), .A2(n863), .B1(n822), .B2(n708), .C(n707), .ZN(
        n723) );
  ND2D2 U34 ( .A1(n839), .A2(n844), .ZN(n760) );
  INVD2 U36 ( .I(a[6]), .ZN(n839) );
  INVD2 U37 ( .I(n450), .ZN(n844) );
  CKND2 U38 ( .I(n673), .ZN(n851) );
  INR4D2 U39 ( .A1(n678), .B1(n677), .B2(n676), .B3(n860), .ZN(n687) );
  OAI222D1 U40 ( .A1(n429), .A2(n777), .B1(a[0]), .B2(n566), .C1(n759), .C2(
        n565), .ZN(n567) );
  BUFFD8 U41 ( .I(n802), .Z(n451) );
  OAI222D1 U42 ( .A1(n537), .A2(n784), .B1(n733), .B2(n634), .C1(n536), .C2(
        n727), .ZN(n549) );
  ND2D2 U43 ( .A1(n447), .A2(n452), .ZN(n781) );
  OAI222D1 U44 ( .A1(n754), .A2(n727), .B1(n778), .B2(n591), .C1(n759), .C2(
        n769), .ZN(n595) );
  CKND2D1 U45 ( .A1(n447), .A2(n825), .ZN(n758) );
  CKND2D1 U46 ( .A1(n819), .A2(n825), .ZN(n764) );
  AOI221D1 U47 ( .A1(n828), .A2(n804), .B1(n836), .B2(n813), .C(n567), .ZN(
        n568) );
  INVD1 U48 ( .I(n455), .ZN(n454) );
  ND2D1 U49 ( .A1(n825), .A2(n832), .ZN(n778) );
  CKND2D0 U50 ( .A1(n442), .A2(a[0]), .ZN(n565) );
  ND2D1 U51 ( .A1(n447), .A2(n832), .ZN(n755) );
  INVD1 U52 ( .I(n781), .ZN(n817) );
  ND2D2 U53 ( .A1(n835), .A2(n853), .ZN(n739) );
  CKBD4 U54 ( .I(a[7]), .Z(n450) );
  AOI221D0 U55 ( .A1(n850), .A2(n618), .B1(n617), .B2(n451), .C(n616), .ZN(
        n631) );
  INVD1 U56 ( .I(n685), .ZN(n824) );
  INVD1 U57 ( .I(n446), .ZN(n807) );
  AOI221D1 U58 ( .A1(n442), .A2(n439), .B1(n814), .B2(n836), .C(n775), .ZN(
        n790) );
  OAI221D0 U59 ( .A1(n747), .A2(n740), .B1(n713), .B2(n753), .C(n602), .ZN(
        n610) );
  AOI221D1 U60 ( .A1(a[0]), .A2(n573), .B1(n847), .B2(n572), .C(n571), .ZN(
        n589) );
  NR2D1 U61 ( .A1(n451), .A2(n447), .ZN(n680) );
  INVD1 U62 ( .I(n755), .ZN(n834) );
  ND2D1 U63 ( .A1(a[0]), .A2(n455), .ZN(n752) );
  CKBD1 U64 ( .I(n807), .Z(n430) );
  INVD1 U65 ( .I(n665), .ZN(n841) );
  ND2D1 U66 ( .A1(n451), .A2(n430), .ZN(n772) );
  ND2D1 U67 ( .A1(a[0]), .A2(n446), .ZN(n769) );
  INVD1 U68 ( .I(n693), .ZN(n820) );
  AOI221D0 U69 ( .A1(n866), .A2(n455), .B1(n848), .B2(n727), .C(n534), .ZN(
        n537) );
  OAI222D0 U70 ( .A1(n816), .A2(n640), .B1(n562), .B2(n542), .C1(n541), .C2(
        n789), .ZN(n548) );
  INVD1 U71 ( .I(n760), .ZN(n850) );
  INVD1 U72 ( .I(n620), .ZN(n835) );
  ND2D2 U73 ( .A1(n448), .A2(n832), .ZN(n620) );
  INVD2 U74 ( .I(n651), .ZN(n822) );
  AN2XD1 U75 ( .A1(n446), .A2(n456), .Z(n40) );
  OA22D0 U76 ( .A1(n479), .A2(n440), .B1(n478), .B2(n769), .Z(n65) );
  AOI22D1 U77 ( .A1(n843), .A2(n40), .B1(n814), .B2(n842), .ZN(n479) );
  INVD3 U78 ( .I(n794), .ZN(n809) );
  OA221D1 U79 ( .A1(n693), .A2(n683), .B1(n682), .B2(n794), .C(n681), .Z(n445)
         );
  OAI21D1 U80 ( .A1(a[0]), .A2(n694), .B(n758), .ZN(n491) );
  ND2D1 U81 ( .A1(n450), .A2(n832), .ZN(n736) );
  INVD6 U82 ( .I(n449), .ZN(n832) );
  AOI221D2 U83 ( .A1(n855), .A2(n815), .B1(n701), .B2(n809), .C(n688), .ZN(
        n725) );
  CKND2D2 U84 ( .A1(n454), .A2(n452), .ZN(n794) );
  AOI22D2 U85 ( .A1(n40), .A2(n832), .B1(n835), .B2(n822), .ZN(n566) );
  OA221D1 U86 ( .A1(n59), .A2(a[1]), .B1(n764), .B2(n64), .C(n65), .Z(n486) );
  OA21D0 U87 ( .A1(n432), .A2(n739), .B(n793), .Z(n59) );
  OA222D0 U89 ( .A1(n481), .A2(n715), .B1(n477), .B2(n713), .C1(n736), .C2(
        n737), .Z(n64) );
  CKND6 U90 ( .I(a[1]), .ZN(n455) );
  INVD2 U91 ( .I(n562), .ZN(n810) );
  NR3D1 U92 ( .A1(n203), .A2(n398), .A3(n653), .ZN(n671) );
  NR4D1 U93 ( .A1(n549), .A2(n548), .A3(n550), .A4(n547), .ZN(n551) );
  AOI211XD1 U94 ( .A1(n864), .A2(n501), .B(n500), .C(n499), .ZN(n515) );
  CKND1 U95 ( .I(n791), .ZN(n823) );
  OAI222D1 U96 ( .A1(n432), .A2(n731), .B1(n599), .B2(n740), .C1(n645), .C2(
        n429), .ZN(n489) );
  OAI22D2 U97 ( .A1(n731), .A2(n761), .B1(n430), .B2(n738), .ZN(n673) );
  CKND2D1 U98 ( .A1(n835), .A2(n847), .ZN(n731) );
  NR2D0 U99 ( .A1(n810), .A2(n812), .ZN(n583) );
  ND4D2 U100 ( .A1(n672), .A2(n671), .A3(n670), .A4(n669), .ZN(d[2]) );
  OAI22D0 U101 ( .A1(n456), .A2(n640), .B1(n639), .B2(n752), .ZN(n641) );
  OAI22D1 U102 ( .A1(n774), .A2(n784), .B1(n453), .B2(n773), .ZN(n775) );
  INVD2 U103 ( .I(n727), .ZN(n803) );
  ND2D2 U104 ( .A1(n454), .A2(a[0]), .ZN(n727) );
  AO31D0 U105 ( .A1(n809), .A2(n864), .A3(n690), .B(n726), .Z(n471) );
  OAI222D1 U106 ( .A1(n767), .A2(n766), .B1(n765), .B2(n764), .C1(a[0]), .C2(
        n763), .ZN(n798) );
  AOI221D1 U107 ( .A1(n472), .A2(n813), .B1(n857), .B2(n823), .C(n471), .ZN(
        n473) );
  AOI221D1 U108 ( .A1(n806), .A2(n696), .B1(n838), .B2(n441), .C(n695), .ZN(
        n697) );
  INVD1 U109 ( .I(n441), .ZN(n733) );
  OA221D1 U110 ( .A1(n755), .A2(n747), .B1(n764), .B2(n429), .C(n445), .Z(n686) );
  CKND2D1 U111 ( .A1(n454), .A2(n446), .ZN(n756) );
  ND2D1 U112 ( .A1(n847), .A2(n679), .ZN(n740) );
  OAI222D1 U113 ( .A1(n733), .A2(n542), .B1(n496), .B2(n760), .C1(n495), .C2(
        n764), .ZN(n500) );
  ND2D2 U114 ( .A1(n809), .A2(n451), .ZN(n562) );
  NR2XD1 U115 ( .A1(a[1]), .A2(n446), .ZN(n442) );
  AOI221D1 U116 ( .A1(n442), .A2(n863), .B1(n815), .B2(n842), .C(n470), .ZN(
        n474) );
  AOI22D1 U117 ( .A1(n814), .A2(n863), .B1(n442), .B2(n842), .ZN(n577) );
  INR2D1 U118 ( .A1(a[0]), .B1(n446), .ZN(n441) );
  BUFFD6 U119 ( .I(a[2]), .Z(n446) );
  CKND2 U120 ( .I(n442), .ZN(n761) );
  CKND2D1 U121 ( .A1(n447), .A2(n449), .ZN(n694) );
  ND2D2 U122 ( .A1(n453), .A2(n451), .ZN(n747) );
  CKND1 U123 ( .I(n455), .ZN(n453) );
  AOI221D1 U124 ( .A1(n852), .A2(n451), .B1(n862), .B2(n453), .C(n649), .ZN(
        n650) );
  OAI33D1 U125 ( .A1(n665), .A2(a[0]), .A3(n430), .B1(n492), .B2(n736), .B3(
        n769), .ZN(n493) );
  CKND1 U126 ( .I(n694), .ZN(n836) );
  ND2D1 U127 ( .A1(n446), .A2(n819), .ZN(n784) );
  OAI222D1 U128 ( .A1(n792), .A2(n591), .B1(n784), .B2(n646), .C1(n503), .C2(
        n772), .ZN(n504) );
  AOI221D1 U129 ( .A1(n847), .A2(n663), .B1(n850), .B2(n662), .C(n661), .ZN(
        n670) );
  AOI221D1 U130 ( .A1(n818), .A2(n580), .B1(n579), .B2(n828), .C(n578), .ZN(
        n588) );
  OAI32D0 U131 ( .A1(n565), .A2(n766), .A3(n755), .B1(n523), .B2(n522), .ZN(
        n524) );
  OAI22D0 U132 ( .A1(n755), .A2(n761), .B1(n774), .B2(n794), .ZN(n695) );
  OA222D0 U133 ( .A1(n756), .A2(n755), .B1(n754), .B2(n753), .C1(n758), .C2(
        n752), .Z(n767) );
  OAI222D1 U134 ( .A1(n570), .A2(n766), .B1(n693), .B2(n569), .C1(n568), .C2(
        n760), .ZN(n571) );
  OAI222D1 U135 ( .A1(n652), .A2(n432), .B1(n769), .B2(n771), .C1(n650), .C2(
        n781), .ZN(n653) );
  ND2D2 U136 ( .A1(n450), .A2(a[6]), .ZN(n713) );
  INVD4 U137 ( .I(n447), .ZN(n819) );
  NR2XD0 U138 ( .A1(n441), .A2(n805), .ZN(n698) );
  ND2D1 U139 ( .A1(n832), .A2(n839), .ZN(n665) );
  ND2D3 U140 ( .A1(n450), .A2(n839), .ZN(n766) );
  ND2D0 U141 ( .A1(n449), .A2(n839), .ZN(n517) );
  AOI211XD0 U142 ( .A1(n824), .A2(a[0]), .B(n822), .C(n815), .ZN(n613) );
  ND4D2 U143 ( .A1(n488), .A2(n487), .A3(n486), .A4(n485), .ZN(d[7]) );
  AOI221D1 U144 ( .A1(n828), .A2(n864), .B1(n817), .B2(n837), .C(n535), .ZN(
        n536) );
  AOI221D1 U145 ( .A1(n861), .A2(n803), .B1(n864), .B2(n700), .C(n699), .ZN(
        n724) );
  OAI211D0 U146 ( .A1(n832), .A2(n764), .B(n781), .C(n759), .ZN(n691) );
  ND2D0 U147 ( .A1(n817), .A2(n453), .ZN(n591) );
  IIND4D2 U148 ( .A1(n801), .A2(n70), .B1(n799), .B2(n800), .ZN(d[0]) );
  AO221D0 U149 ( .A1(n743), .A2(n821), .B1(n820), .B2(n742), .C(n741), .Z(n70)
         );
  AOI33D0 U150 ( .A1(n621), .A2(n839), .A3(n809), .B1(n859), .B2(n819), .B3(
        n806), .ZN(n622) );
  NR2XD0 U151 ( .A1(n448), .A2(n839), .ZN(n472) );
  INVD2 U152 ( .I(n789), .ZN(n847) );
  ND2D1 U153 ( .A1(a[6]), .A2(n844), .ZN(n789) );
  ND4D2 U154 ( .A1(n633), .A2(n632), .A3(n631), .A4(n630), .ZN(d[3]) );
  INVD2 U155 ( .I(n713), .ZN(n853) );
  AOI221D1 U156 ( .A1(n701), .A2(n753), .B1(n453), .B2(n859), .C(n564), .ZN(
        n569) );
  OAI31D0 U157 ( .A1(n713), .A2(n449), .A3(n453), .B(n646), .ZN(n564) );
  INVD6 U158 ( .I(n448), .ZN(n825) );
  ND2D3 U159 ( .A1(n449), .A2(n825), .ZN(n774) );
  AOI221D1 U160 ( .A1(n821), .A2(n610), .B1(n847), .B2(n609), .C(n608), .ZN(
        n632) );
  OAI222D1 U161 ( .A1(a[0]), .A2(n687), .B1(n686), .B2(n760), .C1(n685), .C2(
        n684), .ZN(n688) );
  ND4D2 U162 ( .A1(n516), .A2(n515), .A3(n514), .A4(n513), .ZN(d[6]) );
  CKAN2D1 U163 ( .A1(n847), .A2(n505), .Z(n74) );
  CKAN2D1 U164 ( .A1(n808), .A2(n518), .Z(n192) );
  CKAN2D1 U165 ( .A1(n864), .A2(n654), .Z(n203) );
  CKAN2D1 U166 ( .A1(n861), .A2(n809), .Z(n398) );
  INVD2 U167 ( .I(n766), .ZN(n864) );
  CKAN2D1 U168 ( .A1(n850), .A2(n468), .Z(n399) );
  CKAN2D1 U169 ( .A1(n467), .A2(n451), .Z(n400) );
  NR3D0 U170 ( .A1(n399), .A2(n400), .A3(n466), .ZN(n488) );
  AN2D1 U171 ( .A1(n817), .A2(n837), .Z(n424) );
  CKAN2D1 U172 ( .A1(n820), .A2(n832), .Z(n425) );
  NR2XD1 U173 ( .A1(n424), .A2(n425), .ZN(n773) );
  INVD2 U174 ( .I(n774), .ZN(n837) );
  CKND2D0 U175 ( .A1(n840), .A2(n803), .ZN(n426) );
  CKND2D0 U176 ( .A1(n601), .A2(n455), .ZN(n427) );
  CKND0 U177 ( .I(n743), .ZN(n428) );
  AN3XD1 U178 ( .A1(n426), .A2(n427), .A3(n428), .Z(n602) );
  OAI222D1 U179 ( .A1(n790), .A2(n789), .B1(n447), .B2(n845), .C1(n788), .C2(
        n451), .ZN(n796) );
  CKND2D2 U180 ( .A1(n725), .A2(n444), .ZN(d[1]) );
  NR2XD0 U181 ( .A1(n787), .A2(n786), .ZN(n788) );
  NR4D1 U182 ( .A1(n796), .A2(n797), .A3(n798), .A4(n795), .ZN(n799) );
  CKND2 U183 ( .I(n40), .ZN(n429) );
  CKND0 U184 ( .I(n651), .ZN(n431) );
  CKND2 U185 ( .I(n431), .ZN(n432) );
  ND2D1 U186 ( .A1(n447), .A2(n446), .ZN(n651) );
  ND2D0 U187 ( .A1(n446), .A2(n825), .ZN(n635) );
  ND2D0 U188 ( .A1(n446), .A2(n449), .ZN(n754) );
  CKND2D0 U189 ( .A1(n448), .A2(n446), .ZN(n712) );
  CKND2D1 U190 ( .A1(n679), .A2(n864), .ZN(n783) );
  ND2D0 U191 ( .A1(n834), .A2(n853), .ZN(n606) );
  NR2XD0 U192 ( .A1(n842), .A2(n853), .ZN(n648) );
  CKND0 U193 ( .I(n455), .ZN(n433) );
  NR3D0 U194 ( .A1(n434), .A2(n435), .A3(n475), .ZN(n487) );
  BUFFD6 U195 ( .I(a[5]), .Z(n449) );
  CKND2D0 U196 ( .A1(n827), .A2(n850), .ZN(n678) );
  CKND1 U197 ( .I(n769), .ZN(n815) );
  OAI21D0 U198 ( .A1(n717), .A2(n747), .B(n716), .ZN(n721) );
  IND2D0 U200 ( .A1(n455), .B1(n447), .ZN(n791) );
  CKAN2D1 U201 ( .A1(n433), .A2(n476), .Z(n434) );
  CKAN2D1 U202 ( .A1(n831), .A2(n841), .Z(n435) );
  NR2D0 U203 ( .A1(n474), .A2(n758), .ZN(n436) );
  NR2D0 U204 ( .A1(n694), .A2(n522), .ZN(n437) );
  NR2D0 U205 ( .A1(n473), .A2(n451), .ZN(n438) );
  OR3D1 U206 ( .A1(n436), .A2(n437), .A3(n438), .Z(n475) );
  CKND2D0 U207 ( .A1(n806), .A2(n864), .ZN(n522) );
  INVD1 U208 ( .I(n739), .ZN(n857) );
  CKND2D0 U209 ( .A1(n694), .A2(n758), .ZN(n696) );
  CKND2D0 U210 ( .A1(n791), .A2(n693), .ZN(n531) );
  CKND2D0 U211 ( .A1(n679), .A2(n853), .ZN(n598) );
  AOI21D1 U212 ( .A1(n826), .A2(n867), .B(n854), .ZN(n576) );
  ND2D0 U213 ( .A1(n835), .A2(n455), .ZN(n683) );
  INR2D0 U214 ( .A1(n770), .B1(n507), .ZN(n508) );
  NR2XD0 U216 ( .A1(n865), .A2(n518), .ZN(n519) );
  ND2D0 U217 ( .A1(n449), .A2(n844), .ZN(n715) );
  CKND2D0 U218 ( .A1(n453), .A2(a[6]), .ZN(n492) );
  BUFFD4 U219 ( .I(a[4]), .Z(n448) );
  CKND0 U220 ( .I(n591), .ZN(n818) );
  ND3D0 U221 ( .A1(n822), .A2(n679), .A3(n850), .ZN(n768) );
  CKND0 U222 ( .I(n753), .ZN(n804) );
  AOI22D0 U223 ( .A1(n866), .A2(n809), .B1(n823), .B2(n852), .ZN(n556) );
  ND2D0 U224 ( .A1(n821), .A2(n433), .ZN(n728) );
  NR2D0 U225 ( .A1(n645), .A2(n730), .ZN(n749) );
  NR2D0 U226 ( .A1(n822), .A2(n829), .ZN(n664) );
  CKND2D0 U227 ( .A1(n867), .A2(n439), .ZN(n793) );
  ND2D0 U228 ( .A1(n835), .A2(n864), .ZN(n684) );
  ND2D0 U229 ( .A1(n817), .A2(n859), .ZN(n574) );
  ND2D0 U230 ( .A1(n828), .A2(n867), .ZN(n770) );
  CKND2D0 U231 ( .A1(n840), .A2(n439), .ZN(n542) );
  NR2D0 U232 ( .A1(n726), .A2(n862), .ZN(n734) );
  CKND0 U233 ( .I(n729), .ZN(n849) );
  CKND2D0 U234 ( .A1(n737), .A2(n747), .ZN(n596) );
  NR2D0 U235 ( .A1(n866), .A2(n852), .ZN(n469) );
  AOI21D0 U236 ( .A1(n866), .A2(n822), .B(n860), .ZN(n575) );
  CKND2D0 U237 ( .A1(n441), .A2(n837), .ZN(n655) );
  OAI31D0 U238 ( .A1(n442), .A2(n805), .A3(n817), .B(n865), .ZN(n497) );
  OAI33D0 U239 ( .A1(n764), .A2(n430), .A3(n736), .B1(n665), .B2(n433), .B3(
        n664), .ZN(n668) );
  CKND2D0 U240 ( .A1(n791), .A2(n562), .ZN(n563) );
  NR2D0 U241 ( .A1(n760), .A2(n778), .ZN(n701) );
  NR2XD0 U242 ( .A1(n848), .A2(n859), .ZN(n675) );
  AOI22D0 U243 ( .A1(n857), .A2(n532), .B1(n701), .B2(n531), .ZN(n533) );
  CKND2D0 U244 ( .A1(n759), .A2(n754), .ZN(n558) );
  NR2D0 U245 ( .A1(n837), .A2(n817), .ZN(n523) );
  CKND2D0 U246 ( .A1(n772), .A2(n769), .ZN(n757) );
  OAI22D0 U247 ( .A1(n432), .A2(n752), .B1(n753), .B2(n781), .ZN(n506) );
  OAI31D0 U248 ( .A1(n747), .A2(n829), .A3(n760), .B(n746), .ZN(n751) );
  AOI31D0 U249 ( .A1(n853), .A2(n745), .A3(n829), .B(n744), .ZN(n746) );
  NR2D0 U250 ( .A1(n817), .A2(n811), .ZN(n458) );
  OAI22D0 U251 ( .A1(n456), .A2(n729), .B1(n453), .B2(n645), .ZN(n647) );
  ND2D0 U252 ( .A1(n832), .A2(n844), .ZN(n619) );
  OAI21D0 U253 ( .A1(n759), .A2(n619), .B(n644), .ZN(n518) );
  CKND0 U254 ( .I(n759), .ZN(n829) );
  OAI22D0 U255 ( .A1(n752), .A2(n764), .B1(n611), .B2(n753), .ZN(n618) );
  NR2D0 U256 ( .A1(n830), .A2(n835), .ZN(n611) );
  OAI22D0 U257 ( .A1(n774), .A2(n693), .B1(n698), .B2(n440), .ZN(n463) );
  INR2D0 U258 ( .A1(n529), .B1(n429), .ZN(n719) );
  NR2D0 U259 ( .A1(n517), .A2(n429), .ZN(n579) );
  AOI21D0 U260 ( .A1(n620), .A2(n665), .B(n693), .ZN(n507) );
  CKND2D0 U261 ( .A1(n833), .A2(n853), .ZN(n644) );
  CKND2D0 U262 ( .A1(n690), .A2(n853), .ZN(n640) );
  ND2D0 U263 ( .A1(n430), .A2(n825), .ZN(n561) );
  NR2D0 U264 ( .A1(n811), .A2(n442), .ZN(n481) );
  CKND0 U265 ( .I(n711), .ZN(n867) );
  CKND2D0 U266 ( .A1(n804), .A2(n819), .ZN(n730) );
  NR2D0 U267 ( .A1(n441), .A2(n804), .ZN(n624) );
  ND2D0 U268 ( .A1(n837), .A2(n844), .ZN(n634) );
  CKND2D0 U269 ( .A1(n836), .A2(n853), .ZN(n771) );
  CKND2D0 U270 ( .A1(n828), .A2(n853), .ZN(n615) );
  AOI21D0 U272 ( .A1(n852), .A2(n822), .B(n762), .ZN(n763) );
  CKND2D1 U273 ( .A1(n605), .A2(n604), .ZN(n609) );
  NR2D0 U274 ( .A1(n815), .A2(n813), .ZN(n477) );
  AOI21D0 U275 ( .A1(n812), .A2(n850), .B(n579), .ZN(n520) );
  AOI22D0 U276 ( .A1(n809), .A2(n841), .B1(n817), .B2(n825), .ZN(n780) );
  CKND0 U277 ( .I(n745), .ZN(n816) );
  CKND2D0 U278 ( .A1(n727), .A2(n819), .ZN(n582) );
  CKND2D0 U279 ( .A1(n822), .A2(n825), .ZN(n612) );
  NR2D0 U280 ( .A1(n656), .A2(n776), .ZN(n614) );
  CKND0 U281 ( .I(n646), .ZN(n858) );
  OAI33D0 U282 ( .A1(n432), .A2(n450), .A3(n778), .B1(n711), .B2(n430), .B3(
        n759), .ZN(n543) );
  OAI21D0 U283 ( .A1(n665), .A2(n758), .B(n738), .ZN(n545) );
  ND4D0 U284 ( .A1(n805), .A2(n841), .A3(n448), .A4(n450), .ZN(n735) );
  OAI21D0 U285 ( .A1(n760), .A2(n620), .B(n729), .ZN(n601) );
  AOI21D0 U286 ( .A1(n861), .A2(n433), .B(n701), .ZN(n702) );
  OAI211D0 U287 ( .A1(n711), .A2(n685), .B(n557), .C(n556), .ZN(n573) );
  OAI22D0 U288 ( .A1(n794), .A2(n793), .B1(n792), .B2(n791), .ZN(n795) );
  AOI21D0 U289 ( .A1(n693), .A2(n593), .B(n752), .ZN(n462) );
  OA33D0 U290 ( .A1(n715), .A2(n759), .A3(n752), .B1(n714), .B2(n713), .B3(
        n777), .Z(n716) );
  OAI32D0 U291 ( .A1(n777), .A2(n481), .A3(n713), .B1(n480), .B2(n747), .ZN(
        n484) );
  AOI31D0 U292 ( .A1(n448), .A2(n839), .A3(n817), .B(n703), .ZN(n480) );
  OAI22D0 U293 ( .A1(n450), .A2(n665), .B1(n759), .B2(n736), .ZN(n459) );
  NR2D0 U294 ( .A1(n862), .A2(n701), .ZN(n461) );
  AOI211D0 U295 ( .A1(n785), .A2(n665), .B(n593), .C(n752), .ZN(n482) );
  CKND0 U296 ( .I(n619), .ZN(n846) );
  OAI22D0 U298 ( .A1(n839), .A2(n440), .B1(n825), .B2(n665), .ZN(n657) );
  OAI31D0 U299 ( .A1(n756), .A2(n785), .A3(n758), .B(n622), .ZN(n629) );
  CKND2D0 U300 ( .A1(n448), .A2(n430), .ZN(n593) );
  OAI211D0 U301 ( .A1(n449), .A2(n791), .B(n635), .C(n758), .ZN(n544) );
  CKND2D0 U302 ( .A1(n446), .A2(n747), .ZN(n745) );
  CKND2D1 U303 ( .A1(n782), .A2(n736), .ZN(n580) );
  AOI21D0 U304 ( .A1(n828), .A2(n863), .B(n703), .ZN(n510) );
  NR2D0 U305 ( .A1(n815), .A2(n447), .ZN(n626) );
  CKND2D0 U306 ( .A1(n449), .A2(a[6]), .ZN(n785) );
  AOI32D0 U307 ( .A1(n448), .A2(n844), .A3(n821), .B1(n822), .B2(n555), .ZN(
        n557) );
  OAI22D0 U308 ( .A1(a[6]), .A2(n448), .B1(n449), .B2(n766), .ZN(n555) );
  BUFFD4 U309 ( .I(a[3]), .Z(n447) );
  INVD1 U310 ( .I(n792), .ZN(n852) );
  INVD1 U311 ( .I(n684), .ZN(n866) );
  INVD1 U312 ( .I(n783), .ZN(n865) );
  INVD1 U313 ( .I(n607), .ZN(n831) );
  INVD1 U314 ( .I(n793), .ZN(n868) );
  INVD1 U315 ( .I(n574), .ZN(n860) );
  ND2D1 U316 ( .A1(n850), .A2(n837), .ZN(n792) );
  INVD1 U317 ( .I(n645), .ZN(n859) );
  ND2D1 U318 ( .A1(n803), .A2(n830), .ZN(n607) );
  INVD1 U319 ( .I(n714), .ZN(n814) );
  INVD1 U320 ( .I(n598), .ZN(n862) );
  INVD1 U321 ( .I(n778), .ZN(n833) );
  INVD1 U322 ( .I(n640), .ZN(n855) );
  ND2D1 U323 ( .A1(n826), .A2(n841), .ZN(n710) );
  INVD1 U324 ( .I(n644), .ZN(n861) );
  INVD1 U325 ( .I(n606), .ZN(n856) );
  INVD1 U326 ( .I(n731), .ZN(n848) );
  INVD1 U327 ( .I(n561), .ZN(n826) );
  INVD1 U328 ( .I(n615), .ZN(n854) );
  AOI221D0 U329 ( .A1(n810), .A2(n838), .B1(n833), .B2(n563), .C(n709), .ZN(
        n570) );
  OAI222D0 U330 ( .A1(n733), .A2(n606), .B1(n740), .B2(n685), .C1(n645), .C2(
        n769), .ZN(n554) );
  OAI221D0 U331 ( .A1(n624), .A2(n774), .B1(n759), .B2(n769), .C(n502), .ZN(
        n505) );
  AOI221D0 U332 ( .A1(n841), .A2(n439), .B1(n828), .B2(n580), .C(n856), .ZN(
        n503) );
  OAI222D0 U333 ( .A1(n733), .A2(n758), .B1(n698), .B2(n694), .C1(n764), .C2(
        n562), .ZN(n540) );
  OAI222D0 U334 ( .A1(n736), .A2(n607), .B1(n733), .B2(n771), .C1(n623), .C2(
        n606), .ZN(n608) );
  OAI221D0 U335 ( .A1(n469), .A2(n784), .B1(n729), .B2(n781), .C(n574), .ZN(
        n476) );
  OAI222D0 U336 ( .A1(n769), .A2(n777), .B1(n791), .B2(n655), .C1(n758), .C2(
        n714), .ZN(n663) );
  INVD1 U337 ( .I(n758), .ZN(n828) );
  OAI222D0 U338 ( .A1(n734), .A2(n733), .B1(n732), .B2(n731), .C1(n730), .C2(
        n729), .ZN(n801) );
  NR4D0 U339 ( .A1(n751), .A2(n750), .A3(n749), .A4(n748), .ZN(n800) );
  ND2D1 U340 ( .A1(n847), .A2(n833), .ZN(n729) );
  NR2D1 U341 ( .A1(n629), .A2(n628), .ZN(n630) );
  NR4D0 U342 ( .A1(n668), .A2(n667), .A3(n666), .A4(n750), .ZN(n669) );
  NR4D0 U343 ( .A1(n484), .A2(n483), .A3(n720), .A4(n482), .ZN(n485) );
  AOI221D0 U344 ( .A1(n817), .A2(n849), .B1(n857), .B2(n823), .C(n554), .ZN(
        n590) );
  NR4D0 U345 ( .A1(n586), .A2(n585), .A3(n584), .A4(n748), .ZN(n587) );
  ND2D1 U346 ( .A1(n853), .A2(n837), .ZN(n645) );
  AOI211D1 U347 ( .A1(n867), .A2(n526), .B(n525), .C(n524), .ZN(n553) );
  INR4D0 U348 ( .A1(n768), .B1(n530), .B2(n749), .B3(n719), .ZN(n552) );
  OAI221D0 U349 ( .A1(n433), .A2(n678), .B1(n730), .B2(n684), .C(n533), .ZN(
        n550) );
  INVD1 U350 ( .I(n784), .ZN(n821) );
  NR3D0 U351 ( .A1(n517), .A2(n759), .A3(n794), .ZN(n483) );
  CKND1 U352 ( .I(n443), .ZN(n444) );
  ND2D1 U353 ( .A1(n498), .A2(n497), .ZN(n499) );
  NR2D1 U354 ( .A1(n634), .A2(n752), .ZN(n776) );
  INVD1 U355 ( .I(n752), .ZN(n805) );
  INVD1 U356 ( .I(n736), .ZN(n863) );
  INVD1 U357 ( .I(n756), .ZN(n813) );
  INVD1 U358 ( .I(n777), .ZN(n838) );
  INVD1 U359 ( .I(n737), .ZN(n812) );
  NR2D1 U360 ( .A1(n715), .A2(n718), .ZN(n726) );
  ND2D1 U361 ( .A1(n690), .A2(n850), .ZN(n738) );
  INVD1 U362 ( .I(n712), .ZN(n830) );
  INVD1 U363 ( .I(n517), .ZN(n840) );
  OAI221D0 U364 ( .A1(n458), .A2(n620), .B1(n784), .B2(n727), .C(n457), .ZN(
        n468) );
  OAI221D0 U365 ( .A1(n747), .A2(n693), .B1(n755), .B2(n712), .C(n692), .ZN(
        n700) );
  OAI221D0 U366 ( .A1(n461), .A2(n432), .B1(n781), .B2(n740), .C(n460), .ZN(
        n467) );
  AOI222D0 U367 ( .A1(n813), .A2(n835), .B1(n40), .B2(n491), .C1(n808), .C2(
        n838), .ZN(n496) );
  OAI222D0 U368 ( .A1(n450), .A2(n780), .B1(n779), .B2(n778), .C1(n789), .C2(
        n777), .ZN(n787) );
  NR4D0 U369 ( .A1(n464), .A2(n463), .A3(n538), .A4(n462), .ZN(n465) );
  OAI222D0 U370 ( .A1(n755), .A2(n562), .B1(n651), .B2(n727), .C1(n756), .C2(
        n694), .ZN(n464) );
  OAI222D0 U371 ( .A1(n446), .A2(n660), .B1(n659), .B2(n793), .C1(n658), .C2(
        n792), .ZN(n661) );
  OAI222D0 U372 ( .A1(n739), .A2(n728), .B1(n706), .B2(n451), .C1(n705), .C2(
        n782), .ZN(n707) );
  INVD1 U373 ( .I(n776), .ZN(n845) );
  OAI222D0 U374 ( .A1(n453), .A2(n785), .B1(n753), .B2(n766), .C1(n760), .C2(
        n756), .ZN(n494) );
  OAI222D0 U375 ( .A1(n627), .A2(n783), .B1(n626), .B2(n731), .C1(n625), .C2(
        n764), .ZN(n628) );
  OA22D0 U376 ( .A1(n785), .A2(n752), .B1(n736), .B2(n624), .Z(n625) );
  OAI222D0 U377 ( .A1(n583), .A2(n783), .B1(n792), .B2(n582), .C1(n581), .C2(
        n785), .ZN(n586) );
  OAI222D0 U378 ( .A1(n766), .A2(n635), .B1(n447), .B2(n634), .C1(n760), .C2(
        n777), .ZN(n638) );
  OAI222D0 U379 ( .A1(n645), .A2(n430), .B1(n619), .B2(n612), .C1(n447), .C2(
        n729), .ZN(n617) );
  NR4D0 U380 ( .A1(n778), .A2(n766), .A3(n429), .A4(n447), .ZN(n748) );
  OAI221D0 U381 ( .A1(n747), .A2(n736), .B1(n454), .B2(n792), .C(n735), .ZN(
        n742) );
  NR4D0 U382 ( .A1(n512), .A2(n511), .A3(n527), .A4(n528), .ZN(n513) );
  OAI222D0 U383 ( .A1(n772), .A2(n771), .B1(n770), .B2(n769), .C1(n433), .C2(
        n768), .ZN(n797) );
  OAI221D0 U384 ( .A1(n759), .A2(n761), .B1(n440), .B2(n794), .C(n643), .ZN(
        n654) );
  ND2D1 U385 ( .A1(n449), .A2(n819), .ZN(n777) );
  OAI221D0 U386 ( .A1(n619), .A2(n593), .B1(n447), .B2(n783), .C(n710), .ZN(
        n535) );
  NR3D0 U387 ( .A1(n747), .A2(n448), .A3(n619), .ZN(n656) );
  NR2D1 U388 ( .A1(n447), .A2(n449), .ZN(n690) );
  NR3D0 U389 ( .A1(n713), .A2(n832), .A3(n440), .ZN(n529) );
  NR3D0 U390 ( .A1(n747), .A2(n447), .A3(n774), .ZN(n539) );
  ND2D1 U391 ( .A1(n449), .A2(n450), .ZN(n711) );
  NR3D0 U392 ( .A1(n728), .A2(n448), .A3(n844), .ZN(n667) );
  ND2D1 U393 ( .A1(n448), .A2(n447), .ZN(n759) );
  INVD1 U394 ( .I(n782), .ZN(n842) );
  NR3D0 U395 ( .A1(n784), .A2(n450), .A3(n448), .ZN(n676) );
  AOI221D0 U396 ( .A1(n803), .A2(n820), .B1(n808), .B2(n834), .C(n603), .ZN(
        n604) );
  AOI222D0 U397 ( .A1(n809), .A2(n827), .B1(n829), .B2(n811), .C1(n812), .C2(
        n449), .ZN(n605) );
  INVD1 U398 ( .I(a[0]), .ZN(n802) );
  INVD1 U399 ( .I(n785), .ZN(n843) );
  OAI222D0 U400 ( .A1(n521), .A2(n752), .B1(n520), .B2(n759), .C1(n519), .C2(
        n772), .ZN(n525) );
  OAI222D0 U401 ( .A1(n510), .A2(n753), .B1(n825), .B2(n509), .C1(n508), .C2(
        n727), .ZN(n512) );
  ND2D1 U402 ( .A1(n450), .A2(n506), .ZN(n509) );
  INVD1 U403 ( .I(a[1]), .ZN(n456) );
  NR4D0 U404 ( .A1(a[6]), .A2(n819), .A3(n736), .A4(n769), .ZN(n511) );
  AO221D0 U405 ( .A1(n442), .A2(n838), .B1(n806), .B2(n821), .C(n709), .Z(n662) );
  AOI32D0 U406 ( .A1(n442), .A2(n451), .A3(n838), .B1(n806), .B2(n558), .ZN(
        n560) );
  INVD1 U407 ( .I(n718), .ZN(n439) );
  INVD1 U408 ( .I(n439), .ZN(n440) );
  ND2D1 U409 ( .A1(n448), .A2(n819), .ZN(n718) );
  OA222D0 U410 ( .A1(n756), .A2(n440), .B1(n758), .B2(n733), .C1(n694), .C2(
        n429), .Z(n559) );
  INVD1 U411 ( .I(n565), .ZN(n808) );
  OAI211D1 U412 ( .A1(n561), .A2(n727), .B(n560), .C(n559), .ZN(n572) );
  OAI221D0 U413 ( .A1(n451), .A2(n740), .B1(n713), .B2(n727), .C(n702), .ZN(
        n708) );
  NR3D0 U414 ( .A1(n727), .A2(n825), .A3(n738), .ZN(n584) );
  AOI21D1 U415 ( .A1(n803), .A2(n657), .B(n656), .ZN(n660) );
  NR2D1 U416 ( .A1(n813), .A2(n803), .ZN(n623) );
  NR2D1 U417 ( .A1(n635), .A2(n727), .ZN(n709) );
  AOI31D0 U418 ( .A1(n740), .A2(n739), .A3(n738), .B(n737), .ZN(n741) );
  NR2D0 U419 ( .A1(n739), .A2(n447), .ZN(n703) );
  NR4D0 U420 ( .A1(n440), .A2(n772), .A3(n766), .A4(n832), .ZN(n744) );
  NR4D0 U421 ( .A1(n454), .A2(n844), .A3(n772), .A4(n764), .ZN(n704) );
  INVD1 U422 ( .I(n772), .ZN(n811) );
  OAI222D0 U423 ( .A1(n761), .A2(n770), .B1(n698), .B2(n729), .C1(n697), .C2(
        n789), .ZN(n699) );
  OAI33D0 U424 ( .A1(n761), .A2(n760), .A3(n759), .B1(n782), .B2(n430), .B3(
        n758), .ZN(n762) );
  OAI222D0 U425 ( .A1(n761), .A2(n615), .B1(n614), .B2(n430), .C1(n613), .C2(
        n684), .ZN(n616) );
  OAI22D0 U426 ( .A1(n764), .A2(n761), .B1(n664), .B2(n747), .ZN(n526) );
  OAI222D0 U427 ( .A1(n761), .A2(n694), .B1(n490), .B2(n774), .C1(n433), .C2(
        n759), .ZN(n501) );
  CKND2D0 U428 ( .A1(n733), .A2(n761), .ZN(n532) );
  AOI22D0 U429 ( .A1(n841), .A2(n757), .B1(n843), .B2(n40), .ZN(n765) );
  AOI221D1 U430 ( .A1(n805), .A2(n691), .B1(n690), .B2(n40), .C(n689), .ZN(
        n692) );
  AOI221D0 U431 ( .A1(n40), .A2(n545), .B1(n850), .B2(n544), .C(n543), .ZN(
        n546) );
  AOI32D0 U432 ( .A1(n450), .A2(n825), .A3(n442), .B1(n40), .B2(n459), .ZN(
        n460) );
  AOI22D0 U433 ( .A1(n834), .A2(n40), .B1(n809), .B2(n836), .ZN(n457) );
  AOI21D0 U434 ( .A1(n862), .A2(n823), .B(n703), .ZN(n706) );
  AOI211XD0 U435 ( .A1(n810), .A2(n829), .B(n831), .C(n704), .ZN(n705) );
  OAI222D0 U436 ( .A1(n785), .A2(n794), .B1(n784), .B2(n783), .C1(n782), .C2(
        n781), .ZN(n786) );
  ND3D1 U437 ( .A1(n724), .A2(n723), .A3(n722), .ZN(n443) );
  NR4D0 U438 ( .A1(n721), .A2(n744), .A3(n720), .A4(n719), .ZN(n722) );
  NR4D0 U439 ( .A1(a[0]), .A2(n839), .A3(n778), .A4(n784), .ZN(n585) );
  NR2D1 U440 ( .A1(n451), .A2(n768), .ZN(n750) );
  NR2D1 U441 ( .A1(n768), .A2(a[0]), .ZN(n720) );
  OA21D0 U442 ( .A1(n693), .A2(n451), .B(n623), .Z(n627) );
  OAI22D0 U443 ( .A1(n447), .A2(n620), .B1(n451), .B2(n619), .ZN(n621) );
  AOI22D0 U444 ( .A1(n813), .A2(a[0]), .B1(n453), .B2(n822), .ZN(n490) );
  AN4D1 U445 ( .A1(n679), .A2(n823), .A3(a[0]), .A4(n850), .Z(n527) );
  AOI32D1 U446 ( .A1(n449), .A2(n451), .A3(n823), .B1(n833), .B2(n642), .ZN(
        n643) );
  AOI211D1 U447 ( .A1(n848), .A2(a[0]), .B(n647), .C(n858), .ZN(n652) );
  AOI22D0 U448 ( .A1(n451), .A2(n823), .B1(n819), .B2(n811), .ZN(n599) );
  OAI22D0 U449 ( .A1(n451), .A2(n729), .B1(n456), .B2(n740), .ZN(n534) );
  NR3D0 U450 ( .A1(n451), .A2(n448), .A3(n694), .ZN(n603) );
  AOI22D0 U451 ( .A1(n830), .A2(n804), .B1(n829), .B2(n446), .ZN(n581) );
  AOI31D0 U452 ( .A1(n446), .A2(n832), .A3(n805), .B(n831), .ZN(n502) );
  AOI21D0 U453 ( .A1(n739), .A2(n678), .B(n446), .ZN(n637) );
  OAI31D0 U454 ( .A1(n819), .A2(n810), .A3(n815), .B(n701), .ZN(n498) );
  NR3D0 U455 ( .A1(n680), .A2(n442), .A3(n821), .ZN(n658) );
  INVD1 U456 ( .I(n747), .ZN(n806) );
  INVD1 U457 ( .I(n764), .ZN(n827) );
  NR2XD0 U458 ( .A1(n838), .A2(n834), .ZN(n682) );
  NR3D0 U459 ( .A1(n832), .A2(n454), .A3(n733), .ZN(n538) );
  AOI21D0 U460 ( .A1(n694), .A2(n774), .B(n733), .ZN(n689) );
  OAI22D0 U461 ( .A1(n465), .A2(n789), .B1(n756), .B2(n644), .ZN(n466) );
  NR4D0 U462 ( .A1(n694), .A2(n761), .A3(n789), .A4(n825), .ZN(n666) );
  AOI21D0 U463 ( .A1(n784), .A2(n754), .B(n789), .ZN(n636) );
  AOI21D1 U464 ( .A1(n838), .A2(n847), .B(n856), .ZN(n674) );
endmodule


module aes_sbox_15 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n35, n70, n71, n120, n122, n192, n196, n277, n389, n390, n398, n399,
         n400, n404, n405, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852;

  AN2XD1 U28 ( .A1(n711), .A2(n710), .Z(n715) );
  OA21D1 U35 ( .A1(n695), .A2(n694), .B(n693), .Z(n700) );
  OR3D1 U88 ( .A1(n434), .A2(n801), .A3(n444), .Z(n625) );
  OR4D1 U199 ( .A1(n649), .A2(n568), .A3(n512), .A4(n511), .Z(n514) );
  AN2XD1 U215 ( .A1(n513), .A2(n799), .Z(n512) );
  AN2XD1 U271 ( .A1(n526), .A2(n723), .Z(n464) );
  ND4D2 U1 ( .A1(n500), .A2(n499), .A3(n498), .A4(n497), .ZN(d[6]) );
  AOI221D2 U2 ( .A1(n849), .A2(n440), .B1(n841), .B2(n797), .C(n624), .ZN(n655) );
  IIND4D4 U3 ( .A1(n122), .A2(n192), .B1(n472), .B2(n471), .ZN(d[7]) );
  INVD1 U4 ( .I(n677), .ZN(n820) );
  INVD2 U5 ( .I(n739), .ZN(n812) );
  INVD2 U6 ( .I(n439), .ZN(n828) );
  ND2D1 U7 ( .A1(n437), .A2(n803), .ZN(n701) );
  INVD3 U8 ( .I(n436), .ZN(n803) );
  NR2D1 U9 ( .A1(n462), .A2(n739), .ZN(n425) );
  AOI221D2 U10 ( .A1(n790), .A2(n847), .B1(n799), .B2(n826), .C(n458), .ZN(
        n462) );
  AOI221D1 U11 ( .A1(n684), .A2(n431), .B1(n442), .B2(n843), .C(n548), .ZN(
        n553) );
  OAI22D2 U12 ( .A1(n714), .A2(n742), .B1(n441), .B2(n721), .ZN(n656) );
  ND2D2 U13 ( .A1(n673), .A2(n834), .ZN(n721) );
  CKND2D2 U14 ( .A1(n435), .A2(n443), .ZN(n735) );
  CKND2 U15 ( .I(a[1]), .ZN(n443) );
  OAI222D1 U16 ( .A1(n742), .A2(n598), .B1(n597), .B2(n441), .C1(n596), .C2(
        n667), .ZN(n599) );
  ND2D2 U17 ( .A1(n841), .A2(n440), .ZN(n629) );
  OAI221D1 U18 ( .A1(n730), .A2(n723), .B1(n696), .B2(n431), .C(n585), .ZN(
        n593) );
  CKND3 U19 ( .I(n70), .ZN(n431) );
  INVD4 U20 ( .I(n437), .ZN(n809) );
  BUFFD4 U21 ( .I(n788), .Z(n441) );
  BUFFD6 U22 ( .I(a[0]), .Z(n435) );
  ND2D1 U23 ( .A1(n817), .A2(n823), .ZN(n648) );
  ND2D1 U24 ( .A1(n436), .A2(a[2]), .ZN(n634) );
  ND2D0 U25 ( .A1(n440), .A2(n441), .ZN(n753) );
  CKND2D2 U26 ( .A1(n442), .A2(n440), .ZN(n730) );
  INVD3 U27 ( .I(n443), .ZN(n442) );
  CKND2D1 U29 ( .A1(n803), .A2(n809), .ZN(n745) );
  INVD2 U30 ( .I(n696), .ZN(n837) );
  INVD2 U31 ( .I(n716), .ZN(n789) );
  AO21D1 U32 ( .A1(n786), .A2(n824), .B(n726), .Z(n458) );
  INVD1 U33 ( .I(n735), .ZN(n786) );
  CKND2D1 U34 ( .A1(n436), .A2(n438), .ZN(n677) );
  CKND2D1 U36 ( .A1(n436), .A2(n809), .ZN(n739) );
  BUFFD6 U37 ( .I(a[7]), .Z(n439) );
  NR2D1 U38 ( .A1(n694), .A2(n431), .ZN(n726) );
  OA221D0 U39 ( .A1(n390), .A2(n442), .B1(n745), .B2(n398), .C(n399), .Z(n472)
         );
  NR3D0 U40 ( .A1(n405), .A2(n424), .A3(n488), .ZN(n498) );
  OAI31D2 U41 ( .A1(n808), .A2(n434), .A3(n789), .B(n663), .ZN(n664) );
  ND2D1 U42 ( .A1(n436), .A2(n444), .ZN(n668) );
  AOI221D1 U43 ( .A1(n790), .A2(n814), .B1(n798), .B2(n820), .C(n756), .ZN(
        n771) );
  AN2XD1 U44 ( .A1(n435), .A2(n803), .Z(n434) );
  INVD1 U45 ( .I(n745), .ZN(n811) );
  INVD1 U46 ( .I(n668), .ZN(n808) );
  OAI32D1 U47 ( .A1(n577), .A2(n431), .A3(n677), .B1(n576), .B2(n755), .ZN(
        n578) );
  AOI21D1 U48 ( .A1(n804), .A2(n442), .B(n793), .ZN(n576) );
  INVD1 U49 ( .I(n648), .ZN(n825) );
  INVD1 U50 ( .I(n750), .ZN(n799) );
  ND2D1 U51 ( .A1(n435), .A2(a[2]), .ZN(n750) );
  INVD1 U52 ( .I(a[1]), .ZN(n444) );
  ND2D1 U53 ( .A1(n809), .A2(n817), .ZN(n759) );
  INVD2 U54 ( .I(n657), .ZN(n795) );
  ND2D2 U55 ( .A1(a[1]), .A2(n441), .ZN(n775) );
  ND2D2 U56 ( .A1(n439), .A2(n823), .ZN(n747) );
  ND2D1 U57 ( .A1(n837), .A2(n821), .ZN(n628) );
  INVD1 U58 ( .I(n676), .ZN(n804) );
  NR3D0 U59 ( .A1(n428), .A2(n429), .A3(n726), .ZN(n585) );
  NR4D0 U60 ( .A1(n452), .A2(n451), .A3(n522), .A4(n450), .ZN(n453) );
  INVD1 U61 ( .I(n442), .ZN(n71) );
  NR3D1 U62 ( .A1(n425), .A2(n426), .A3(n427), .ZN(n389) );
  NR4D0 U63 ( .A1(n524), .A2(n523), .A3(n522), .A4(n586), .ZN(n525) );
  MAOI22D1 U64 ( .A1(n846), .A2(n803), .B1(n618), .B2(n763), .ZN(n505) );
  ND4D3 U65 ( .A1(n654), .A2(n655), .A3(n653), .A4(n652), .ZN(d[2]) );
  NR2D1 U66 ( .A1(n612), .A2(n611), .ZN(n613) );
  CKND2 U67 ( .I(n656), .ZN(n835) );
  INR4D2 U68 ( .A1(n662), .B1(n661), .B2(n660), .B3(n844), .ZN(n670) );
  ND2D1 U69 ( .A1(a[1]), .A2(n435), .ZN(n710) );
  AN2XD1 U70 ( .A1(n436), .A2(n817), .Z(n35) );
  AN2XD1 U71 ( .A1(n440), .A2(n443), .Z(n70) );
  AOI211XD0 U72 ( .A1(n852), .A2(n798), .B(n473), .C(n656), .ZN(n500) );
  OAI222D0 U73 ( .A1(n634), .A2(n714), .B1(n583), .B2(n723), .C1(n628), .C2(
        n657), .ZN(n473) );
  OA221D0 U74 ( .A1(n457), .A2(n765), .B1(n712), .B2(n762), .C(n558), .Z(n120)
         );
  AO221D1 U75 ( .A1(n834), .A2(n456), .B1(n455), .B2(n440), .C(n454), .Z(n122)
         );
  OAI221D1 U76 ( .A1(n71), .A2(n120), .B1(n590), .B2(n648), .C(n389), .ZN(n192) );
  AOI221D2 U77 ( .A1(n848), .A2(n637), .B1(n845), .B2(n792), .C(n636), .ZN(
        n654) );
  OAI221D1 U78 ( .A1(n740), .A2(n742), .B1(n701), .B2(n775), .C(n626), .ZN(
        n637) );
  AN2XD1 U79 ( .A1(n831), .A2(n489), .Z(n405) );
  AOI211XD0 U80 ( .A1(n793), .A2(n813), .B(n816), .C(n687), .ZN(n688) );
  AOI221D1 U81 ( .A1(n795), .A2(n529), .B1(n834), .B2(n528), .C(n527), .ZN(
        n530) );
  AOI221D1 U82 ( .A1(n787), .A2(n679), .B1(n822), .B2(n789), .C(n678), .ZN(
        n680) );
  CKBD4 U83 ( .I(a[6]), .Z(n196) );
  OA221D1 U84 ( .A1(n432), .A2(n730), .B1(n745), .B2(n657), .C(n433), .Z(n669)
         );
  OA221D1 U85 ( .A1(n549), .A2(n623), .B1(n710), .B2(n774), .C(n277), .Z(n616)
         );
  OA222D1 U86 ( .A1(n634), .A2(n627), .B1(n583), .B2(n582), .C1(n747), .C2(
        n581), .Z(n277) );
  AOI221D1 U87 ( .A1(n850), .A2(n443), .B1(n832), .B2(n710), .C(n518), .ZN(
        n521) );
  AOI211XD0 U89 ( .A1(n848), .A2(n485), .B(n484), .C(n483), .ZN(n499) );
  OAI22D0 U90 ( .A1(n444), .A2(n623), .B1(n622), .B2(n735), .ZN(n624) );
  OAI222D1 U91 ( .A1(n657), .A2(n758), .B1(n435), .B2(n550), .C1(n740), .C2(
        n549), .ZN(n551) );
  ND2D1 U92 ( .A1(n790), .A2(n435), .ZN(n549) );
  OA21D0 U93 ( .A1(n634), .A2(n722), .B(n774), .Z(n390) );
  OA222D0 U94 ( .A1(n467), .A2(n698), .B1(n463), .B2(n696), .C1(n719), .C2(
        n720), .Z(n398) );
  OA22D0 U95 ( .A1(n465), .A2(n701), .B1(n464), .B2(n750), .Z(n399) );
  ND2D1 U96 ( .A1(n35), .A2(n837), .ZN(n589) );
  OAI221D2 U97 ( .A1(n659), .A2(n668), .B1(n658), .B2(n657), .C(n835), .ZN(
        n661) );
  ND4D2 U98 ( .A1(n616), .A2(n615), .A3(n614), .A4(n613), .ZN(d[3]) );
  AOI221D1 U99 ( .A1(n805), .A2(n593), .B1(n831), .B2(n592), .C(n591), .ZN(
        n615) );
  OAI222D1 U100 ( .A1(n716), .A2(n739), .B1(n681), .B2(n677), .C1(n745), .C2(
        n546), .ZN(n524) );
  ND2D2 U101 ( .A1(n435), .A2(n441), .ZN(n716) );
  AOI211XD1 U102 ( .A1(n35), .A2(n580), .B(n578), .C(n579), .ZN(n581) );
  AOI211XD0 U103 ( .A1(n832), .A2(n435), .B(n630), .C(n842), .ZN(n635) );
  OAI222D1 U104 ( .A1(n716), .A2(n526), .B1(n480), .B2(n741), .C1(n479), .C2(
        n745), .ZN(n484) );
  INVD1 U105 ( .I(n629), .ZN(n842) );
  CKND2D1 U106 ( .A1(n801), .A2(n442), .ZN(n575) );
  AOI221D1 U107 ( .A1(n692), .A2(n847), .B1(n806), .B2(n691), .C(n690), .ZN(
        n706) );
  OAI222D1 U108 ( .A1(n635), .A2(n634), .B1(n750), .B2(n752), .C1(n633), .C2(
        n762), .ZN(n636) );
  ND2D2 U109 ( .A1(n439), .A2(n196), .ZN(n696) );
  AOI211XD0 U110 ( .A1(n808), .A2(n435), .B(n806), .C(n799), .ZN(n596) );
  AOI222D1 U111 ( .A1(n797), .A2(n819), .B1(n795), .B2(n475), .C1(n791), .C2(
        n822), .ZN(n480) );
  OAI21D0 U112 ( .A1(n648), .A2(n739), .B(n721), .ZN(n529) );
  NR3D1 U113 ( .A1(n555), .A2(n404), .A3(n400), .ZN(n573) );
  OAI222D1 U114 ( .A1(n554), .A2(n747), .B1(n553), .B2(n676), .C1(n552), .C2(
        n741), .ZN(n555) );
  CKND2D1 U115 ( .A1(n439), .A2(n817), .ZN(n719) );
  INVD2 U116 ( .I(n763), .ZN(n826) );
  ND2D2 U117 ( .A1(n196), .A2(n817), .ZN(n763) );
  INVD3 U118 ( .I(n770), .ZN(n831) );
  ND2D1 U119 ( .A1(n196), .A2(n828), .ZN(n770) );
  AOI21D0 U120 ( .A1(n765), .A2(n736), .B(n770), .ZN(n619) );
  OAI222D1 U121 ( .A1(n771), .A2(n770), .B1(n436), .B2(n829), .C1(n769), .C2(
        n440), .ZN(n777) );
  ND2D2 U122 ( .A1(n819), .A2(n831), .ZN(n714) );
  OAI222D1 U123 ( .A1(n736), .A2(n710), .B1(n759), .B2(n575), .C1(n740), .C2(
        n750), .ZN(n579) );
  ND2D1 U124 ( .A1(n831), .A2(n818), .ZN(n712) );
  AOI221D1 U125 ( .A1(n460), .A2(n797), .B1(n841), .B2(n807), .C(n459), .ZN(
        n461) );
  AO31D1 U126 ( .A1(n792), .A2(n848), .A3(n673), .B(n709), .Z(n459) );
  OAI222D1 U127 ( .A1(n521), .A2(n765), .B1(n716), .B2(n617), .C1(n520), .C2(
        n710), .ZN(n533) );
  NR4D1 U128 ( .A1(n777), .A2(n778), .A3(n779), .A4(n776), .ZN(n780) );
  OA21D0 U129 ( .A1(n676), .A2(n440), .B(n606), .Z(n610) );
  OAI22D1 U130 ( .A1(n755), .A2(n765), .B1(n442), .B2(n754), .ZN(n756) );
  OA221D1 U131 ( .A1(n676), .A2(n666), .B1(n665), .B2(n775), .C(n664), .Z(n433) );
  AOI221D1 U132 ( .A1(n836), .A2(n440), .B1(n846), .B2(n442), .C(n632), .ZN(
        n633) );
  OAI22D0 U133 ( .A1(n431), .A2(n698), .B1(n631), .B2(n730), .ZN(n632) );
  ND2D3 U134 ( .A1(n823), .A2(n828), .ZN(n741) );
  BUFFD8 U135 ( .I(a[3]), .Z(n436) );
  NR2D1 U136 ( .A1(n789), .A2(n786), .ZN(n681) );
  NR2D1 U137 ( .A1(n617), .A2(n735), .ZN(n757) );
  CKAN2D1 U138 ( .A1(n435), .A2(n557), .Z(n400) );
  CKAN2D1 U139 ( .A1(n831), .A2(n556), .Z(n404) );
  OAI211D0 U140 ( .A1(n545), .A2(n710), .B(n544), .C(n543), .ZN(n556) );
  AOI221D1 U141 ( .A1(n845), .A2(n430), .B1(n848), .B2(n683), .C(n682), .ZN(
        n707) );
  ND2D2 U142 ( .A1(n792), .A2(n440), .ZN(n546) );
  INVD4 U143 ( .I(n775), .ZN(n792) );
  ND2D2 U144 ( .A1(a[2]), .A2(n444), .ZN(n657) );
  INVD2 U145 ( .I(n742), .ZN(n790) );
  NR4D1 U146 ( .A1(n534), .A2(n533), .A3(n532), .A4(n531), .ZN(n535) );
  AOI221D1 U147 ( .A1(n812), .A2(n848), .B1(n801), .B2(n821), .C(n519), .ZN(
        n520) );
  INVD4 U148 ( .I(n196), .ZN(n823) );
  ND2D4 U149 ( .A1(n438), .A2(n809), .ZN(n755) );
  INVD2 U150 ( .I(n755), .ZN(n821) );
  AOI221D1 U151 ( .A1(n802), .A2(n564), .B1(n563), .B2(n812), .C(n562), .ZN(
        n572) );
  OAI22D0 U152 ( .A1(n453), .A2(n770), .B1(n737), .B2(n627), .ZN(n454) );
  CKAN2D1 U153 ( .A1(n791), .A2(n502), .Z(n424) );
  INVD1 U154 ( .I(n549), .ZN(n791) );
  NR2D0 U155 ( .A1(n677), .A2(n506), .ZN(n426) );
  NR2D0 U156 ( .A1(n461), .A2(n440), .ZN(n427) );
  CKND2D0 U157 ( .A1(n787), .A2(n848), .ZN(n506) );
  CKAN2D1 U158 ( .A1(n824), .A2(n430), .Z(n428) );
  AN2XD1 U159 ( .A1(n584), .A2(n443), .Z(n429) );
  AOI221D1 U160 ( .A1(n812), .A2(n785), .B1(n820), .B2(n797), .C(n551), .ZN(
        n552) );
  CKND2D1 U161 ( .A1(n441), .A2(n803), .ZN(n676) );
  OAI222D1 U162 ( .A1(n435), .A2(n670), .B1(n741), .B2(n669), .C1(n668), .C2(
        n667), .ZN(n671) );
  INVD1 U163 ( .I(n710), .ZN(n430) );
  ND2D1 U164 ( .A1(n797), .A2(n440), .ZN(n697) );
  BUFFD8 U165 ( .I(n784), .Z(n440) );
  AOI221D1 U166 ( .A1(n839), .A2(n799), .B1(n684), .B2(n792), .C(n671), .ZN(
        n708) );
  INVD2 U167 ( .I(n759), .ZN(n818) );
  NR2D1 U168 ( .A1(n741), .A2(n759), .ZN(n684) );
  OAI33D0 U169 ( .A1(n634), .A2(n439), .A3(n759), .B1(n694), .B2(n441), .B3(
        n740), .ZN(n527) );
  ND2D0 U170 ( .A1(n436), .A2(n817), .ZN(n432) );
  INVD4 U171 ( .I(n438), .ZN(n817) );
  OAI31D0 U172 ( .A1(n696), .A2(n438), .A3(n442), .B(n629), .ZN(n548) );
  ND2D1 U173 ( .A1(n442), .A2(n436), .ZN(n772) );
  ND2D0 U174 ( .A1(n438), .A2(n828), .ZN(n698) );
  CKND2D0 U175 ( .A1(n824), .A2(n814), .ZN(n526) );
  CKND2D0 U176 ( .A1(n811), .A2(n834), .ZN(n662) );
  ND2D0 U177 ( .A1(n442), .A2(n196), .ZN(n476) );
  INVD1 U178 ( .I(n773), .ZN(n836) );
  CKND0 U179 ( .I(n575), .ZN(n802) );
  CKND2D0 U180 ( .A1(n819), .A2(n848), .ZN(n667) );
  CKND2D0 U181 ( .A1(n817), .A2(n828), .ZN(n602) );
  NR2D0 U182 ( .A1(n797), .A2(n430), .ZN(n606) );
  CKND2D0 U183 ( .A1(n819), .A2(n443), .ZN(n666) );
  ND2D1 U184 ( .A1(n439), .A2(n490), .ZN(n493) );
  INVD0 U185 ( .I(n765), .ZN(n805) );
  ND2D0 U186 ( .A1(n435), .A2(n795), .ZN(n720) );
  ND2D0 U187 ( .A1(n438), .A2(n823), .ZN(n501) );
  ND2D0 U188 ( .A1(n441), .A2(n809), .ZN(n545) );
  CKND2D0 U189 ( .A1(n763), .A2(n719), .ZN(n564) );
  ND2D0 U190 ( .A1(n438), .A2(n196), .ZN(n766) );
  OAI31D0 U191 ( .A1(n790), .A2(n786), .A3(n801), .B(n849), .ZN(n481) );
  CKND0 U192 ( .I(n431), .ZN(n785) );
  AOI22D0 U193 ( .A1(n850), .A2(n792), .B1(n807), .B2(n836), .ZN(n540) );
  CKND2D0 U194 ( .A1(n851), .A2(n814), .ZN(n774) );
  NR2D0 U195 ( .A1(n794), .A2(n790), .ZN(n467) );
  CKND2D0 U196 ( .A1(n801), .A2(n843), .ZN(n558) );
  ND2D0 U197 ( .A1(n812), .A2(n851), .ZN(n751) );
  CKND0 U198 ( .I(n764), .ZN(n849) );
  NR2D0 U200 ( .A1(n709), .A2(n846), .ZN(n717) );
  AOI22D0 U201 ( .A1(n798), .A2(n847), .B1(n790), .B2(n826), .ZN(n561) );
  AOI22D0 U202 ( .A1(n841), .A2(n516), .B1(n684), .B2(n515), .ZN(n517) );
  CKND2D0 U203 ( .A1(n716), .A2(n742), .ZN(n516) );
  CKND2D0 U204 ( .A1(n772), .A2(n676), .ZN(n515) );
  OAI32D0 U205 ( .A1(n549), .A2(n747), .A3(n432), .B1(n507), .B2(n506), .ZN(
        n508) );
  NR2D0 U206 ( .A1(n821), .A2(n801), .ZN(n507) );
  CKND2D1 U207 ( .A1(n482), .A2(n481), .ZN(n483) );
  OAI22D0 U208 ( .A1(n745), .A2(n742), .B1(n647), .B2(n730), .ZN(n510) );
  NR2D0 U209 ( .A1(n826), .A2(n837), .ZN(n631) );
  AOI22D0 U210 ( .A1(n440), .A2(n807), .B1(n803), .B2(n794), .ZN(n583) );
  OAI21D0 U211 ( .A1(n740), .A2(n602), .B(n627), .ZN(n502) );
  CKND0 U212 ( .I(n740), .ZN(n813) );
  OAI22D0 U213 ( .A1(n735), .A2(n745), .B1(n594), .B2(n431), .ZN(n601) );
  NR2D0 U214 ( .A1(n815), .A2(n819), .ZN(n594) );
  NR2D0 U216 ( .A1(n440), .A2(n749), .ZN(n733) );
  AOI21D0 U217 ( .A1(n603), .A2(n648), .B(n676), .ZN(n491) );
  AOI31D0 U218 ( .A1(n723), .A2(n722), .A3(n721), .B(n720), .ZN(n724) );
  NR2D0 U219 ( .A1(n806), .A2(n813), .ZN(n647) );
  CKND2D0 U220 ( .A1(n818), .A2(n837), .ZN(n627) );
  CKND2D0 U221 ( .A1(n805), .A2(n442), .ZN(n711) );
  CKND2D0 U222 ( .A1(n673), .A2(n837), .ZN(n623) );
  CKND2D0 U223 ( .A1(n785), .A2(n803), .ZN(n713) );
  CKND0 U224 ( .I(n694), .ZN(n851) );
  CKND2D0 U225 ( .A1(n821), .A2(n828), .ZN(n617) );
  CKND2D0 U226 ( .A1(n820), .A2(n837), .ZN(n752) );
  CKND2D0 U227 ( .A1(n812), .A2(n837), .ZN(n598) );
  CKND2D1 U228 ( .A1(n588), .A2(n587), .ZN(n592) );
  OAI21D0 U229 ( .A1(n435), .A2(n677), .B(n739), .ZN(n475) );
  NR2D0 U230 ( .A1(n799), .A2(n797), .ZN(n463) );
  NR2D0 U231 ( .A1(n799), .A2(n436), .ZN(n609) );
  AOI21D0 U232 ( .A1(n812), .A2(n847), .B(n686), .ZN(n494) );
  AOI31D0 U233 ( .A1(n437), .A2(n823), .A3(n801), .B(n686), .ZN(n466) );
  CKND2D0 U234 ( .A1(n806), .A2(n809), .ZN(n595) );
  NR2XD0 U235 ( .A1(n639), .A2(n757), .ZN(n597) );
  CKND2D0 U236 ( .A1(n677), .A2(n739), .ZN(n679) );
  AOI22D0 U237 ( .A1(n819), .A2(n806), .B1(n795), .B2(n817), .ZN(n550) );
  OAI22D0 U238 ( .A1(n440), .A2(n712), .B1(n444), .B2(n723), .ZN(n518) );
  OAI33D0 U239 ( .A1(n745), .A2(n441), .A3(n719), .B1(n648), .B2(n442), .B3(
        n647), .ZN(n651) );
  OAI211D0 U240 ( .A1(n817), .A2(n745), .B(n762), .C(n740), .ZN(n674) );
  AOI21D0 U241 ( .A1(n845), .A2(n442), .B(n684), .ZN(n685) );
  ND4D0 U242 ( .A1(n786), .A2(n825), .A3(n437), .A4(n439), .ZN(n718) );
  OAI21D0 U243 ( .A1(n741), .A2(n603), .B(n712), .ZN(n584) );
  NR2D0 U244 ( .A1(n801), .A2(n794), .ZN(n446) );
  NR2D0 U245 ( .A1(n850), .A2(n836), .ZN(n457) );
  CKND2D0 U246 ( .A1(n720), .A2(n730), .ZN(n580) );
  OAI22D0 U247 ( .A1(n439), .A2(n648), .B1(n740), .B2(n719), .ZN(n447) );
  NR2D0 U248 ( .A1(n846), .A2(n684), .ZN(n449) );
  AOI32D0 U249 ( .A1(n439), .A2(n809), .A3(n790), .B1(n795), .B2(n447), .ZN(
        n448) );
  NR2D0 U250 ( .A1(n437), .A2(n823), .ZN(n460) );
  AOI211D0 U251 ( .A1(n766), .A2(n648), .B(n577), .C(n735), .ZN(n468) );
  CKND2D0 U252 ( .A1(n753), .A2(n750), .ZN(n738) );
  OAI22D0 U253 ( .A1(n436), .A2(n603), .B1(n440), .B2(n602), .ZN(n604) );
  AOI33D0 U254 ( .A1(n604), .A2(n823), .A3(n792), .B1(n843), .B2(n803), .B3(
        n787), .ZN(n605) );
  AOI211XD0 U255 ( .A1(n830), .A2(n798), .B(n478), .C(n477), .ZN(n479) );
  CKND0 U256 ( .I(n602), .ZN(n830) );
  AOI32D0 U257 ( .A1(n790), .A2(n440), .A3(n822), .B1(n787), .B2(n542), .ZN(
        n544) );
  CKND2D0 U258 ( .A1(n740), .A2(n736), .ZN(n542) );
  NR2D0 U259 ( .A1(n722), .A2(n436), .ZN(n686) );
  OAI22D0 U260 ( .A1(n823), .A2(n701), .B1(n809), .B2(n648), .ZN(n640) );
  AOI22D0 U261 ( .A1(n801), .A2(n821), .B1(n804), .B2(n817), .ZN(n754) );
  AOI32D0 U262 ( .A1(n438), .A2(n440), .A3(n807), .B1(n818), .B2(n625), .ZN(
        n626) );
  NR2D0 U263 ( .A1(n749), .A2(n435), .ZN(n703) );
  OAI22D0 U264 ( .A1(n755), .A2(n676), .B1(n681), .B2(n701), .ZN(n451) );
  AOI21D0 U265 ( .A1(n676), .A2(n577), .B(n735), .ZN(n450) );
  AOI22D0 U266 ( .A1(n797), .A2(n435), .B1(n442), .B2(n806), .ZN(n474) );
  OAI31D0 U267 ( .A1(n730), .A2(n813), .A3(n741), .B(n729), .ZN(n734) );
  OAI21D0 U268 ( .A1(n700), .A2(n730), .B(n699), .ZN(n704) );
  AOI21D0 U269 ( .A1(n436), .A2(n848), .B(n808), .ZN(n760) );
  AOI21D0 U270 ( .A1(n836), .A2(n806), .B(n743), .ZN(n744) );
  OAI33D0 U272 ( .A1(n742), .A2(n741), .A3(n740), .B1(n763), .B2(n441), .B3(
        n739), .ZN(n743) );
  AOI21D0 U273 ( .A1(n796), .A2(n834), .B(n563), .ZN(n504) );
  CKND2D0 U274 ( .A1(n710), .A2(n803), .ZN(n566) );
  AOI32D0 U275 ( .A1(n437), .A2(n828), .A3(n805), .B1(n806), .B2(n539), .ZN(
        n541) );
  OAI22D0 U276 ( .A1(n196), .A2(n437), .B1(n438), .B2(n747), .ZN(n539) );
  INVD1 U277 ( .I(a[2]), .ZN(n788) );
  BUFFD4 U278 ( .I(a[4]), .Z(n437) );
  BUFFD4 U279 ( .I(a[5]), .Z(n438) );
  INVD1 U280 ( .I(n667), .ZN(n850) );
  INVD1 U281 ( .I(n558), .ZN(n844) );
  INVD1 U282 ( .I(n774), .ZN(n852) );
  INVD1 U283 ( .I(n582), .ZN(n846) );
  INVD1 U284 ( .I(n627), .ZN(n845) );
  INVD1 U285 ( .I(n697), .ZN(n798) );
  INVD1 U286 ( .I(n628), .ZN(n843) );
  INVD1 U287 ( .I(n714), .ZN(n832) );
  INVD1 U288 ( .I(n623), .ZN(n839) );
  INVD1 U289 ( .I(n712), .ZN(n833) );
  INVD1 U290 ( .I(n590), .ZN(n816) );
  ND2D1 U291 ( .A1(n810), .A2(n825), .ZN(n693) );
  INVD1 U292 ( .I(n722), .ZN(n841) );
  INVD1 U293 ( .I(n589), .ZN(n840) );
  INVD1 U294 ( .I(n598), .ZN(n838) );
  OAI222D0 U295 ( .A1(n561), .A2(n701), .B1(n560), .B2(n735), .C1(n442), .C2(
        n559), .ZN(n562) );
  AOI21D1 U296 ( .A1(n810), .A2(n851), .B(n838), .ZN(n560) );
  AOI21D1 U297 ( .A1(n850), .A2(n806), .B(n844), .ZN(n559) );
  IND4D1 U298 ( .A1(n783), .B1(n782), .B2(n781), .B3(n780), .ZN(d[0]) );
  OAI222D0 U299 ( .A1(n717), .A2(n716), .B1(n715), .B2(n714), .C1(n713), .C2(
        n712), .ZN(n783) );
  NR4D0 U300 ( .A1(n734), .A2(n733), .A3(n732), .A4(n731), .ZN(n781) );
  NR4D0 U301 ( .A1(n701), .A2(n753), .A3(n747), .A4(n817), .ZN(n727) );
  AOI221D0 U302 ( .A1(n834), .A2(n601), .B1(n600), .B2(n440), .C(n599), .ZN(
        n614) );
  ND3D1 U303 ( .A1(n537), .A2(n536), .A3(n535), .ZN(d[5]) );
  AOI211D1 U304 ( .A1(n851), .A2(n510), .B(n509), .C(n508), .ZN(n537) );
  INR4D0 U305 ( .A1(n749), .B1(n514), .B2(n732), .B3(n702), .ZN(n536) );
  INVD1 U306 ( .I(n772), .ZN(n807) );
  OAI221D0 U307 ( .A1(n442), .A2(n662), .B1(n713), .B2(n667), .C(n517), .ZN(
        n534) );
  OAI222D0 U308 ( .A1(n742), .A2(n677), .B1(n474), .B2(n755), .C1(n442), .C2(
        n740), .ZN(n485) );
  NR4D0 U309 ( .A1(n470), .A2(n469), .A3(n703), .A4(n468), .ZN(n471) );
  ND4D1 U310 ( .A1(n708), .A2(n707), .A3(n706), .A4(n705), .ZN(d[1]) );
  NR4D0 U311 ( .A1(n704), .A2(n727), .A3(n703), .A4(n702), .ZN(n705) );
  ND2D1 U312 ( .A1(n663), .A2(n848), .ZN(n764) );
  NR3D0 U313 ( .A1(n710), .A2(n809), .A3(n721), .ZN(n568) );
  INVD1 U314 ( .I(n701), .ZN(n814) );
  INVD1 U315 ( .I(n719), .ZN(n847) );
  NR2D1 U316 ( .A1(n698), .A2(n701), .ZN(n709) );
  INVD1 U317 ( .I(n762), .ZN(n801) );
  INVD1 U318 ( .I(n753), .ZN(n794) );
  INVD1 U319 ( .I(n747), .ZN(n848) );
  INVD1 U320 ( .I(n603), .ZN(n819) );
  ND2D1 U321 ( .A1(n430), .A2(n815), .ZN(n590) );
  AO221D0 U322 ( .A1(n790), .A2(n822), .B1(n787), .B2(n805), .C(n692), .Z(n645) );
  INVD1 U323 ( .I(n758), .ZN(n822) );
  ND2D1 U324 ( .A1(n819), .A2(n837), .ZN(n722) );
  INVD1 U325 ( .I(n720), .ZN(n796) );
  INVD1 U326 ( .I(n501), .ZN(n824) );
  INVD1 U327 ( .I(n741), .ZN(n834) );
  INVD1 U328 ( .I(n545), .ZN(n810) );
  AOI221D0 U329 ( .A1(n793), .A2(n822), .B1(n818), .B2(n547), .C(n692), .ZN(
        n554) );
  ND2D1 U330 ( .A1(n772), .A2(n546), .ZN(n547) );
  OAI222D0 U331 ( .A1(n719), .A2(n590), .B1(n716), .B2(n752), .C1(n606), .C2(
        n589), .ZN(n591) );
  OAI222D0 U332 ( .A1(n628), .A2(n441), .B1(n602), .B2(n595), .C1(n436), .C2(
        n712), .ZN(n600) );
  AOI221D0 U333 ( .A1(n825), .A2(n814), .B1(n812), .B2(n564), .C(n840), .ZN(
        n487) );
  OAI222D0 U334 ( .A1(n742), .A2(n751), .B1(n681), .B2(n712), .C1(n680), .C2(
        n770), .ZN(n682) );
  OAI221D0 U335 ( .A1(n730), .A2(n676), .B1(n432), .B2(n695), .C(n675), .ZN(
        n683) );
  AOI221D0 U336 ( .A1(n786), .A2(n674), .B1(n673), .B2(n795), .C(n672), .ZN(
        n675) );
  OAI222D0 U337 ( .A1(n722), .A2(n711), .B1(n689), .B2(n440), .C1(n688), .C2(
        n763), .ZN(n690) );
  AOI21D1 U338 ( .A1(n846), .A2(n807), .B(n686), .ZN(n689) );
  NR4D0 U339 ( .A1(n442), .A2(n828), .A3(n753), .A4(n745), .ZN(n687) );
  OAI222D0 U340 ( .A1(n800), .A2(n623), .B1(n546), .B2(n526), .C1(n525), .C2(
        n770), .ZN(n532) );
  NR3D0 U341 ( .A1(n730), .A2(n436), .A3(n755), .ZN(n523) );
  OAI222D0 U342 ( .A1(n697), .A2(n723), .B1(n435), .B2(n530), .C1(n775), .C2(
        n764), .ZN(n531) );
  OAI222D0 U343 ( .A1(n505), .A2(n735), .B1(n504), .B2(n740), .C1(n503), .C2(
        n753), .ZN(n509) );
  NR2D1 U344 ( .A1(n849), .A2(n502), .ZN(n503) );
  OAI222D0 U345 ( .A1(n610), .A2(n764), .B1(n609), .B2(n714), .C1(n608), .C2(
        n745), .ZN(n611) );
  OA22D0 U346 ( .A1(n766), .A2(n735), .B1(n719), .B2(n607), .Z(n608) );
  NR3D0 U347 ( .A1(n440), .A2(n437), .A3(n677), .ZN(n586) );
  NR2D1 U348 ( .A1(n436), .A2(n438), .ZN(n673) );
  OAI221D0 U349 ( .A1(n602), .A2(n577), .B1(n436), .B2(n764), .C(n693), .ZN(
        n519) );
  OAI222D0 U350 ( .A1(n748), .A2(n747), .B1(n746), .B2(n745), .C1(n435), .C2(
        n744), .ZN(n779) );
  OAI221D0 U351 ( .A1(n440), .A2(n723), .B1(n696), .B2(n710), .C(n685), .ZN(
        n691) );
  NR4D0 U352 ( .A1(n677), .A2(n742), .A3(n770), .A4(n809), .ZN(n649) );
  NR4D0 U353 ( .A1(n651), .A2(n650), .A3(n649), .A4(n733), .ZN(n652) );
  NR4D0 U354 ( .A1(n496), .A2(n495), .A3(n511), .A4(n512), .ZN(n497) );
  NR2XD0 U355 ( .A1(n832), .A2(n843), .ZN(n659) );
  INVD1 U356 ( .I(n757), .ZN(n829) );
  NR2XD0 U357 ( .A1(n768), .A2(n767), .ZN(n769) );
  NR3D0 U358 ( .A1(n730), .A2(n437), .A3(n602), .ZN(n639) );
  NR4D0 U359 ( .A1(n570), .A2(n569), .A3(n568), .A4(n731), .ZN(n571) );
  AOI221D0 U360 ( .A1(n801), .A2(n833), .B1(n841), .B2(n807), .C(n538), .ZN(
        n574) );
  ND2D1 U361 ( .A1(n436), .A2(n441), .ZN(n762) );
  OAI222D0 U362 ( .A1(n442), .A2(n766), .B1(n431), .B2(n747), .C1(n741), .C2(
        n737), .ZN(n478) );
  OAI221D0 U363 ( .A1(n730), .A2(n719), .B1(n442), .B2(n773), .C(n718), .ZN(
        n725) );
  OAI222D0 U364 ( .A1(n439), .A2(n761), .B1(n760), .B2(n759), .C1(n770), .C2(
        n758), .ZN(n768) );
  ND2D1 U365 ( .A1(n438), .A2(n803), .ZN(n758) );
  ND2D1 U366 ( .A1(n444), .A2(n441), .ZN(n742) );
  INVD1 U367 ( .I(n737), .ZN(n797) );
  NR3D0 U368 ( .A1(n696), .A2(n817), .A3(n701), .ZN(n513) );
  ND2D1 U369 ( .A1(n438), .A2(n439), .ZN(n694) );
  ND2D1 U370 ( .A1(n437), .A2(n441), .ZN(n577) );
  NR3D0 U371 ( .A1(n711), .A2(n437), .A3(n828), .ZN(n650) );
  AN2XD1 U372 ( .A1(n437), .A2(n438), .Z(n663) );
  ND2D1 U373 ( .A1(n437), .A2(n436), .ZN(n740) );
  INVD1 U374 ( .I(n435), .ZN(n784) );
  INVD1 U375 ( .I(n634), .ZN(n806) );
  AOI221D0 U376 ( .A1(n430), .A2(n804), .B1(n791), .B2(n35), .C(n586), .ZN(
        n587) );
  AOI222D0 U377 ( .A1(n792), .A2(n811), .B1(n813), .B2(n794), .C1(n796), .C2(
        n438), .ZN(n588) );
  OAI222D0 U378 ( .A1(n494), .A2(n431), .B1(n809), .B2(n493), .C1(n492), .C2(
        n710), .ZN(n496) );
  INR2D1 U379 ( .A1(n751), .B1(n491), .ZN(n492) );
  ND2D1 U380 ( .A1(n437), .A2(n817), .ZN(n603) );
  INVD1 U381 ( .I(n766), .ZN(n827) );
  AOI21D1 U382 ( .A1(n430), .A2(n640), .B(n639), .ZN(n643) );
  OAI221D0 U383 ( .A1(n607), .A2(n755), .B1(n740), .B2(n750), .C(n486), .ZN(
        n489) );
  NR4D0 U384 ( .A1(n621), .A2(n620), .A3(n838), .A4(n619), .ZN(n622) );
  AOI22D1 U385 ( .A1(n792), .A2(n825), .B1(n801), .B2(n809), .ZN(n761) );
  NR2D1 U386 ( .A1(n628), .A2(n713), .ZN(n732) );
  OAI22D0 U387 ( .A1(n444), .A2(n712), .B1(n442), .B2(n628), .ZN(n630) );
  INVD1 U388 ( .I(n730), .ZN(n787) );
  AOI22D0 U389 ( .A1(n825), .A2(n738), .B1(n827), .B2(n795), .ZN(n746) );
  AOI22D0 U390 ( .A1(n827), .A2(n795), .B1(n798), .B2(n826), .ZN(n465) );
  AOI22D0 U391 ( .A1(n35), .A2(n795), .B1(n792), .B2(n820), .ZN(n445) );
  NR2D1 U392 ( .A1(n785), .A2(n795), .ZN(n642) );
  NR2D1 U393 ( .A1(n789), .A2(n785), .ZN(n607) );
  AOI222D0 U394 ( .A1(n797), .A2(n814), .B1(n812), .B2(n789), .C1(n820), .C2(
        n795), .ZN(n543) );
  CKND2D0 U395 ( .A1(n789), .A2(n821), .ZN(n638) );
  OAI211D0 U396 ( .A1(n694), .A2(n668), .B(n541), .C(n540), .ZN(n557) );
  OAI222D0 U397 ( .A1(n716), .A2(n589), .B1(n723), .B2(n668), .C1(n628), .C2(
        n750), .ZN(n538) );
  NR3D0 U398 ( .A1(n501), .A2(n740), .A3(n775), .ZN(n469) );
  OAI22D0 U399 ( .A1(n775), .A2(n774), .B1(n773), .B2(n772), .ZN(n776) );
  OAI22D0 U400 ( .A1(n432), .A2(n742), .B1(n755), .B2(n775), .ZN(n678) );
  CKND2D1 U401 ( .A1(n834), .A2(n821), .ZN(n773) );
  ND2D1 U402 ( .A1(n442), .A2(a[2]), .ZN(n737) );
  ND2D0 U403 ( .A1(n437), .A2(a[2]), .ZN(n695) );
  CKND2D1 U404 ( .A1(a[2]), .A2(n809), .ZN(n618) );
  ND2D1 U405 ( .A1(a[2]), .A2(n803), .ZN(n765) );
  CKND2D0 U406 ( .A1(a[2]), .A2(n438), .ZN(n736) );
  OAI222D0 U407 ( .A1(a[2]), .A2(n643), .B1(n642), .B2(n774), .C1(n641), .C2(
        n773), .ZN(n644) );
  CKND2D0 U408 ( .A1(a[2]), .A2(n730), .ZN(n728) );
  OAI222D0 U409 ( .A1(n432), .A2(n546), .B1(n634), .B2(n710), .C1(n737), .C2(
        n677), .ZN(n452) );
  OA222D0 U410 ( .A1(n737), .A2(n432), .B1(n736), .B2(n431), .C1(n739), .C2(
        n735), .Z(n748) );
  OAI22D0 U411 ( .A1(n634), .A2(n735), .B1(n431), .B2(n762), .ZN(n490) );
  OAI221D0 U412 ( .A1(n449), .A2(n634), .B1(n762), .B2(n723), .C(n448), .ZN(
        n455) );
  OAI222D0 U413 ( .A1(n567), .A2(n764), .B1(n773), .B2(n566), .C1(n565), .C2(
        n766), .ZN(n570) );
  OAI31D1 U414 ( .A1(n737), .A2(n766), .A3(n739), .B(n605), .ZN(n612) );
  NR4D0 U415 ( .A1(n759), .A2(n747), .A3(n657), .A4(n436), .ZN(n731) );
  INR2D1 U416 ( .A1(n513), .B1(n657), .ZN(n702) );
  NR2D1 U417 ( .A1(n501), .A2(n657), .ZN(n563) );
  INVD1 U418 ( .I(n695), .ZN(n815) );
  NR2D0 U419 ( .A1(n618), .A2(n710), .ZN(n692) );
  OAI211D0 U420 ( .A1(n438), .A2(n772), .B(n618), .C(n739), .ZN(n528) );
  OAI222D0 U421 ( .A1(n753), .A2(n752), .B1(n751), .B2(n750), .C1(n442), .C2(
        n749), .ZN(n778) );
  NR4D0 U422 ( .A1(n196), .A2(n803), .A3(n719), .A4(n750), .ZN(n495) );
  OAI33D0 U423 ( .A1(n648), .A2(n435), .A3(n441), .B1(n476), .B2(n719), .B3(
        n750), .ZN(n477) );
  OAI222D0 U424 ( .A1(n766), .A2(n775), .B1(n765), .B2(n764), .C1(n763), .C2(
        n762), .ZN(n767) );
  NR3D0 U425 ( .A1(n765), .A2(n439), .A3(n437), .ZN(n660) );
  NR4D0 U426 ( .A1(n435), .A2(n823), .A3(n759), .A4(n765), .ZN(n569) );
  OAI222D0 U427 ( .A1(n773), .A2(n575), .B1(n765), .B2(n629), .C1(n487), .C2(
        n753), .ZN(n488) );
  OAI221D0 U428 ( .A1(n446), .A2(n603), .B1(n765), .B2(n710), .C(n445), .ZN(
        n456) );
  INVD1 U429 ( .I(n728), .ZN(n800) );
  AOI31D1 U430 ( .A1(n837), .A2(n728), .A3(n813), .B(n727), .ZN(n729) );
  AOI221D0 U431 ( .A1(n726), .A2(n805), .B1(n804), .B2(n725), .C(n724), .ZN(
        n782) );
  AN4D1 U432 ( .A1(n663), .A2(n807), .A3(n435), .A4(n834), .Z(n511) );
  ND3D0 U433 ( .A1(n806), .A2(n663), .A3(n834), .ZN(n749) );
  CKND2D0 U434 ( .A1(n663), .A2(n837), .ZN(n582) );
  ND2D1 U435 ( .A1(n831), .A2(n663), .ZN(n723) );
  OAI32D0 U436 ( .A1(n758), .A2(n467), .A3(n696), .B1(n466), .B2(n730), .ZN(
        n470) );
  OAI222D0 U437 ( .A1(n750), .A2(n758), .B1(n772), .B2(n638), .C1(n739), .C2(
        n697), .ZN(n646) );
  OA33D0 U438 ( .A1(n698), .A2(n740), .A3(n735), .B1(n697), .B2(n696), .B3(
        n758), .Z(n699) );
  OAI222D0 U439 ( .A1(n747), .A2(n618), .B1(n436), .B2(n617), .C1(n741), .C2(
        n758), .ZN(n621) );
  NR2D1 U440 ( .A1(n793), .A2(n796), .ZN(n567) );
  OAI31D0 U441 ( .A1(n803), .A2(n793), .A3(n799), .B(n684), .ZN(n482) );
  INVD1 U442 ( .I(n546), .ZN(n793) );
  NR3D0 U443 ( .A1(n434), .A2(n790), .A3(n805), .ZN(n641) );
  AOI22D0 U444 ( .A1(n815), .A2(n785), .B1(n813), .B2(a[2]), .ZN(n565) );
  AOI31D0 U445 ( .A1(a[2]), .A2(n817), .A3(n786), .B(n816), .ZN(n486) );
  AOI21D0 U446 ( .A1(n722), .A2(n662), .B(a[2]), .ZN(n620) );
  NR2XD0 U447 ( .A1(n822), .A2(n35), .ZN(n665) );
  ND4D1 U448 ( .A1(n574), .A2(n573), .A3(n572), .A4(n571), .ZN(d[4]) );
  NR3D0 U449 ( .A1(n817), .A2(n442), .A3(n716), .ZN(n522) );
  AOI21D0 U450 ( .A1(n677), .A2(n755), .B(n716), .ZN(n672) );
  AOI221D1 U451 ( .A1(n831), .A2(n646), .B1(n834), .B2(n645), .C(n644), .ZN(
        n653) );
  AOI21D1 U452 ( .A1(n822), .A2(n831), .B(n840), .ZN(n658) );
endmodule


module aes_sbox_14 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   N169, n70, n277, n342, n410, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864;

  OA21D1 U35 ( .A1(n703), .A2(n702), .B(n701), .Z(n708) );
  OR4D1 U199 ( .A1(n655), .A2(n574), .A3(n519), .A4(n518), .Z(n521) );
  MAOI22D1 U209 ( .A1(n858), .A2(n814), .B1(n624), .B2(n773), .ZN(n512) );
  AN2XD1 U215 ( .A1(n520), .A2(n810), .Z(n519) );
  AN2XD1 U271 ( .A1(n532), .A2(n731), .Z(n466) );
  ND2D2 U339 ( .A1(a[6]), .A2(n840), .ZN(n780) );
  AOI221D2 U1 ( .A1(n692), .A2(n430), .B1(a[1]), .B2(n855), .C(n554), .ZN(n559) );
  AOI221D1 U2 ( .A1(n846), .A2(n607), .B1(n606), .B2(n443), .C(n605), .ZN(n620) );
  AOI22D1 U3 ( .A1(n803), .A2(n837), .B1(n812), .B2(n820), .ZN(n771) );
  INVD2 U4 ( .I(a[1]), .ZN(n445) );
  NR2XD0 U5 ( .A1(n778), .A2(n777), .ZN(n779) );
  CKBD4 U6 ( .I(n794), .Z(n443) );
  ND2D0 U7 ( .A1(n441), .A2(n814), .ZN(n768) );
  AOI221D1 U8 ( .A1(n836), .A2(n795), .B1(n590), .B2(n444), .C(n734), .ZN(n591) );
  CKND2D1 U9 ( .A1(n814), .A2(n820), .ZN(n755) );
  NR2D2 U10 ( .A1(n800), .A2(n797), .ZN(n689) );
  NR4D1 U11 ( .A1(n530), .A2(n529), .A3(n528), .A4(n592), .ZN(n531) );
  OAI221D1 U12 ( .A1(n738), .A2(n684), .B1(n746), .B2(n703), .C(n683), .ZN(
        n691) );
  OAI22D1 U13 ( .A1(n430), .A2(n706), .B1(n637), .B2(n738), .ZN(n638) );
  OA221D1 U14 ( .A1(n749), .A2(n757), .B1(n772), .B2(n765), .C(n277), .Z(n526)
         );
  AOI221D1 U15 ( .A1(n470), .A2(n444), .B1(n822), .B2(n469), .C(n468), .ZN(
        n477) );
  OAI22D0 U16 ( .A1(n467), .A2(n709), .B1(n466), .B2(n760), .ZN(n468) );
  AOI221D1 U17 ( .A1(n813), .A2(n570), .B1(n569), .B2(n823), .C(n568), .ZN(
        n578) );
  AOI21D1 U18 ( .A1(n730), .A2(n668), .B(n438), .ZN(n626) );
  NR2D0 U19 ( .A1(n730), .A2(n439), .ZN(n694) );
  INVD2 U20 ( .I(n730), .ZN(n853) );
  ND2D3 U21 ( .A1(n831), .A2(n849), .ZN(n730) );
  INVD2 U22 ( .I(n785), .ZN(n803) );
  ND2D2 U23 ( .A1(a[1]), .A2(n799), .ZN(n785) );
  ND2D2 U24 ( .A1(n445), .A2(n799), .ZN(n752) );
  CKND2D0 U25 ( .A1(n799), .A2(n820), .ZN(n551) );
  INVD6 U26 ( .I(n438), .ZN(n799) );
  OAI222D1 U27 ( .A1(n724), .A2(n532), .B1(n487), .B2(n751), .C1(n486), .C2(
        n755), .ZN(n491) );
  CKND2D1 U28 ( .A1(n820), .A2(n828), .ZN(n769) );
  CKND2D1 U29 ( .A1(n439), .A2(n441), .ZN(n685) );
  INVD1 U30 ( .I(n747), .ZN(n808) );
  BUFFD6 U31 ( .I(a[2]), .Z(n438) );
  INVD1 U32 ( .I(a[6]), .ZN(n835) );
  ND2D0 U33 ( .A1(a[1]), .A2(n438), .ZN(n747) );
  INVD1 U34 ( .I(a[1]), .ZN(n444) );
  BUFFD6 U36 ( .I(a[3]), .Z(n439) );
  CKND2D1 U37 ( .A1(n828), .A2(n835), .ZN(n654) );
  INVD2 U38 ( .I(n663), .ZN(n806) );
  CKND2D1 U39 ( .A1(n439), .A2(n820), .ZN(n749) );
  ND2D1 U40 ( .A1(n437), .A2(n444), .ZN(n743) );
  ND2D2 U41 ( .A1(a[1]), .A2(n443), .ZN(n738) );
  INVD2 U42 ( .I(n772), .ZN(n812) );
  ND2D1 U43 ( .A1(n437), .A2(n799), .ZN(n724) );
  ND2D1 U44 ( .A1(n439), .A2(n445), .ZN(n676) );
  INVD1 U45 ( .I(n718), .ZN(n795) );
  ND2D1 U46 ( .A1(n853), .A2(n443), .ZN(n635) );
  ND2D1 U47 ( .A1(n442), .A2(a[6]), .ZN(n704) );
  ND2D2 U48 ( .A1(n440), .A2(n814), .ZN(n709) );
  ND2D1 U49 ( .A1(n439), .A2(n799), .ZN(n772) );
  ND2D1 U50 ( .A1(n681), .A2(n846), .ZN(n729) );
  ND2D1 U51 ( .A1(n799), .A2(n814), .ZN(n684) );
  ND2D1 U52 ( .A1(n443), .A2(n799), .ZN(n763) );
  OAI222D0 U53 ( .A1(n745), .A2(n718), .B1(n769), .B2(n581), .C1(n750), .C2(
        n760), .ZN(n585) );
  ND2D1 U54 ( .A1(a[1]), .A2(n437), .ZN(n718) );
  INVD1 U55 ( .I(n684), .ZN(n815) );
  ND2D1 U56 ( .A1(n846), .A2(n833), .ZN(n783) );
  INVD2 U57 ( .I(n751), .ZN(n846) );
  AOI21D2 U58 ( .A1(n815), .A2(a[1]), .B(n804), .ZN(n582) );
  INVD2 U59 ( .I(n704), .ZN(n849) );
  OAI31D1 U60 ( .A1(n704), .A2(n441), .A3(a[1]), .B(n635), .ZN(n554) );
  AOI21D1 U61 ( .A1(n797), .A2(n836), .B(n734), .ZN(n70) );
  OAI222D1 U62 ( .A1(a[1]), .A2(n776), .B1(n431), .B2(n757), .C1(n751), .C2(
        n747), .ZN(n485) );
  CKND2D1 U63 ( .A1(n849), .A2(n833), .ZN(n634) );
  ND2D1 U64 ( .A1(n830), .A2(n849), .ZN(n595) );
  NR2D1 U65 ( .A1(n461), .A2(n443), .ZN(n427) );
  CKND2D1 U66 ( .A1(n443), .A2(n444), .ZN(n430) );
  AOI22D2 U67 ( .A1(n831), .A2(n817), .B1(n806), .B2(n828), .ZN(n556) );
  CKND2D2 U68 ( .A1(n442), .A2(n835), .ZN(n757) );
  CKND2D1 U69 ( .A1(n443), .A2(n444), .ZN(n744) );
  ND2D1 U70 ( .A1(n831), .A2(n843), .ZN(n722) );
  AOI221D1 U71 ( .A1(n798), .A2(n687), .B1(n834), .B2(n800), .C(n686), .ZN(
        n688) );
  OA221D0 U72 ( .A1(n608), .A2(n583), .B1(n439), .B2(n774), .C(n701), .Z(n277)
         );
  CKND2 U73 ( .I(n765), .ZN(n833) );
  INVD2 U74 ( .I(n609), .ZN(n831) );
  INVD2 U75 ( .I(n780), .ZN(n843) );
  ND2D0 U76 ( .A1(n808), .A2(n443), .ZN(n705) );
  AOI211XD0 U77 ( .A1(n804), .A2(n824), .B(n827), .C(n695), .ZN(n696) );
  OA221D1 U78 ( .A1(n555), .A2(n629), .B1(n718), .B2(n784), .C(n342), .Z(n622)
         );
  OA222D1 U79 ( .A1(n640), .A2(n633), .B1(n589), .B2(n588), .C1(n587), .C2(
        n757), .Z(n342) );
  AO31D1 U80 ( .A1(n803), .A2(n860), .A3(n681), .B(n717), .Z(n459) );
  AOI221D1 U81 ( .A1(n862), .A2(n444), .B1(n844), .B2(n718), .C(n525), .ZN(
        n527) );
  INVD2 U82 ( .I(n757), .ZN(n860) );
  AOI221D1 U83 ( .A1(n861), .A2(n443), .B1(n853), .B2(n808), .C(n630), .ZN(
        n661) );
  OAI222D1 U84 ( .A1(n783), .A2(n581), .B1(n775), .B2(n635), .C1(n494), .C2(
        n763), .ZN(n495) );
  ND2D1 U85 ( .A1(n438), .A2(n814), .ZN(n775) );
  INVD3 U86 ( .I(n439), .ZN(n814) );
  AOI211XD1 U87 ( .A1(n830), .A2(n586), .B(n584), .C(n585), .ZN(n587) );
  CKND2D0 U88 ( .A1(n669), .A2(n849), .ZN(n588) );
  CKND2 U89 ( .I(N169), .ZN(n410) );
  INVD2 U90 ( .I(n410), .ZN(d[7]) );
  OAI22D1 U91 ( .A1(n445), .A2(n629), .B1(n628), .B2(n743), .ZN(n630) );
  ND4D2 U92 ( .A1(n478), .A2(n479), .A3(n477), .A4(n476), .ZN(N169) );
  AOI211XD0 U93 ( .A1(n844), .A2(n437), .B(n636), .C(n854), .ZN(n641) );
  OAI222D1 U94 ( .A1(n663), .A2(n768), .B1(n437), .B2(n556), .C1(n750), .C2(
        n555), .ZN(n557) );
  OR3D0 U95 ( .A1(n670), .A2(n812), .A3(n445), .Z(n631) );
  OAI221D1 U96 ( .A1(n665), .A2(n676), .B1(n664), .B2(n663), .C(n847), .ZN(
        n667) );
  ND2D1 U97 ( .A1(n443), .A2(n444), .ZN(n431) );
  AOI211XD0 U98 ( .A1(n864), .A2(n809), .B(n480), .C(n662), .ZN(n507) );
  OAI31D1 U99 ( .A1(n670), .A2(n800), .A3(n819), .B(n669), .ZN(n671) );
  OR2D0 U100 ( .A1(n677), .A2(n751), .Z(n433) );
  AOI221D1 U101 ( .A1(n848), .A2(n443), .B1(n858), .B2(a[1]), .C(n638), .ZN(
        n639) );
  AOI22D1 U102 ( .A1(n839), .A2(n806), .B1(n809), .B2(n838), .ZN(n467) );
  AOI221D1 U103 ( .A1(n700), .A2(n859), .B1(n817), .B2(n699), .C(n698), .ZN(
        n714) );
  AOI222D1 U104 ( .A1(n808), .A2(n831), .B1(n806), .B2(n482), .C1(n802), .C2(
        n834), .ZN(n487) );
  AOI221D1 U105 ( .A1(n857), .A2(n795), .B1(n860), .B2(n691), .C(n690), .ZN(
        n715) );
  OAI222D0 U106 ( .A1(n752), .A2(n761), .B1(n689), .B2(n720), .C1(n688), .C2(
        n780), .ZN(n690) );
  AOI221D2 U107 ( .A1(a[1]), .A2(n464), .B1(n827), .B2(n837), .C(n463), .ZN(
        n478) );
  OAI221D1 U108 ( .A1(n684), .A2(n673), .B1(n672), .B2(n785), .C(n671), .ZN(
        n674) );
  OA21D0 U109 ( .A1(n684), .A2(n443), .B(n612), .Z(n616) );
  OAI222D1 U110 ( .A1(n527), .A2(n775), .B1(n724), .B2(n623), .C1(n718), .C2(
        n526), .ZN(n539) );
  AOI221D1 U111 ( .A1(n830), .A2(n798), .B1(n822), .B2(n806), .C(n674), .ZN(
        n677) );
  CKND2D1 U112 ( .A1(n442), .A2(n828), .ZN(n727) );
  AOI221D1 U113 ( .A1(n837), .A2(n825), .B1(n823), .B2(n570), .C(n852), .ZN(
        n494) );
  INVD2 U114 ( .I(n752), .ZN(n801) );
  INVD0 U115 ( .I(n555), .ZN(n802) );
  ND4D2 U116 ( .A1(n716), .A2(n715), .A3(n714), .A4(n713), .ZN(d[1]) );
  CKND2D2 U117 ( .A1(n835), .A2(n840), .ZN(n751) );
  NR3D1 U118 ( .A1(n435), .A2(n436), .A3(n679), .ZN(n716) );
  AOI22D1 U119 ( .A1(n812), .A2(n833), .B1(n815), .B2(n828), .ZN(n764) );
  ND2D3 U120 ( .A1(n439), .A2(n438), .ZN(n640) );
  ND2D1 U121 ( .A1(n801), .A2(n437), .ZN(n555) );
  AOI32D0 U122 ( .A1(n442), .A2(n820), .A3(n801), .B1(n806), .B2(n448), .ZN(
        n449) );
  OAI33D0 U123 ( .A1(n752), .A2(n751), .A3(n750), .B1(n773), .B2(n799), .B3(
        n749), .ZN(n753) );
  ND2D0 U124 ( .A1(n801), .A2(n859), .ZN(n428) );
  ND2D2 U125 ( .A1(n438), .A2(n445), .ZN(n663) );
  ND2D2 U126 ( .A1(n437), .A2(n438), .ZN(n760) );
  INVD6 U127 ( .I(n440), .ZN(n820) );
  BUFFD8 U128 ( .I(a[4]), .Z(n440) );
  OAI222D1 U129 ( .A1(n567), .A2(n709), .B1(n566), .B2(n743), .C1(a[1]), .C2(
        n565), .ZN(n568) );
  AOI221D1 U130 ( .A1(n460), .A2(n808), .B1(n853), .B2(n818), .C(n459), .ZN(
        n461) );
  OAI222D1 U131 ( .A1(n811), .A2(n629), .B1(n552), .B2(n532), .C1(n531), .C2(
        n780), .ZN(n538) );
  IND4D2 U132 ( .A1(n793), .B1(n792), .B2(n791), .B3(n790), .ZN(d[0]) );
  ND4D2 U133 ( .A1(n622), .A2(n621), .A3(n620), .A4(n619), .ZN(d[3]) );
  ND2D1 U134 ( .A1(n439), .A2(n828), .ZN(n746) );
  INVD6 U135 ( .I(n441), .ZN(n828) );
  ND2D1 U136 ( .A1(a[6]), .A2(n828), .ZN(n773) );
  OAI222D1 U137 ( .A1(n560), .A2(n757), .B1(n684), .B2(n559), .C1(n751), .C2(
        n558), .ZN(n561) );
  NR4D1 U138 ( .A1(n539), .A2(n540), .A3(n538), .A4(n537), .ZN(n541) );
  OAI222D1 U139 ( .A1(n641), .A2(n640), .B1(n760), .B2(n762), .C1(n639), .C2(
        n772), .ZN(n642) );
  AOI221D1 U140 ( .A1(n846), .A2(n457), .B1(n456), .B2(n443), .C(n455), .ZN(
        n479) );
  AOI221D1 U141 ( .A1(n816), .A2(n599), .B1(n843), .B2(n598), .C(n597), .ZN(
        n621) );
  OAI221D1 U142 ( .A1(n738), .A2(n731), .B1(n704), .B2(n431), .C(n591), .ZN(
        n599) );
  NR4D1 U143 ( .A1(n789), .A2(n788), .A3(n787), .A4(n786), .ZN(n790) );
  OAI222D1 U144 ( .A1(n781), .A2(n780), .B1(n439), .B2(n841), .C1(n779), .C2(
        n443), .ZN(n787) );
  AOI221D1 U145 ( .A1(n823), .A2(n796), .B1(n832), .B2(n808), .C(n557), .ZN(
        n558) );
  ND4D2 U146 ( .A1(n507), .A2(n506), .A3(n505), .A4(n504), .ZN(d[6]) );
  AOI221D1 U147 ( .A1(n843), .A2(n496), .B1(n802), .B2(n509), .C(n495), .ZN(
        n505) );
  OAI33D0 U148 ( .A1(n654), .A2(n437), .A3(n799), .B1(n483), .B2(n727), .B3(
        n760), .ZN(n484) );
  CKAN2D0 U149 ( .A1(n719), .A2(n718), .Z(n723) );
  NR2D0 U150 ( .A1(n624), .A2(n718), .ZN(n700) );
  AOI221D1 U151 ( .A1(n801), .A2(n825), .B1(n809), .B2(n832), .C(n766), .ZN(
        n781) );
  AOI221D1 U152 ( .A1(n437), .A2(n563), .B1(n843), .B2(n562), .C(n561), .ZN(
        n579) );
  NR2D1 U153 ( .A1(n462), .A2(n749), .ZN(n425) );
  NR2D0 U154 ( .A1(n685), .A2(n513), .ZN(n426) );
  OR3D1 U155 ( .A1(n425), .A2(n426), .A3(n427), .Z(n463) );
  ND2D0 U156 ( .A1(n810), .A2(n838), .ZN(n429) );
  AN3XD1 U157 ( .A1(n428), .A2(n429), .A3(n70), .Z(n462) );
  INVD1 U158 ( .I(n760), .ZN(n810) );
  CKND2D0 U159 ( .A1(n800), .A2(n833), .ZN(n644) );
  OR2D0 U160 ( .A1(n437), .A2(n678), .Z(n432) );
  OR2D0 U161 ( .A1(n676), .A2(n675), .Z(n434) );
  ND2D0 U162 ( .A1(n831), .A2(n860), .ZN(n675) );
  NR2D0 U163 ( .A1(n751), .A2(n769), .ZN(n692) );
  ND3D1 U164 ( .A1(n432), .A2(n433), .A3(n434), .ZN(n679) );
  CKAN2D1 U165 ( .A1(n851), .A2(n810), .Z(n435) );
  CKAN2D1 U166 ( .A1(n692), .A2(n803), .Z(n436) );
  ND2D0 U167 ( .A1(n833), .A2(n840), .ZN(n623) );
  OAI22D0 U168 ( .A1(n765), .A2(n775), .B1(a[1]), .B2(n764), .ZN(n766) );
  AOI221D1 U169 ( .A1(n860), .A2(n643), .B1(n857), .B2(n803), .C(n642), .ZN(
        n660) );
  ND2D0 U170 ( .A1(a[1]), .A2(n439), .ZN(n782) );
  OAI22D0 U171 ( .A1(n765), .A2(n684), .B1(n689), .B2(n709), .ZN(n452) );
  CKBD4 U172 ( .I(a[7]), .Z(n442) );
  INVD1 U173 ( .I(n596), .ZN(n827) );
  CKND2D0 U174 ( .A1(n836), .A2(n825), .ZN(n532) );
  NR2D0 U175 ( .A1(n808), .A2(n795), .ZN(n612) );
  ND2D1 U176 ( .A1(n812), .A2(a[1]), .ZN(n581) );
  AOI21D1 U177 ( .A1(n862), .A2(n817), .B(n856), .ZN(n565) );
  INVD1 U178 ( .I(n640), .ZN(n817) );
  NR2XD0 U179 ( .A1(n834), .A2(n830), .ZN(n672) );
  CKND2D0 U180 ( .A1(n829), .A2(n849), .ZN(n633) );
  INVD0 U181 ( .I(n685), .ZN(n832) );
  NR2D0 U182 ( .A1(n623), .A2(n743), .ZN(n767) );
  AOI22D0 U183 ( .A1(n853), .A2(n523), .B1(n692), .B2(n522), .ZN(n524) );
  CKND2D0 U184 ( .A1(n823), .A2(n849), .ZN(n604) );
  INR2XD0 U185 ( .A1(n761), .B1(n498), .ZN(n499) );
  ND2D0 U186 ( .A1(n438), .A2(n820), .ZN(n624) );
  ND2D0 U187 ( .A1(n437), .A2(n806), .ZN(n728) );
  ND2D0 U188 ( .A1(n441), .A2(n840), .ZN(n706) );
  ND2D0 U189 ( .A1(n441), .A2(n835), .ZN(n508) );
  CKND2D0 U190 ( .A1(n773), .A2(n727), .ZN(n570) );
  INVD1 U191 ( .I(n635), .ZN(n854) );
  ND2D0 U192 ( .A1(n441), .A2(a[6]), .ZN(n776) );
  OAI33D0 U193 ( .A1(n755), .A2(n799), .A3(n727), .B1(n654), .B2(a[1]), .B3(
        n653), .ZN(n657) );
  AOI21D0 U194 ( .A1(n857), .A2(a[1]), .B(n692), .ZN(n693) );
  CKND2D0 U195 ( .A1(n816), .A2(a[1]), .ZN(n719) );
  NR2D0 U196 ( .A1(n805), .A2(n801), .ZN(n472) );
  CKND0 U197 ( .I(n774), .ZN(n861) );
  CKND0 U198 ( .I(n581), .ZN(n813) );
  OAI31D0 U200 ( .A1(n801), .A2(n797), .A3(n812), .B(n861), .ZN(n488) );
  AOI22D0 U201 ( .A1(n862), .A2(n803), .B1(n818), .B2(n848), .ZN(n546) );
  ND2D0 U202 ( .A1(n812), .A2(n855), .ZN(n564) );
  NR2D0 U203 ( .A1(n800), .A2(n796), .ZN(n613) );
  ND2D0 U204 ( .A1(n823), .A2(n863), .ZN(n761) );
  CKND2D0 U205 ( .A1(n822), .A2(n846), .ZN(n668) );
  ND2D0 U206 ( .A1(n798), .A2(n860), .ZN(n513) );
  NR2D0 U207 ( .A1(n717), .A2(n858), .ZN(n725) );
  CKND0 U208 ( .I(n720), .ZN(n845) );
  AOI211XD0 U210 ( .A1(n860), .A2(n492), .B(n491), .C(n490), .ZN(n506) );
  AOI21D0 U211 ( .A1(n821), .A2(n863), .B(n850), .ZN(n566) );
  AOI22D0 U212 ( .A1(n809), .A2(n859), .B1(n801), .B2(n838), .ZN(n567) );
  CKND2D0 U213 ( .A1(n728), .A2(n738), .ZN(n586) );
  NR2XD0 U214 ( .A1(n838), .A2(n849), .ZN(n637) );
  OAI22D0 U216 ( .A1(n443), .A2(n720), .B1(n445), .B2(n731), .ZN(n525) );
  CKND2D0 U217 ( .A1(n782), .A2(n552), .ZN(n553) );
  NR2D0 U218 ( .A1(n862), .A2(n848), .ZN(n458) );
  OAI211D0 U219 ( .A1(n828), .A2(n755), .B(n772), .C(n750), .ZN(n682) );
  CKND2D0 U220 ( .A1(n782), .A2(n684), .ZN(n522) );
  NR2XD0 U221 ( .A1(n844), .A2(n855), .ZN(n665) );
  OAI32D0 U222 ( .A1(n555), .A2(n757), .A3(n746), .B1(n514), .B2(n513), .ZN(
        n515) );
  NR2D0 U223 ( .A1(n833), .A2(n812), .ZN(n514) );
  ND2D0 U224 ( .A1(n843), .A2(n669), .ZN(n731) );
  CKND2D0 U225 ( .A1(n763), .A2(n760), .ZN(n748) );
  OAI22D0 U226 ( .A1(n640), .A2(n743), .B1(n430), .B2(n772), .ZN(n497) );
  OAI31D0 U227 ( .A1(n738), .A2(n824), .A3(n751), .B(n737), .ZN(n742) );
  AOI31D0 U228 ( .A1(n849), .A2(n736), .A3(n824), .B(n735), .ZN(n737) );
  NR2D0 U229 ( .A1(n812), .A2(n805), .ZN(n447) );
  OAI31D0 U230 ( .A1(n814), .A2(n804), .A3(n810), .B(n692), .ZN(n489) );
  AOI22D0 U231 ( .A1(n443), .A2(n818), .B1(n814), .B2(n805), .ZN(n589) );
  ND2D0 U232 ( .A1(n828), .A2(n840), .ZN(n608) );
  OAI21D0 U233 ( .A1(n750), .A2(n608), .B(n633), .ZN(n509) );
  CKND0 U234 ( .I(n750), .ZN(n824) );
  AOI32D0 U235 ( .A1(n801), .A2(n443), .A3(n834), .B1(n798), .B2(n548), .ZN(
        n550) );
  CKND2D0 U236 ( .A1(n750), .A2(n745), .ZN(n548) );
  OAI22D0 U237 ( .A1(n743), .A2(n755), .B1(n600), .B2(n430), .ZN(n607) );
  NR2D0 U238 ( .A1(n826), .A2(n831), .ZN(n600) );
  CKND2D0 U239 ( .A1(n831), .A2(n444), .ZN(n673) );
  NR2D0 U240 ( .A1(n443), .A2(n759), .ZN(n741) );
  CKND0 U241 ( .I(n709), .ZN(n825) );
  CKND2D0 U242 ( .A1(n681), .A2(n849), .ZN(n629) );
  CKND2D0 U243 ( .A1(n796), .A2(n814), .ZN(n721) );
  CKND0 U244 ( .I(n702), .ZN(n863) );
  CKND2D0 U245 ( .A1(n832), .A2(n849), .ZN(n762) );
  AOI21D0 U246 ( .A1(n807), .A2(n846), .B(n569), .ZN(n511) );
  NR2D0 U247 ( .A1(n440), .A2(n835), .ZN(n460) );
  CKND2D0 U248 ( .A1(n718), .A2(n814), .ZN(n572) );
  NR2D0 U249 ( .A1(n804), .A2(n807), .ZN(n573) );
  AOI22D0 U250 ( .A1(n826), .A2(n796), .B1(n824), .B2(n438), .ZN(n571) );
  CKND0 U251 ( .I(n736), .ZN(n811) );
  CKND2D0 U252 ( .A1(n817), .A2(n820), .ZN(n601) );
  AOI211D0 U253 ( .A1(n819), .A2(n437), .B(n817), .C(n810), .ZN(n602) );
  NR2XD0 U254 ( .A1(n645), .A2(n767), .ZN(n603) );
  AOI21D0 U255 ( .A1(n858), .A2(n818), .B(n694), .ZN(n697) );
  CKND2D0 U256 ( .A1(n685), .A2(n749), .ZN(n687) );
  OAI33D0 U257 ( .A1(n640), .A2(n442), .A3(n769), .B1(n702), .B2(n799), .B3(
        n750), .ZN(n533) );
  ND4D0 U258 ( .A1(n797), .A2(n837), .A3(n440), .A4(n442), .ZN(n726) );
  AOI31D0 U259 ( .A1(n438), .A2(n828), .A3(n797), .B(n827), .ZN(n493) );
  OAI211D0 U260 ( .A1(n702), .A2(n676), .B(n547), .C(n546), .ZN(n563) );
  OAI211D0 U261 ( .A1(n551), .A2(n718), .B(n550), .C(n549), .ZN(n562) );
  OAI32D0 U262 ( .A1(n768), .A2(n472), .A3(n704), .B1(n471), .B2(n738), .ZN(
        n475) );
  AOI31D0 U263 ( .A1(n440), .A2(n835), .A3(n812), .B(n694), .ZN(n471) );
  AOI21D0 U264 ( .A1(n775), .A2(n745), .B(n780), .ZN(n625) );
  AOI211D0 U265 ( .A1(n776), .A2(n654), .B(n583), .C(n743), .ZN(n473) );
  AOI33D0 U266 ( .A1(n610), .A2(n835), .A3(n803), .B1(n855), .B2(n814), .B3(
        n798), .ZN(n611) );
  OAI31D0 U267 ( .A1(n747), .A2(n776), .A3(n749), .B(n611), .ZN(n618) );
  OAI21D0 U268 ( .A1(n654), .A2(n749), .B(n729), .ZN(n535) );
  OAI22D0 U269 ( .A1(n445), .A2(n720), .B1(a[1]), .B2(n634), .ZN(n636) );
  OAI22D0 U270 ( .A1(n835), .A2(n709), .B1(n820), .B2(n654), .ZN(n646) );
  NR2D0 U272 ( .A1(n759), .A2(n437), .ZN(n711) );
  CKND0 U273 ( .I(n608), .ZN(n842) );
  OAI22D0 U274 ( .A1(n454), .A2(n780), .B1(n747), .B2(n633), .ZN(n455) );
  AOI21D0 U275 ( .A1(n684), .A2(n583), .B(n743), .ZN(n451) );
  AOI22D0 U276 ( .A1(n808), .A2(n437), .B1(a[1]), .B2(n817), .ZN(n481) );
  OAI22D0 U277 ( .A1(n442), .A2(n654), .B1(n750), .B2(n727), .ZN(n448) );
  NR2D0 U278 ( .A1(n858), .A2(n692), .ZN(n450) );
  CKND2D0 U279 ( .A1(n440), .A2(n799), .ZN(n583) );
  OAI21D0 U280 ( .A1(n708), .A2(n738), .B(n707), .ZN(n712) );
  CKND2D0 U281 ( .A1(n438), .A2(n738), .ZN(n736) );
  AOI21D0 U282 ( .A1(n439), .A2(n860), .B(n819), .ZN(n770) );
  CKND2D1 U283 ( .A1(n594), .A2(n593), .ZN(n598) );
  AOI21D0 U284 ( .A1(n848), .A2(n817), .B(n753), .ZN(n754) );
  NR2D0 U285 ( .A1(n810), .A2(n439), .ZN(n615) );
  AOI21D0 U286 ( .A1(n823), .A2(n859), .B(n694), .ZN(n501) );
  AOI32D0 U287 ( .A1(n440), .A2(n840), .A3(n816), .B1(n817), .B2(n545), .ZN(
        n547) );
  ND2D0 U288 ( .A1(a[1]), .A2(a[6]), .ZN(n483) );
  BUFFD4 U289 ( .I(a[5]), .Z(n441) );
  CKBD4 U290 ( .I(a[0]), .Z(n437) );
  INVD1 U291 ( .I(n783), .ZN(n848) );
  INVD1 U292 ( .I(n675), .ZN(n862) );
  INVD1 U293 ( .I(n564), .ZN(n856) );
  INVD1 U294 ( .I(n784), .ZN(n864) );
  ND2D1 U295 ( .A1(n669), .A2(n860), .ZN(n774) );
  NR2D1 U296 ( .A1(n634), .A2(n721), .ZN(n740) );
  INVD1 U297 ( .I(n588), .ZN(n858) );
  INVD1 U298 ( .I(n738), .ZN(n798) );
  AO221D0 U299 ( .A1(n801), .A2(n834), .B1(n798), .B2(n816), .C(n700), .Z(n651) );
  INVD1 U300 ( .I(n633), .ZN(n857) );
  INVD1 U301 ( .I(n763), .ZN(n805) );
  INVD1 U302 ( .I(n629), .ZN(n851) );
  INVD1 U303 ( .I(n431), .ZN(n796) );
  NR2D1 U304 ( .A1(n810), .A2(n808), .ZN(n465) );
  INVD1 U305 ( .I(n705), .ZN(n809) );
  ND2D1 U306 ( .A1(n863), .A2(n825), .ZN(n784) );
  INVD1 U307 ( .I(n634), .ZN(n855) );
  INVD1 U308 ( .I(n769), .ZN(n829) );
  INVD1 U309 ( .I(n755), .ZN(n822) );
  INVD1 U310 ( .I(n722), .ZN(n844) );
  ND2D1 U311 ( .A1(n795), .A2(n826), .ZN(n596) );
  ND2D1 U312 ( .A1(n821), .A2(n837), .ZN(n701) );
  NR2D1 U313 ( .A1(n817), .A2(n824), .ZN(n653) );
  INVD1 U314 ( .I(n595), .ZN(n852) );
  INVD1 U315 ( .I(n552), .ZN(n804) );
  INVD1 U316 ( .I(n551), .ZN(n821) );
  INVD1 U317 ( .I(n604), .ZN(n850) );
  OAI222D0 U318 ( .A1(n724), .A2(n749), .B1(n689), .B2(n685), .C1(n755), .C2(
        n552), .ZN(n530) );
  NR4D0 U319 ( .A1(n709), .A2(n763), .A3(n757), .A4(n828), .ZN(n735) );
  OAI32D1 U320 ( .A1(n583), .A2(n431), .A3(n685), .B1(n582), .B2(n765), .ZN(
        n584) );
  NR4D0 U321 ( .A1(n742), .A2(n741), .A3(n740), .A4(n739), .ZN(n791) );
  ND4D1 U322 ( .A1(n579), .A2(n580), .A3(n578), .A4(n577), .ZN(d[4]) );
  NR4D0 U323 ( .A1(n576), .A2(n575), .A3(n574), .A4(n739), .ZN(n577) );
  AOI221D0 U324 ( .A1(n812), .A2(n845), .B1(n853), .B2(n818), .C(n544), .ZN(
        n580) );
  INVD1 U325 ( .I(n749), .ZN(n823) );
  ND3D1 U326 ( .A1(n543), .A2(n542), .A3(n541), .ZN(d[5]) );
  AOI211D1 U327 ( .A1(n863), .A2(n517), .B(n516), .C(n515), .ZN(n543) );
  INR4D0 U328 ( .A1(n759), .B1(n521), .B2(n740), .B3(n710), .ZN(n542) );
  AOI221D0 U329 ( .A1(n843), .A2(n652), .B1(n846), .B2(n651), .C(n650), .ZN(
        n659) );
  NR4D0 U330 ( .A1(n657), .A2(n656), .A3(n655), .A4(n741), .ZN(n658) );
  ND2D1 U331 ( .A1(n489), .A2(n488), .ZN(n490) );
  OAI222D0 U332 ( .A1(n752), .A2(n685), .B1(n481), .B2(n765), .C1(a[1]), .C2(
        n750), .ZN(n492) );
  NR4D0 U333 ( .A1(n712), .A2(n735), .A3(n711), .A4(n710), .ZN(n713) );
  OAI221D0 U334 ( .A1(a[1]), .A2(n668), .B1(n721), .B2(n675), .C(n524), .ZN(
        n540) );
  INVD1 U335 ( .I(n782), .ZN(n818) );
  INVD1 U336 ( .I(n654), .ZN(n837) );
  ND2D1 U337 ( .A1(n843), .A2(n829), .ZN(n720) );
  NR4D0 U338 ( .A1(n475), .A2(n474), .A3(n711), .A4(n473), .ZN(n476) );
  NR2D1 U340 ( .A1(n618), .A2(n617), .ZN(n619) );
  NR3D0 U341 ( .A1(n718), .A2(n820), .A3(n729), .ZN(n574) );
  INVD1 U342 ( .I(n746), .ZN(n830) );
  INVD1 U343 ( .I(n727), .ZN(n859) );
  INVD1 U344 ( .I(n775), .ZN(n816) );
  INVD1 U345 ( .I(n743), .ZN(n797) );
  INVD1 U346 ( .I(n768), .ZN(n834) );
  NR2D1 U347 ( .A1(n706), .A2(n709), .ZN(n717) );
  NR2D1 U348 ( .A1(n702), .A2(n744), .ZN(n734) );
  INVD1 U349 ( .I(n676), .ZN(n819) );
  ND2D1 U350 ( .A1(n803), .A2(n443), .ZN(n552) );
  OAI221D0 U351 ( .A1(n458), .A2(n775), .B1(n720), .B2(n772), .C(n564), .ZN(
        n464) );
  INVD1 U352 ( .I(n703), .ZN(n826) );
  INVD1 U353 ( .I(n728), .ZN(n807) );
  INVD1 U354 ( .I(n508), .ZN(n836) );
  OAI222D0 U355 ( .A1(n760), .A2(n768), .B1(n782), .B2(n644), .C1(n749), .C2(
        n705), .ZN(n652) );
  OAI221D0 U356 ( .A1(n447), .A2(n609), .B1(n775), .B2(n718), .C(n446), .ZN(
        n457) );
  AOI221D0 U357 ( .A1(n797), .A2(n682), .B1(n681), .B2(n806), .C(n680), .ZN(
        n683) );
  INVD1 U358 ( .I(n724), .ZN(n800) );
  OAI222D0 U359 ( .A1(n746), .A2(n552), .B1(n640), .B2(n718), .C1(n747), .C2(
        n685), .ZN(n453) );
  NR3D0 U360 ( .A1(n738), .A2(n439), .A3(n765), .ZN(n529) );
  OAI222D0 U361 ( .A1(n730), .A2(n719), .B1(n697), .B2(n443), .C1(n696), .C2(
        n773), .ZN(n698) );
  NR4D0 U362 ( .A1(a[1]), .A2(n840), .A3(n763), .A4(n755), .ZN(n695) );
  INVD1 U363 ( .I(n767), .ZN(n841) );
  AOI221D0 U364 ( .A1(n795), .A2(n815), .B1(n802), .B2(n830), .C(n592), .ZN(
        n593) );
  AOI222D0 U365 ( .A1(n803), .A2(n822), .B1(n824), .B2(n805), .C1(n807), .C2(
        n441), .ZN(n594) );
  OAI222D0 U366 ( .A1(n472), .A2(n706), .B1(n465), .B2(n704), .C1(n727), .C2(
        n728), .ZN(n469) );
  OAI222D0 U367 ( .A1(n438), .A2(n649), .B1(n648), .B2(n784), .C1(n647), .C2(
        n783), .ZN(n650) );
  AOI21D1 U368 ( .A1(n795), .A2(n646), .B(n645), .ZN(n649) );
  OAI222D0 U369 ( .A1(n705), .A2(n731), .B1(n437), .B2(n536), .C1(n785), .C2(
        n774), .ZN(n537) );
  AOI221D0 U370 ( .A1(n806), .A2(n535), .B1(n846), .B2(n534), .C(n533), .ZN(
        n536) );
  OAI21D1 U371 ( .A1(n437), .A2(n685), .B(n749), .ZN(n482) );
  OAI222D0 U372 ( .A1(n442), .A2(n771), .B1(n770), .B2(n769), .C1(n780), .C2(
        n768), .ZN(n778) );
  OAI222D0 U373 ( .A1(n776), .A2(n785), .B1(n775), .B2(n774), .C1(n773), .C2(
        n772), .ZN(n777) );
  OAI222D0 U374 ( .A1(n512), .A2(n743), .B1(n511), .B2(n750), .C1(n510), .C2(
        n763), .ZN(n516) );
  NR2D1 U375 ( .A1(n861), .A2(n509), .ZN(n510) );
  OAI222D0 U376 ( .A1(n501), .A2(n431), .B1(n820), .B2(n500), .C1(n499), .C2(
        n718), .ZN(n503) );
  ND2D1 U377 ( .A1(n442), .A2(n497), .ZN(n500) );
  OAI221D0 U378 ( .A1(n613), .A2(n765), .B1(n750), .B2(n760), .C(n493), .ZN(
        n496) );
  NR4D0 U379 ( .A1(n453), .A2(n452), .A3(n528), .A4(n451), .ZN(n454) );
  OAI221D0 U380 ( .A1(n450), .A2(n640), .B1(n772), .B2(n731), .C(n449), .ZN(
        n456) );
  INR4D0 U381 ( .A1(n668), .B1(n667), .B2(n666), .B3(n856), .ZN(n678) );
  OAI221D0 U382 ( .A1(n750), .A2(n752), .B1(n709), .B2(n785), .C(n632), .ZN(
        n643) );
  OAI221D0 U383 ( .A1(n443), .A2(n731), .B1(n704), .B2(n718), .C(n693), .ZN(
        n699) );
  NR4D0 U384 ( .A1(n503), .A2(n502), .A3(n518), .A4(n519), .ZN(n504) );
  OAI222D0 U385 ( .A1(n758), .A2(n757), .B1(n756), .B2(n755), .C1(n437), .C2(
        n754), .ZN(n789) );
  OAI222D0 U386 ( .A1(n763), .A2(n762), .B1(n761), .B2(n760), .C1(a[1]), .C2(
        n759), .ZN(n788) );
  NR4D0 U387 ( .A1(n627), .A2(n626), .A3(n850), .A4(n625), .ZN(n628) );
  NR3D0 U388 ( .A1(n738), .A2(n440), .A3(n608), .ZN(n645) );
  ND2D1 U389 ( .A1(n441), .A2(n442), .ZN(n702) );
  NR4D0 U390 ( .A1(n437), .A2(n835), .A3(n769), .A4(n775), .ZN(n575) );
  NR3D0 U391 ( .A1(n775), .A2(n442), .A3(n440), .ZN(n666) );
  ND2D1 U392 ( .A1(n441), .A2(n820), .ZN(n765) );
  NR3D0 U393 ( .A1(n443), .A2(n440), .A3(n685), .ZN(n592) );
  OAI221D0 U394 ( .A1(n738), .A2(n727), .B1(a[1]), .B2(n783), .C(n726), .ZN(
        n733) );
  NR3D0 U395 ( .A1(n704), .A2(n828), .A3(n709), .ZN(n520) );
  OAI222D0 U396 ( .A1(n573), .A2(n774), .B1(n783), .B2(n572), .C1(n571), .C2(
        n776), .ZN(n576) );
  ND2D1 U397 ( .A1(n438), .A2(n441), .ZN(n745) );
  AOI211XD0 U398 ( .A1(n842), .A2(n809), .B(n485), .C(n484), .ZN(n486) );
  NR3D0 U399 ( .A1(n719), .A2(n440), .A3(n840), .ZN(n656) );
  ND2D1 U400 ( .A1(n440), .A2(n439), .ZN(n750) );
  ND2D1 U401 ( .A1(n440), .A2(n828), .ZN(n609) );
  INVD1 U402 ( .I(n437), .ZN(n794) );
  INVD1 U403 ( .I(n773), .ZN(n838) );
  OAI222D0 U404 ( .A1(n616), .A2(n774), .B1(n615), .B2(n722), .C1(n614), .C2(
        n755), .ZN(n617) );
  OA22D0 U405 ( .A1(n776), .A2(n743), .B1(n727), .B2(n613), .Z(n614) );
  ND2D1 U406 ( .A1(n440), .A2(n438), .ZN(n703) );
  OAI222D0 U407 ( .A1(n634), .A2(n799), .B1(n608), .B2(n601), .C1(n439), .C2(
        n720), .ZN(n606) );
  INVD1 U408 ( .I(n776), .ZN(n839) );
  INVD1 U409 ( .I(n442), .ZN(n840) );
  OAI222D0 U410 ( .A1(n757), .A2(n624), .B1(n439), .B2(n623), .C1(n751), .C2(
        n768), .ZN(n627) );
  NR4D0 U411 ( .A1(a[6]), .A2(n814), .A3(n727), .A4(n760), .ZN(n502) );
  OAI222D0 U412 ( .A1(n640), .A2(n722), .B1(n589), .B2(n731), .C1(n634), .C2(
        n663), .ZN(n480) );
  ND4D1 U413 ( .A1(n660), .A2(n661), .A3(n659), .A4(n658), .ZN(d[2]) );
  AN2XD1 U414 ( .A1(n437), .A2(n814), .Z(n670) );
  NR3D0 U415 ( .A1(n670), .A2(n801), .A3(n816), .ZN(n647) );
  OAI22D0 U416 ( .A1(n755), .A2(n752), .B1(n653), .B2(n738), .ZN(n517) );
  OAI222D0 U417 ( .A1(n752), .A2(n604), .B1(n603), .B2(n799), .C1(n602), .C2(
        n675), .ZN(n605) );
  NR4D0 U418 ( .A1(n685), .A2(n752), .A3(n780), .A4(n820), .ZN(n655) );
  OA33D0 U419 ( .A1(n706), .A2(n750), .A3(n743), .B1(n705), .B2(n704), .B3(
        n768), .Z(n707) );
  ND3D0 U420 ( .A1(n817), .A2(n669), .A3(n846), .ZN(n759) );
  AN4D1 U421 ( .A1(n669), .A2(n818), .A3(n437), .A4(n846), .Z(n518) );
  NR2D1 U422 ( .A1(n820), .A2(n828), .ZN(n669) );
  NR3D0 U423 ( .A1(n508), .A2(n750), .A3(n785), .ZN(n474) );
  OAI22D0 U424 ( .A1(n785), .A2(n784), .B1(n783), .B2(n782), .ZN(n786) );
  OAI222D0 U425 ( .A1(n725), .A2(n724), .B1(n723), .B2(n722), .C1(n721), .C2(
        n720), .ZN(n793) );
  AOI21D0 U426 ( .A1(n685), .A2(n765), .B(n724), .ZN(n680) );
  OAI222D0 U427 ( .A1(n727), .A2(n596), .B1(n724), .B2(n762), .C1(n612), .C2(
        n595), .ZN(n597) );
  OAI222D0 U428 ( .A1(n724), .A2(n595), .B1(n731), .B2(n676), .C1(n634), .C2(
        n760), .ZN(n544) );
  CKND2D0 U429 ( .A1(n724), .A2(n752), .ZN(n523) );
  NR3D0 U430 ( .A1(n828), .A2(a[1]), .A3(n724), .ZN(n528) );
  AOI221D0 U431 ( .A1(n734), .A2(n816), .B1(n815), .B2(n733), .C(n732), .ZN(
        n792) );
  AOI221D0 U432 ( .A1(n804), .A2(n834), .B1(n829), .B2(n553), .C(n700), .ZN(
        n560) );
  INR2D1 U433 ( .A1(n520), .B1(n663), .ZN(n710) );
  NR4D0 U434 ( .A1(n769), .A2(n757), .A3(n663), .A4(n439), .ZN(n739) );
  AOI22D0 U435 ( .A1(n837), .A2(n748), .B1(n839), .B2(n806), .ZN(n756) );
  NR2D1 U436 ( .A1(n508), .A2(n663), .ZN(n569) );
  NR2D1 U437 ( .A1(n796), .A2(n806), .ZN(n648) );
  CKND1 U438 ( .I(n662), .ZN(n847) );
  AOI32D1 U439 ( .A1(n441), .A2(n443), .A3(n818), .B1(n829), .B2(n631), .ZN(
        n632) );
  OA222D0 U440 ( .A1(n747), .A2(n746), .B1(n745), .B2(n431), .C1(n749), .C2(
        n743), .Z(n758) );
  AOI22D0 U441 ( .A1(n830), .A2(n806), .B1(n803), .B2(n832), .ZN(n446) );
  OAI22D0 U442 ( .A1(a[6]), .A2(n440), .B1(n441), .B2(n757), .ZN(n545) );
  OAI211D0 U443 ( .A1(n441), .A2(n782), .B(n624), .C(n749), .ZN(n534) );
  OAI22D0 U444 ( .A1(n746), .A2(n752), .B1(n765), .B2(n785), .ZN(n686) );
  NR2D1 U445 ( .A1(n439), .A2(n441), .ZN(n681) );
  AOI222D0 U446 ( .A1(n808), .A2(n825), .B1(n823), .B2(n800), .C1(n832), .C2(
        n806), .ZN(n549) );
  AOI21D1 U447 ( .A1(n834), .A2(n843), .B(n852), .ZN(n664) );
  OAI22D1 U448 ( .A1(n722), .A2(n752), .B1(n799), .B2(n729), .ZN(n662) );
  OAI21D0 U449 ( .A1(n640), .A2(n730), .B(n784), .ZN(n470) );
  AOI31D0 U450 ( .A1(n731), .A2(n730), .A3(n729), .B(n728), .ZN(n732) );
  OAI22D0 U451 ( .A1(n439), .A2(n609), .B1(n443), .B2(n608), .ZN(n610) );
  AOI21D0 U452 ( .A1(n609), .A2(n654), .B(n684), .ZN(n498) );
  OAI21D0 U453 ( .A1(n751), .A2(n609), .B(n720), .ZN(n590) );
endmodule


module aes_sbox_13 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n18, n68, n70, n74, n77, n78, n79, n80, n100, n123, n196, n204, n245,
         n277, n287, n304, n305, n306, n405, n408, n409, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862;

  AN2XD1 U28 ( .A1(n726), .A2(n725), .Z(n730) );
  OA21D1 U35 ( .A1(n710), .A2(n709), .B(n708), .Z(n715) );
  OR4D1 U199 ( .A1(n664), .A2(n585), .A3(n532), .A4(n531), .Z(n534) );
  AN2XD1 U215 ( .A1(n533), .A2(n809), .Z(n532) );
  AN2XD1 U271 ( .A1(n546), .A2(n738), .Z(n479) );
  AO21D1 U297 ( .A1(n80), .A2(n835), .B(n741), .Z(n474) );
  AOI211XD0 U1 ( .A1(n858), .A2(n505), .B(n504), .C(n503), .ZN(n519) );
  ND2D2 U2 ( .A1(n851), .A2(n456), .ZN(n644) );
  AOI221D1 U3 ( .A1(n699), .A2(n750), .B1(n457), .B2(n853), .C(n568), .ZN(n573) );
  ND4D2 U4 ( .A1(n669), .A2(n670), .A3(n668), .A4(n667), .ZN(d[2]) );
  INVD1 U5 ( .I(n777), .ZN(n811) );
  OA221D1 U6 ( .A1(n758), .A2(n716), .B1(n712), .B2(n692), .C(n196), .Z(n786)
         );
  OAI221D1 U7 ( .A1(n465), .A2(n440), .B1(n777), .B2(n738), .C(n464), .ZN(n471) );
  ND2D3 U8 ( .A1(n456), .A2(n459), .ZN(n750) );
  OAI31D2 U9 ( .A1(n444), .A2(n799), .A3(n818), .B(n677), .ZN(n678) );
  AOI221D0 U10 ( .A1(n797), .A2(n694), .B1(n833), .B2(n799), .C(n693), .ZN(
        n695) );
  CKND2D0 U11 ( .A1(n799), .A2(n832), .ZN(n653) );
  INVD2 U12 ( .I(n731), .ZN(n799) );
  OAI221D1 U13 ( .A1(n70), .A2(n680), .B1(n679), .B2(n790), .C(n678), .ZN(n681) );
  INVD1 U14 ( .I(n671), .ZN(n805) );
  CKND2D1 U15 ( .A1(n451), .A2(n460), .ZN(n671) );
  ND2D2 U16 ( .A1(n802), .A2(n456), .ZN(n566) );
  OAI22D1 U17 ( .A1(n469), .A2(n785), .B1(n753), .B2(n642), .ZN(n470) );
  AOI21D2 U18 ( .A1(n814), .A2(n457), .B(n803), .ZN(n592) );
  AOI221D2 U19 ( .A1(n849), .A2(n809), .B1(n699), .B2(n802), .C(n686), .ZN(
        n723) );
  ND2D2 U20 ( .A1(n834), .A2(n839), .ZN(n757) );
  ND2D0 U21 ( .A1(n454), .A2(n839), .ZN(n713) );
  CKND2D0 U22 ( .A1(n827), .A2(n839), .ZN(n618) );
  CKND2D0 U23 ( .A1(n832), .A2(n839), .ZN(n632) );
  INVD2 U24 ( .I(n757), .ZN(n845) );
  AOI221D1 U25 ( .A1(n812), .A2(n581), .B1(n580), .B2(n822), .C(n579), .ZN(
        n589) );
  NR4D1 U26 ( .A1(n468), .A2(n467), .A3(n542), .A4(n466), .ZN(n469) );
  INR4D2 U27 ( .A1(n676), .B1(n674), .B2(n675), .B3(n854), .ZN(n685) );
  ND4D2 U29 ( .A1(n723), .A2(n722), .A3(n721), .A4(n720), .ZN(d[1]) );
  AOI221D1 U30 ( .A1(n835), .A2(n795), .B1(n600), .B2(n459), .C(n741), .ZN(
        n601) );
  OAI21D0 U31 ( .A1(n757), .A2(n619), .B(n727), .ZN(n600) );
  OAI221D2 U32 ( .A1(n673), .A2(n683), .B1(n672), .B2(n671), .C(n439), .ZN(
        n675) );
  OA22D2 U33 ( .A1(n729), .A2(n758), .B1(n798), .B2(n736), .Z(n439) );
  INVD2 U34 ( .I(n691), .ZN(n18) );
  CKND2 U36 ( .I(n18), .ZN(n68) );
  CKND0 U37 ( .I(n18), .ZN(n70) );
  CKND0 U38 ( .I(n18), .ZN(n74) );
  CKBD1 U39 ( .I(n755), .Z(n77) );
  CKBD0 U40 ( .I(n755), .Z(n78) );
  BUFFD1 U41 ( .I(n755), .Z(n79) );
  INVD2 U42 ( .I(n711), .ZN(n847) );
  INVD1 U43 ( .I(n766), .ZN(n809) );
  CKND1 U44 ( .I(a[1]), .ZN(n460) );
  ND2D1 U45 ( .A1(n813), .A2(n819), .ZN(n761) );
  INVD1 U46 ( .I(n758), .ZN(n800) );
  INVD2 U47 ( .I(n790), .ZN(n802) );
  ND2D0 U48 ( .A1(n452), .A2(n819), .ZN(n755) );
  CKND2D1 U49 ( .A1(n455), .A2(n827), .ZN(n734) );
  AOI221D1 U50 ( .A1(n845), .A2(n617), .B1(n616), .B2(n456), .C(n615), .ZN(
        n630) );
  CKBD4 U51 ( .I(n794), .Z(n456) );
  NR3D0 U52 ( .A1(n571), .A2(n434), .A3(n433), .ZN(n572) );
  INVD1 U53 ( .I(n773), .ZN(n833) );
  INVD1 U54 ( .I(n455), .ZN(n839) );
  INVD2 U55 ( .I(n619), .ZN(n830) );
  CKND2D1 U56 ( .A1(n450), .A2(n798), .ZN(n731) );
  OAI222D0 U57 ( .A1(n751), .A2(n725), .B1(n774), .B2(n591), .C1(n756), .C2(
        n766), .ZN(n595) );
  INVD1 U58 ( .I(n643), .ZN(n853) );
  BUFFD3 U59 ( .I(a[7]), .Z(n455) );
  ND2D0 U60 ( .A1(n811), .A2(n853), .ZN(n575) );
  ND2D1 U61 ( .A1(n827), .A2(n834), .ZN(n663) );
  ND2D2 U62 ( .A1(n455), .A2(a[6]), .ZN(n711) );
  INVD1 U63 ( .I(n753), .ZN(n807) );
  OAI221D0 U64 ( .A1(n756), .A2(n758), .B1(n716), .B2(n790), .C(n641), .ZN(
        n652) );
  ND4D1 U65 ( .A1(n520), .A2(n519), .A3(n518), .A4(n517), .ZN(d[6]) );
  OA221D1 U66 ( .A1(n569), .A2(n638), .B1(n725), .B2(n789), .C(n408), .Z(n631)
         );
  OAI22D1 U67 ( .A1(n750), .A2(n713), .B1(n646), .B2(n745), .ZN(n647) );
  OA22D0 U68 ( .A1(n771), .A2(n780), .B1(n457), .B2(n770), .Z(n196) );
  AOI22D1 U69 ( .A1(n811), .A2(n832), .B1(n814), .B2(n827), .ZN(n770) );
  OAI222D0 U70 ( .A1(n455), .A2(n776), .B1(n775), .B2(n774), .C1(n785), .C2(
        n773), .ZN(n783) );
  AOI221D0 U71 ( .A1(n795), .A2(n814), .B1(n801), .B2(n829), .C(n602), .ZN(
        n603) );
  ND2D1 U72 ( .A1(n819), .A2(n827), .ZN(n774) );
  INVD1 U73 ( .I(n771), .ZN(n832) );
  ND2D1 U74 ( .A1(n452), .A2(n827), .ZN(n752) );
  ND2D1 U75 ( .A1(n847), .A2(n832), .ZN(n643) );
  AOI222D1 U76 ( .A1(n807), .A2(n830), .B1(n805), .B2(n495), .C1(n801), .C2(
        n833), .ZN(n500) );
  ND2D2 U77 ( .A1(n454), .A2(n819), .ZN(n771) );
  OAI222D0 U78 ( .A1(n752), .A2(n566), .B1(n440), .B2(n725), .C1(n753), .C2(
        n692), .ZN(n468) );
  ND2D1 U79 ( .A1(n453), .A2(n827), .ZN(n619) );
  OR2D1 U80 ( .A1(n453), .A2(n834), .Z(n204) );
  NR3D0 U81 ( .A1(n409), .A2(n424), .A3(n474), .ZN(n476) );
  ND2D2 U82 ( .A1(n457), .A2(n456), .ZN(n745) );
  OAI222D0 U83 ( .A1(n578), .A2(n716), .B1(n577), .B2(n435), .C1(n457), .C2(
        n576), .ZN(n579) );
  OA221D0 U84 ( .A1(n456), .A2(n441), .B1(n785), .B2(n442), .C(n443), .Z(n590)
         );
  INVD1 U85 ( .I(n68), .ZN(n814) );
  NR3D0 U86 ( .A1(n425), .A2(n426), .A3(n427), .ZN(n408) );
  ND2D1 U87 ( .A1(n458), .A2(n450), .ZN(n725) );
  MAOI22D1 U88 ( .A1(n856), .A2(n813), .B1(n633), .B2(n778), .ZN(n525) );
  OAI222D0 U89 ( .A1(n485), .A2(n713), .B1(n478), .B2(n711), .C1(n734), .C2(
        n735), .ZN(n482) );
  INVD1 U90 ( .I(n80), .ZN(n435) );
  ND2D1 U91 ( .A1(n460), .A2(n798), .ZN(n758) );
  AN2XD1 U92 ( .A1(n450), .A2(n459), .Z(n80) );
  AO221D1 U93 ( .A1(n815), .A2(n609), .B1(n842), .B2(n608), .C(n607), .Z(n100)
         );
  BUFFD2 U94 ( .I(n649), .Z(n440) );
  NR2XD0 U95 ( .A1(n783), .A2(n782), .ZN(n784) );
  NR2D1 U96 ( .A1(n784), .A2(n456), .ZN(n432) );
  BUFFD1 U97 ( .I(n731), .Z(n123) );
  INVD2 U98 ( .I(n452), .ZN(n813) );
  AN4XD1 U99 ( .A1(n277), .A2(n287), .A3(n304), .A4(n305), .Z(n791) );
  INVD2 U100 ( .I(n440), .ZN(n816) );
  NR2D1 U101 ( .A1(n794), .A2(n452), .ZN(n444) );
  ND4D2 U102 ( .A1(n492), .A2(n491), .A3(n490), .A4(n489), .ZN(d[7]) );
  AOI31D1 U103 ( .A1(n802), .A2(n858), .A3(n688), .B(n724), .ZN(n245) );
  CKND2D1 U104 ( .A1(n452), .A2(n460), .ZN(n683) );
  INVD1 U105 ( .I(n683), .ZN(n818) );
  CKND2D0 U106 ( .A1(n457), .A2(n452), .ZN(n787) );
  INVD2 U107 ( .I(n459), .ZN(n457) );
  OAI211D1 U108 ( .A1(n454), .A2(n787), .B(n633), .C(n78), .ZN(n548) );
  NR2XD0 U109 ( .A1(n799), .A2(n80), .ZN(n696) );
  OAI222D0 U110 ( .A1(n731), .A2(n79), .B1(n696), .B2(n692), .C1(n761), .C2(
        n566), .ZN(n544) );
  OA211D0 U111 ( .A1(n709), .A2(n683), .B(n561), .C(n560), .Z(n441) );
  OA221D1 U112 ( .A1(n204), .A2(n753), .B1(n737), .B2(n787), .C(n245), .Z(n475) );
  INVD1 U113 ( .I(n787), .ZN(n817) );
  NR3D1 U114 ( .A1(n430), .A2(n431), .A3(n432), .ZN(n304) );
  CKND2D0 U115 ( .A1(n123), .A2(n758), .ZN(n536) );
  ND2D0 U116 ( .A1(n456), .A2(n798), .ZN(n769) );
  CKND2D1 U117 ( .A1(n451), .A2(n813), .ZN(n780) );
  IND4D1 U118 ( .A1(n449), .B1(n590), .B2(n589), .B3(n588), .ZN(d[4]) );
  AOI221D1 U119 ( .A1(n858), .A2(n652), .B1(n855), .B2(n802), .C(n651), .ZN(
        n669) );
  INVD2 U120 ( .I(n737), .ZN(n851) );
  ND2D2 U121 ( .A1(n830), .A2(n847), .ZN(n737) );
  OA222D0 U122 ( .A1(n764), .A2(n763), .B1(n762), .B2(n761), .C1(n450), .C2(
        n760), .Z(n277) );
  OA222D0 U123 ( .A1(n769), .A2(n768), .B1(n767), .B2(n766), .C1(n457), .C2(
        n765), .Z(n287) );
  OA22D0 U124 ( .A1(n790), .A2(n789), .B1(n788), .B2(n787), .Z(n305) );
  CKND2 U125 ( .I(n100), .ZN(n306) );
  ND4D4 U126 ( .A1(n631), .A2(n306), .A3(n630), .A4(n629), .ZN(d[3]) );
  INVD1 U127 ( .I(n569), .ZN(n801) );
  OAI33D0 U128 ( .A1(n761), .A2(n798), .A3(n734), .B1(n663), .B2(n457), .B3(
        n662), .ZN(n666) );
  ND2D1 U129 ( .A1(n454), .A2(n813), .ZN(n773) );
  INVD2 U130 ( .I(n451), .ZN(n798) );
  OAI222D0 U131 ( .A1(n758), .A2(n614), .B1(n613), .B2(n798), .C1(n612), .C2(
        n682), .ZN(n615) );
  ND2D0 U132 ( .A1(n450), .A2(n805), .ZN(n735) );
  NR2XD0 U133 ( .A1(n804), .A2(n800), .ZN(n485) );
  IIND4D2 U134 ( .A1(n793), .A2(n405), .B1(n791), .B2(n792), .ZN(d[0]) );
  AO221D0 U135 ( .A1(n741), .A2(n815), .B1(n814), .B2(n740), .C(n739), .Z(n405) );
  NR2D1 U136 ( .A1(n597), .A2(n763), .ZN(n427) );
  OAI222D1 U137 ( .A1(n541), .A2(n780), .B1(n123), .B2(n632), .C1(n540), .C2(
        n725), .ZN(n553) );
  AOI221D1 U138 ( .A1(n707), .A2(n857), .B1(n816), .B2(n706), .C(n705), .ZN(
        n721) );
  OAI222D1 U139 ( .A1(n123), .A2(n546), .B1(n500), .B2(n757), .C1(n499), .C2(
        n761), .ZN(n504) );
  NR2D1 U140 ( .A1(n819), .A2(n827), .ZN(n677) );
  CKND2D0 U141 ( .A1(n787), .A2(n74), .ZN(n535) );
  AOI221D1 U142 ( .A1(n805), .A2(n549), .B1(n845), .B2(n548), .C(n547), .ZN(
        n550) );
  AOI221D1 U143 ( .A1(n842), .A2(n661), .B1(n845), .B2(n660), .C(n659), .ZN(
        n668) );
  OA222D0 U144 ( .A1(n753), .A2(n752), .B1(n751), .B2(n750), .C1(n78), .C2(
        n435), .Z(n764) );
  ND2D1 U145 ( .A1(n458), .A2(n451), .ZN(n753) );
  AOI211D1 U146 ( .A1(n841), .A2(n808), .B(n498), .C(n497), .ZN(n499) );
  AN2D1 U147 ( .A1(n822), .A2(n796), .Z(n433) );
  ND2D1 U148 ( .A1(n822), .A2(n847), .ZN(n614) );
  ND2D1 U149 ( .A1(n822), .A2(n861), .ZN(n767) );
  ND2D1 U150 ( .A1(n452), .A2(n798), .ZN(n777) );
  ND2D1 U151 ( .A1(n798), .A2(n813), .ZN(n691) );
  AOI211XD0 U152 ( .A1(n862), .A2(n808), .B(n493), .C(n445), .ZN(n520) );
  OR3D1 U153 ( .A1(n444), .A2(n811), .A3(n460), .Z(n640) );
  ND2D1 U154 ( .A1(n811), .A2(n457), .ZN(n591) );
  NR2D0 U155 ( .A1(n811), .A2(n804), .ZN(n462) );
  NR2D0 U156 ( .A1(n832), .A2(n811), .ZN(n527) );
  OAI222D1 U157 ( .A1(n671), .A2(n773), .B1(n450), .B2(n570), .C1(n756), .C2(
        n569), .ZN(n571) );
  OAI31D1 U158 ( .A1(n711), .A2(n454), .A3(n457), .B(n644), .ZN(n568) );
  AOI221D1 U159 ( .A1(n803), .A2(n833), .B1(n828), .B2(n567), .C(n707), .ZN(
        n574) );
  NR4D1 U160 ( .A1(n552), .A2(n553), .A3(n554), .A4(n551), .ZN(n555) );
  ND3D2 U161 ( .A1(n555), .A2(n556), .A3(n557), .ZN(d[5]) );
  NR2D1 U162 ( .A1(n786), .A2(n785), .ZN(n430) );
  AOI211XD1 U163 ( .A1(n829), .A2(n596), .B(n595), .C(n594), .ZN(n597) );
  OR2XD1 U164 ( .A1(n475), .A2(n456), .Z(n448) );
  AOI221D1 U165 ( .A1(n845), .A2(n472), .B1(n471), .B2(n456), .C(n470), .ZN(
        n492) );
  AOI222D1 U166 ( .A1(n802), .A2(n821), .B1(n823), .B2(n804), .C1(n806), .C2(
        n454), .ZN(n604) );
  AOI22D1 U167 ( .A1(n456), .A2(n817), .B1(n813), .B2(n804), .ZN(n599) );
  AOI221D1 U168 ( .A1(n846), .A2(n456), .B1(n856), .B2(n457), .C(n647), .ZN(
        n648) );
  AOI221D1 U169 ( .A1(n855), .A2(n795), .B1(n858), .B2(n698), .C(n697), .ZN(
        n722) );
  AOI221D1 U170 ( .A1(n483), .A2(n459), .B1(n821), .B2(n482), .C(n481), .ZN(
        n490) );
  CKND4 U171 ( .I(a[1]), .ZN(n459) );
  INVD3 U172 ( .I(n459), .ZN(n458) );
  OAI222D1 U173 ( .A1(n650), .A2(n440), .B1(n766), .B2(n768), .C1(n648), .C2(
        n777), .ZN(n651) );
  OA21D0 U174 ( .A1(n74), .A2(n456), .B(n622), .Z(n626) );
  AOI221D1 U175 ( .A1(n829), .A2(n797), .B1(n821), .B2(n805), .C(n681), .ZN(
        n684) );
  INVD4 U176 ( .I(n453), .ZN(n819) );
  AOI221D1 U177 ( .A1(n859), .A2(n456), .B1(n851), .B2(n807), .C(n639), .ZN(
        n670) );
  OAI22D0 U178 ( .A1(n460), .A2(n638), .B1(n637), .B2(n435), .ZN(n639) );
  INVD6 U179 ( .I(n454), .ZN(n827) );
  OAI222D1 U180 ( .A1(n450), .A2(n685), .B1(n757), .B2(n684), .C1(n683), .C2(
        n682), .ZN(n686) );
  AN2D1 U181 ( .A1(n800), .A2(n857), .Z(n409) );
  CKAN2D1 U182 ( .A1(n809), .A2(n837), .Z(n424) );
  CKND0 U183 ( .I(n734), .ZN(n857) );
  OR2D0 U184 ( .A1(n476), .A2(n78), .Z(n446) );
  NR2D0 U185 ( .A1(n440), .A2(n642), .ZN(n425) );
  NR2D0 U186 ( .A1(n599), .A2(n598), .ZN(n426) );
  ND2D1 U187 ( .A1(n828), .A2(n847), .ZN(n642) );
  ND2D2 U188 ( .A1(n455), .A2(n834), .ZN(n763) );
  CKAN2D1 U189 ( .A1(n842), .A2(n509), .Z(n428) );
  CKAN2D1 U190 ( .A1(n801), .A2(n522), .Z(n429) );
  NR3D0 U191 ( .A1(n428), .A2(n429), .A3(n508), .ZN(n518) );
  INVD4 U192 ( .I(n785), .ZN(n842) );
  NR2D0 U193 ( .A1(n452), .A2(n840), .ZN(n431) );
  ND2D2 U194 ( .A1(a[6]), .A2(n839), .ZN(n785) );
  CKND0 U195 ( .I(n772), .ZN(n840) );
  CKAN2D1 U196 ( .A1(n831), .A2(n807), .Z(n434) );
  CKND1 U197 ( .I(n750), .ZN(n796) );
  CKND1 U198 ( .I(n692), .ZN(n831) );
  AN4D1 U200 ( .A1(n677), .A2(n817), .A3(n450), .A4(n845), .Z(n531) );
  ND2D0 U201 ( .A1(n677), .A2(n847), .ZN(n598) );
  ND3D1 U202 ( .A1(n816), .A2(n677), .A3(n845), .ZN(n765) );
  ND2D1 U203 ( .A1(n842), .A2(n677), .ZN(n738) );
  ND2D0 U204 ( .A1(n457), .A2(n477), .ZN(n436) );
  CKND2D0 U205 ( .A1(n826), .A2(n836), .ZN(n437) );
  OAI22D0 U206 ( .A1(n480), .A2(n716), .B1(n479), .B2(n766), .ZN(n481) );
  AOI22D0 U207 ( .A1(n838), .A2(n805), .B1(n808), .B2(n837), .ZN(n480) );
  BUFFD4 U208 ( .I(a[0]), .Z(n450) );
  AOI21D1 U209 ( .A1(n833), .A2(n842), .B(n850), .ZN(n672) );
  ND2D1 U210 ( .A1(n830), .A2(n842), .ZN(n729) );
  AOI211D0 U211 ( .A1(n818), .A2(n450), .B(n816), .C(n809), .ZN(n612) );
  ND2D0 U212 ( .A1(n455), .A2(n510), .ZN(n513) );
  CKND2D0 U213 ( .A1(n457), .A2(a[6]), .ZN(n496) );
  BUFFD4 U214 ( .I(a[2]), .Z(n451) );
  CKND2D0 U216 ( .A1(n835), .A2(n824), .ZN(n546) );
  NR2D0 U217 ( .A1(n807), .A2(n795), .ZN(n622) );
  AOI21D1 U218 ( .A1(n820), .A2(n861), .B(n848), .ZN(n577) );
  NR2D1 U219 ( .A1(n709), .A2(n750), .ZN(n741) );
  NR2XD0 U220 ( .A1(n833), .A2(n829), .ZN(n679) );
  CKND2D0 U221 ( .A1(n756), .A2(n751), .ZN(n562) );
  NR2D0 U222 ( .A1(n632), .A2(n435), .ZN(n772) );
  CKND2D0 U223 ( .A1(n688), .A2(n847), .ZN(n638) );
  NR2D0 U224 ( .A1(n809), .A2(n807), .ZN(n478) );
  OAI21D0 U225 ( .A1(n450), .A2(n692), .B(n79), .ZN(n495) );
  ND2D0 U226 ( .A1(n451), .A2(n819), .ZN(n633) );
  CKND2D1 U227 ( .A1(n778), .A2(n734), .ZN(n581) );
  NR2XD0 U228 ( .A1(n859), .A2(n522), .ZN(n523) );
  BUFFD4 U229 ( .I(a[4]), .Z(n453) );
  BUFFD4 U230 ( .I(a[3]), .Z(n452) );
  BUFFD4 U231 ( .I(a[5]), .Z(n454) );
  CKND0 U232 ( .I(n745), .ZN(n797) );
  CKND0 U233 ( .I(n779), .ZN(n859) );
  CKND0 U234 ( .I(n591), .ZN(n812) );
  OAI22D0 U235 ( .A1(n761), .A2(n758), .B1(n662), .B2(n745), .ZN(n530) );
  AOI22D0 U236 ( .A1(n860), .A2(n802), .B1(n817), .B2(n846), .ZN(n560) );
  NR2D0 U237 ( .A1(n816), .A2(n823), .ZN(n662) );
  ND2D0 U238 ( .A1(n815), .A2(n457), .ZN(n726) );
  ND2D0 U239 ( .A1(n830), .A2(n858), .ZN(n682) );
  OAI21D0 U240 ( .A1(n440), .A2(n737), .B(n789), .ZN(n483) );
  CKND2D0 U241 ( .A1(n821), .A2(n845), .ZN(n676) );
  NR2D0 U242 ( .A1(n724), .A2(n856), .ZN(n732) );
  CKND2D0 U243 ( .A1(n787), .A2(n566), .ZN(n567) );
  AOI22D0 U244 ( .A1(n808), .A2(n857), .B1(n800), .B2(n837), .ZN(n578) );
  AOI31D0 U245 ( .A1(n847), .A2(n743), .A3(n823), .B(n742), .ZN(n744) );
  NR2D0 U246 ( .A1(n860), .A2(n846), .ZN(n473) );
  CKND2D0 U247 ( .A1(n830), .A2(n459), .ZN(n680) );
  NR2XD0 U248 ( .A1(n843), .A2(n853), .ZN(n673) );
  CKND2D0 U249 ( .A1(n735), .A2(n745), .ZN(n596) );
  OAI32D0 U250 ( .A1(n569), .A2(n763), .A3(n752), .B1(n527), .B2(n526), .ZN(
        n528) );
  CKND2D0 U251 ( .A1(n769), .A2(n766), .ZN(n754) );
  NR2XD0 U252 ( .A1(n837), .A2(n847), .ZN(n646) );
  OAI21D0 U253 ( .A1(n756), .A2(n618), .B(n642), .ZN(n522) );
  OAI22D0 U254 ( .A1(n435), .A2(n761), .B1(n610), .B2(n750), .ZN(n617) );
  NR2D0 U255 ( .A1(n825), .A2(n830), .ZN(n610) );
  CKND0 U256 ( .I(n756), .ZN(n823) );
  AOI31D0 U257 ( .A1(n738), .A2(n737), .A3(n736), .B(n735), .ZN(n739) );
  CKND0 U258 ( .I(n716), .ZN(n824) );
  ND2D0 U259 ( .A1(n798), .A2(n819), .ZN(n565) );
  CKND2D0 U260 ( .A1(n796), .A2(n813), .ZN(n728) );
  CKND0 U261 ( .I(n709), .ZN(n861) );
  CKND2D0 U262 ( .A1(n831), .A2(n847), .ZN(n768) );
  AOI21D0 U263 ( .A1(n846), .A2(n816), .B(n759), .ZN(n760) );
  AOI22D0 U264 ( .A1(n807), .A2(n450), .B1(n457), .B2(n816), .ZN(n494) );
  AOI21D0 U265 ( .A1(n806), .A2(n845), .B(n580), .ZN(n524) );
  AOI21D0 U266 ( .A1(n822), .A2(n857), .B(n701), .ZN(n514) );
  CKND0 U267 ( .I(n743), .ZN(n810) );
  CKND2D0 U268 ( .A1(n816), .A2(n819), .ZN(n611) );
  NR2XD0 U269 ( .A1(n654), .A2(n772), .ZN(n613) );
  OAI33D0 U270 ( .A1(n440), .A2(n455), .A3(n774), .B1(n709), .B2(n798), .B3(
        n756), .ZN(n547) );
  AOI32D0 U272 ( .A1(n454), .A2(n456), .A3(n817), .B1(n828), .B2(n640), .ZN(
        n641) );
  OAI32D0 U273 ( .A1(n773), .A2(n485), .A3(n711), .B1(n484), .B2(n745), .ZN(
        n488) );
  NR2D0 U274 ( .A1(n856), .A2(n699), .ZN(n465) );
  OAI31D0 U275 ( .A1(n753), .A2(n781), .A3(n78), .B(n621), .ZN(n628) );
  AOI33D0 U276 ( .A1(n620), .A2(n834), .A3(n802), .B1(n853), .B2(n813), .B3(
        n797), .ZN(n621) );
  OAI22D0 U277 ( .A1(n452), .A2(n619), .B1(n456), .B2(n618), .ZN(n620) );
  AOI21D0 U278 ( .A1(n452), .A2(n858), .B(n818), .ZN(n775) );
  NR2D0 U279 ( .A1(n803), .A2(n806), .ZN(n584) );
  CKND2D0 U280 ( .A1(n725), .A2(n813), .ZN(n583) );
  OAI22D0 U281 ( .A1(n771), .A2(n74), .B1(n696), .B2(n716), .ZN(n467) );
  AOI21D0 U282 ( .A1(n70), .A2(n593), .B(n435), .ZN(n466) );
  NR2D0 U283 ( .A1(n737), .A2(n452), .ZN(n701) );
  AOI21D0 U284 ( .A1(n856), .A2(n817), .B(n701), .ZN(n704) );
  CKND2D0 U285 ( .A1(n453), .A2(n798), .ZN(n593) );
  CKND2D0 U286 ( .A1(n451), .A2(n745), .ZN(n743) );
  OAI21D0 U287 ( .A1(n715), .A2(n745), .B(n714), .ZN(n719) );
  OA33D0 U288 ( .A1(n713), .A2(n756), .A3(n435), .B1(n712), .B2(n711), .B3(
        n773), .Z(n714) );
  CKND2D1 U289 ( .A1(n604), .A2(n603), .ZN(n608) );
  CKND2D0 U290 ( .A1(n454), .A2(n834), .ZN(n521) );
  NR2D0 U291 ( .A1(n809), .A2(n452), .ZN(n625) );
  OAI33D0 U292 ( .A1(n663), .A2(n450), .A3(n798), .B1(n496), .B2(n734), .B3(
        n766), .ZN(n497) );
  CKND2D0 U293 ( .A1(n454), .A2(a[6]), .ZN(n781) );
  INVD1 U294 ( .I(n788), .ZN(n846) );
  INVD1 U295 ( .I(n712), .ZN(n808) );
  INVD1 U296 ( .I(n682), .ZN(n860) );
  INVD1 U298 ( .I(n789), .ZN(n862) );
  INVD1 U299 ( .I(n575), .ZN(n854) );
  INVD1 U300 ( .I(n566), .ZN(n803) );
  INVD1 U301 ( .I(n606), .ZN(n826) );
  INVD1 U302 ( .I(n644), .ZN(n852) );
  ND2D1 U303 ( .A1(n677), .A2(n858), .ZN(n779) );
  ND2D1 U304 ( .A1(n845), .A2(n832), .ZN(n788) );
  NR2D1 U305 ( .A1(n643), .A2(n728), .ZN(n747) );
  INVD1 U306 ( .I(n761), .ZN(n821) );
  INVD1 U307 ( .I(n598), .ZN(n856) );
  ND2D1 U308 ( .A1(n861), .A2(n824), .ZN(n789) );
  ND2D1 U309 ( .A1(n807), .A2(n456), .ZN(n712) );
  INVD1 U310 ( .I(n642), .ZN(n855) );
  INVD1 U311 ( .I(n769), .ZN(n804) );
  NR2D1 U312 ( .A1(n456), .A2(n765), .ZN(n748) );
  INVD1 U313 ( .I(n774), .ZN(n828) );
  INVD1 U314 ( .I(n638), .ZN(n849) );
  ND2D1 U315 ( .A1(n795), .A2(n825), .ZN(n606) );
  ND2D1 U316 ( .A1(n820), .A2(n836), .ZN(n708) );
  INVD1 U317 ( .I(n605), .ZN(n850) );
  INVD1 U318 ( .I(n729), .ZN(n843) );
  INVD1 U319 ( .I(n618), .ZN(n841) );
  INVD1 U320 ( .I(n565), .ZN(n820) );
  INVD1 U321 ( .I(n614), .ZN(n848) );
  OAI222D0 U322 ( .A1(n788), .A2(n591), .B1(n780), .B2(n644), .C1(n507), .C2(
        n769), .ZN(n508) );
  OAI221D0 U323 ( .A1(n623), .A2(n771), .B1(n756), .B2(n766), .C(n506), .ZN(
        n509) );
  AOI221D0 U324 ( .A1(n836), .A2(n824), .B1(n822), .B2(n581), .C(n850), .ZN(
        n507) );
  AOI221D0 U325 ( .A1(n860), .A2(n459), .B1(n843), .B2(n725), .C(n538), .ZN(
        n541) );
  AOI221D0 U326 ( .A1(n822), .A2(n858), .B1(n811), .B2(n832), .C(n539), .ZN(
        n540) );
  NR4D0 U327 ( .A1(n716), .A2(n769), .A3(n763), .A4(n827), .ZN(n742) );
  OAI32D1 U328 ( .A1(n593), .A2(n750), .A3(n692), .B1(n592), .B2(n771), .ZN(
        n594) );
  NR2D1 U329 ( .A1(n628), .A2(n627), .ZN(n629) );
  NR4D0 U330 ( .A1(n666), .A2(n665), .A3(n664), .A4(n748), .ZN(n667) );
  NR4D0 U331 ( .A1(n488), .A2(n487), .A3(n718), .A4(n486), .ZN(n489) );
  OAI221D0 U332 ( .A1(n462), .A2(n619), .B1(n780), .B2(n725), .C(n461), .ZN(
        n472) );
  OAI221D0 U333 ( .A1(n745), .A2(n74), .B1(n752), .B2(n710), .C(n690), .ZN(
        n698) );
  AOI221D0 U334 ( .A1(n80), .A2(n689), .B1(n688), .B2(n805), .C(n687), .ZN(
        n690) );
  NR4D0 U335 ( .A1(n749), .A2(n748), .A3(n747), .A4(n746), .ZN(n792) );
  INVD1 U336 ( .I(n725), .ZN(n795) );
  INVD1 U337 ( .I(n79), .ZN(n822) );
  OAI221D0 U338 ( .A1(n457), .A2(n676), .B1(n728), .B2(n682), .C(n537), .ZN(
        n554) );
  AOI22D1 U339 ( .A1(n851), .A2(n536), .B1(n699), .B2(n535), .ZN(n537) );
  NR4D0 U340 ( .A1(n719), .A2(n742), .A3(n718), .A4(n717), .ZN(n720) );
  AOI211D1 U341 ( .A1(n861), .A2(n530), .B(n529), .C(n528), .ZN(n557) );
  INR4D0 U342 ( .A1(n765), .B1(n534), .B2(n747), .B3(n717), .ZN(n556) );
  NR3D0 U343 ( .A1(n725), .A2(n819), .A3(n736), .ZN(n585) );
  NR2D1 U344 ( .A1(n633), .A2(n725), .ZN(n707) );
  AN3XD1 U345 ( .A1(n436), .A2(n437), .A3(n438), .Z(n491) );
  AN3XD1 U346 ( .A1(n446), .A2(n447), .A3(n448), .Z(n438) );
  NR4D0 U347 ( .A1(n587), .A2(n586), .A3(n585), .A4(n746), .ZN(n588) );
  NR3D0 U348 ( .A1(n521), .A2(n756), .A3(n790), .ZN(n487) );
  AOI21D1 U349 ( .A1(n860), .A2(n816), .B(n854), .ZN(n576) );
  ND2D1 U350 ( .A1(n688), .A2(n845), .ZN(n736) );
  ND2D1 U351 ( .A1(n842), .A2(n828), .ZN(n727) );
  ND2D1 U352 ( .A1(n502), .A2(n501), .ZN(n503) );
  INVD1 U353 ( .I(n752), .ZN(n829) );
  INVD1 U354 ( .I(n780), .ZN(n815) );
  ND2D1 U355 ( .A1(n458), .A2(n798), .ZN(n790) );
  NR2D1 U356 ( .A1(n713), .A2(n716), .ZN(n724) );
  INVD1 U357 ( .I(n710), .ZN(n825) );
  INVD1 U358 ( .I(n763), .ZN(n858) );
  INVD1 U359 ( .I(n735), .ZN(n806) );
  INVD1 U360 ( .I(n521), .ZN(n835) );
  ND2D1 U361 ( .A1(n829), .A2(n847), .ZN(n605) );
  AOI211XD0 U362 ( .A1(n843), .A2(n450), .B(n645), .C(n852), .ZN(n650) );
  OAI222D0 U363 ( .A1(n737), .A2(n726), .B1(n704), .B2(n456), .C1(n703), .C2(
        n778), .ZN(n705) );
  OAI222D0 U364 ( .A1(n781), .A2(n790), .B1(n780), .B2(n779), .C1(n778), .C2(
        n777), .ZN(n782) );
  OAI222D0 U365 ( .A1(n810), .A2(n638), .B1(n566), .B2(n546), .C1(n545), .C2(
        n785), .ZN(n552) );
  NR4D0 U366 ( .A1(n544), .A2(n543), .A3(n542), .A4(n602), .ZN(n545) );
  NR3D0 U367 ( .A1(n745), .A2(n452), .A3(n771), .ZN(n543) );
  NR4D0 U368 ( .A1(n516), .A2(n515), .A3(n531), .A4(n532), .ZN(n517) );
  OAI222D0 U369 ( .A1(n525), .A2(n435), .B1(n524), .B2(n756), .C1(n523), .C2(
        n769), .ZN(n529) );
  OAI222D0 U370 ( .A1(n766), .A2(n773), .B1(n787), .B2(n653), .C1(n79), .C2(
        n712), .ZN(n661) );
  AO221D0 U371 ( .A1(n800), .A2(n833), .B1(n797), .B2(n815), .C(n707), .Z(n660) );
  OAI222D0 U372 ( .A1(n451), .A2(n658), .B1(n657), .B2(n789), .C1(n656), .C2(
        n788), .ZN(n659) );
  OAI222D0 U373 ( .A1(n758), .A2(n692), .B1(n494), .B2(n771), .C1(n457), .C2(
        n756), .ZN(n505) );
  OAI222D0 U374 ( .A1(n626), .A2(n779), .B1(n625), .B2(n729), .C1(n624), .C2(
        n761), .ZN(n627) );
  OA22D0 U375 ( .A1(n781), .A2(n435), .B1(n734), .B2(n623), .Z(n624) );
  OAI222D0 U376 ( .A1(n584), .A2(n779), .B1(n788), .B2(n583), .C1(n582), .C2(
        n781), .ZN(n587) );
  OAI222D0 U377 ( .A1(n514), .A2(n750), .B1(n819), .B2(n513), .C1(n512), .C2(
        n725), .ZN(n516) );
  INR2D1 U378 ( .A1(n767), .B1(n511), .ZN(n512) );
  ND2D1 U379 ( .A1(n452), .A2(n454), .ZN(n692) );
  OAI222D0 U380 ( .A1(n712), .A2(n738), .B1(n450), .B2(n550), .C1(n790), .C2(
        n779), .ZN(n551) );
  OAI221D0 U381 ( .A1(n745), .A2(n734), .B1(n458), .B2(n788), .C(n733), .ZN(
        n740) );
  OAI221D0 U382 ( .A1(n456), .A2(n738), .B1(n711), .B2(n725), .C(n700), .ZN(
        n706) );
  AOI21D1 U383 ( .A1(n855), .A2(n457), .B(n699), .ZN(n700) );
  NR4D0 U384 ( .A1(n636), .A2(n635), .A3(n848), .A4(n634), .ZN(n637) );
  ND2D1 U385 ( .A1(n453), .A2(n452), .ZN(n756) );
  OAI221D0 U386 ( .A1(n745), .A2(n738), .B1(n711), .B2(n750), .C(n601), .ZN(
        n609) );
  NR4D0 U387 ( .A1(n450), .A2(n834), .A3(n774), .A4(n780), .ZN(n586) );
  OAI221D0 U388 ( .A1(n618), .A2(n593), .B1(n452), .B2(n779), .C(n708), .ZN(
        n539) );
  ND2D1 U389 ( .A1(n450), .A2(n451), .ZN(n766) );
  ND2D1 U390 ( .A1(n453), .A2(n813), .ZN(n716) );
  NR2D1 U391 ( .A1(n452), .A2(n454), .ZN(n688) );
  NR3D0 U392 ( .A1(n711), .A2(n827), .A3(n716), .ZN(n533) );
  ND2D1 U393 ( .A1(n454), .A2(n455), .ZN(n709) );
  ND2D1 U394 ( .A1(n451), .A2(n454), .ZN(n751) );
  NR2D1 U395 ( .A1(n765), .A2(n450), .ZN(n718) );
  AOI21D1 U396 ( .A1(n795), .A2(n655), .B(n654), .ZN(n658) );
  ND2D1 U397 ( .A1(n800), .A2(n450), .ZN(n569) );
  INVD1 U398 ( .I(n778), .ZN(n837) );
  OAI222D0 U399 ( .A1(n758), .A2(n767), .B1(n696), .B2(n727), .C1(n695), .C2(
        n785), .ZN(n697) );
  ND2D1 U400 ( .A1(n692), .A2(n78), .ZN(n694) );
  OAI222D0 U401 ( .A1(n643), .A2(n798), .B1(n618), .B2(n611), .C1(n452), .C2(
        n727), .ZN(n616) );
  INVD1 U402 ( .I(n781), .ZN(n838) );
  INVD1 U403 ( .I(n450), .ZN(n794) );
  NR4D0 U404 ( .A1(a[6]), .A2(n813), .A3(n734), .A4(n766), .ZN(n515) );
  ND2D1 U405 ( .A1(a[6]), .A2(n827), .ZN(n778) );
  INVD2 U406 ( .I(a[6]), .ZN(n834) );
  OAI222D0 U407 ( .A1(n732), .A2(n123), .B1(n730), .B2(n729), .C1(n728), .C2(
        n727), .ZN(n793) );
  OAI222D0 U408 ( .A1(n734), .A2(n606), .B1(n123), .B2(n768), .C1(n622), .C2(
        n605), .ZN(n607) );
  OAI222D0 U409 ( .A1(n123), .A2(n605), .B1(n738), .B2(n683), .C1(n643), .C2(
        n766), .ZN(n558) );
  NR3D0 U410 ( .A1(n827), .A2(n458), .A3(n731), .ZN(n542) );
  AOI21D0 U411 ( .A1(n692), .A2(n771), .B(n731), .ZN(n687) );
  AOI32D0 U412 ( .A1(n453), .A2(n839), .A3(n815), .B1(n816), .B2(n559), .ZN(
        n561) );
  ND4D1 U413 ( .A1(n80), .A2(n836), .A3(n453), .A4(n455), .ZN(n733) );
  OAI22D0 U414 ( .A1(a[6]), .A2(n453), .B1(n454), .B2(n763), .ZN(n559) );
  NR3D0 U415 ( .A1(n780), .A2(n455), .A3(n453), .ZN(n674) );
  NR3D0 U416 ( .A1(n456), .A2(n453), .A3(n692), .ZN(n602) );
  NR3D0 U417 ( .A1(n745), .A2(n453), .A3(n618), .ZN(n654) );
  ND2D1 U418 ( .A1(n453), .A2(n451), .ZN(n710) );
  ND2D1 U419 ( .A1(n452), .A2(n451), .ZN(n649) );
  OA211D0 U420 ( .A1(n565), .A2(n725), .B(n564), .C(n563), .Z(n442) );
  OA222D1 U421 ( .A1(n574), .A2(n763), .B1(n70), .B2(n573), .C1(n757), .C2(
        n572), .Z(n443) );
  NR2D0 U422 ( .A1(n799), .A2(n796), .ZN(n623) );
  AOI222D0 U423 ( .A1(n807), .A2(n824), .B1(n822), .B2(n799), .C1(n831), .C2(
        n805), .ZN(n563) );
  OAI33D0 U424 ( .A1(n758), .A2(n757), .A3(n756), .B1(n778), .B2(n798), .B3(
        n77), .ZN(n759) );
  OAI31D0 U425 ( .A1(n745), .A2(n823), .A3(n757), .B(n744), .ZN(n749) );
  OAI222D0 U426 ( .A1(n763), .A2(n633), .B1(n452), .B2(n632), .C1(n757), .C2(
        n773), .ZN(n636) );
  OAI222D0 U427 ( .A1(n457), .A2(n781), .B1(n750), .B2(n763), .C1(n757), .C2(
        n753), .ZN(n498) );
  NR2XD0 U428 ( .A1(n757), .A2(n774), .ZN(n699) );
  AOI211XD0 U429 ( .A1(n803), .A2(n823), .B(n826), .C(n702), .ZN(n703) );
  OAI31D0 U430 ( .A1(n813), .A2(n803), .A3(n809), .B(n699), .ZN(n502) );
  CKND0 U431 ( .I(n439), .ZN(n445) );
  OAI22D0 U432 ( .A1(n752), .A2(n758), .B1(n771), .B2(n790), .ZN(n693) );
  NR3D0 U433 ( .A1(n444), .A2(n800), .A3(n815), .ZN(n656) );
  INR2D0 U434 ( .A1(n533), .B1(n671), .ZN(n717) );
  OAI222D0 U435 ( .A1(n440), .A2(n729), .B1(n599), .B2(n738), .C1(n643), .C2(
        n671), .ZN(n493) );
  NR4D0 U436 ( .A1(n774), .A2(n763), .A3(n671), .A4(n452), .ZN(n746) );
  NR2D0 U437 ( .A1(n521), .A2(n671), .ZN(n580) );
  OR2D1 U438 ( .A1(n692), .A2(n526), .Z(n447) );
  OAI221D0 U439 ( .A1(n473), .A2(n780), .B1(n727), .B2(n777), .C(n575), .ZN(
        n477) );
  INVD1 U440 ( .I(n663), .ZN(n836) );
  ND2D1 U441 ( .A1(n797), .A2(n858), .ZN(n526) );
  AOI32D0 U442 ( .A1(n800), .A2(n456), .A3(n833), .B1(n797), .B2(n562), .ZN(
        n564) );
  AOI22D0 U443 ( .A1(n825), .A2(n796), .B1(n823), .B2(n451), .ZN(n582) );
  AOI31D0 U444 ( .A1(n451), .A2(n827), .A3(n80), .B(n826), .ZN(n506) );
  AOI21D0 U445 ( .A1(n737), .A2(n676), .B(n451), .ZN(n635) );
  NR3D0 U446 ( .A1(n726), .A2(n453), .A3(n839), .ZN(n665) );
  INVD1 U447 ( .I(n727), .ZN(n844) );
  OAI22D0 U448 ( .A1(n456), .A2(n727), .B1(n460), .B2(n738), .ZN(n538) );
  OAI22D1 U449 ( .A1(n460), .A2(n727), .B1(n457), .B2(n643), .ZN(n645) );
  NR4D0 U450 ( .A1(n458), .A2(n839), .A3(n769), .A4(n761), .ZN(n702) );
  MAOI22D1 U451 ( .A1(n805), .A2(n827), .B1(n619), .B2(n440), .ZN(n570) );
  AOI211D1 U452 ( .A1(n781), .A2(n663), .B(n593), .C(n435), .ZN(n486) );
  AOI21D0 U453 ( .A1(n619), .A2(n663), .B(n70), .ZN(n511) );
  OAI21D0 U454 ( .A1(n663), .A2(n79), .B(n736), .ZN(n549) );
  OAI22D0 U455 ( .A1(n834), .A2(n716), .B1(n819), .B2(n663), .ZN(n655) );
  OAI22D0 U456 ( .A1(n455), .A2(n663), .B1(n756), .B2(n734), .ZN(n463) );
  OAI31D0 U457 ( .A1(n800), .A2(n80), .A3(n811), .B(n859), .ZN(n501) );
  AOI31D0 U458 ( .A1(n453), .A2(n834), .A3(n811), .B(n701), .ZN(n484) );
  OAI22D0 U459 ( .A1(n440), .A2(n435), .B1(n750), .B2(n777), .ZN(n510) );
  OAI211D0 U460 ( .A1(n827), .A2(n761), .B(n777), .C(n756), .ZN(n689) );
  AOI22D0 U461 ( .A1(n802), .A2(n836), .B1(n811), .B2(n819), .ZN(n776) );
  AOI22D0 U462 ( .A1(n836), .A2(n754), .B1(n838), .B2(n805), .ZN(n762) );
  NR2D0 U463 ( .A1(n796), .A2(n805), .ZN(n657) );
  AOI32D0 U464 ( .A1(n455), .A2(n819), .A3(n800), .B1(n805), .B2(n463), .ZN(
        n464) );
  AOI22D0 U465 ( .A1(n829), .A2(n805), .B1(n802), .B2(n831), .ZN(n461) );
  AO221D0 U466 ( .A1(n811), .A2(n844), .B1(n851), .B2(n817), .C(n558), .Z(n449) );
  AOI21D0 U467 ( .A1(n780), .A2(n751), .B(n785), .ZN(n634) );
  NR4D0 U468 ( .A1(n692), .A2(n758), .A3(n785), .A4(n819), .ZN(n664) );
endmodule


module aes_sbox_12 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n31, n70, n192, n223, n224, n410, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869;

  AN2XD1 U28 ( .A1(n725), .A2(n724), .Z(n729) );
  OA21D1 U35 ( .A1(n709), .A2(n708), .B(n707), .Z(n714) );
  OR4D1 U199 ( .A1(n662), .A2(n582), .A3(n526), .A4(n525), .Z(n528) );
  AN2XD1 U215 ( .A1(n527), .A2(n816), .Z(n526) );
  AO31D1 U286 ( .A1(n809), .A2(n865), .A3(n687), .B(n723), .Z(n466) );
  BUFFD6 U1 ( .I(a[3]), .Z(n445) );
  BUFFD6 U2 ( .I(a[2]), .Z(n444) );
  OAI222D1 U3 ( .A1(n670), .A2(n774), .B1(n443), .B2(n564), .C1(n756), .C2(
        n563), .ZN(n565) );
  ND2D1 U4 ( .A1(n839), .A2(n845), .ZN(n632) );
  AOI221D1 U5 ( .A1(n866), .A2(n449), .B1(n858), .B2(n814), .C(n639), .ZN(n668) );
  INVD2 U6 ( .I(n649), .ZN(n823) );
  OAI221D0 U7 ( .A1(n457), .A2(n649), .B1(n778), .B2(n737), .C(n456), .ZN(n463) );
  AN2D2 U8 ( .A1(n443), .A2(n820), .Z(n677) );
  ND2D1 U9 ( .A1(n834), .A2(n840), .ZN(n661) );
  OAI31D1 U10 ( .A1(n710), .A2(n447), .A3(n433), .B(n644), .ZN(n562) );
  ND2D1 U11 ( .A1(n858), .A2(n449), .ZN(n644) );
  ND2D1 U12 ( .A1(a[6]), .A2(n845), .ZN(n786) );
  CKND2 U13 ( .I(n448), .ZN(n845) );
  INVD2 U14 ( .I(n730), .ZN(n806) );
  AOI22D2 U15 ( .A1(n837), .A2(n823), .B1(n812), .B2(n834), .ZN(n564) );
  AOI221D2 U16 ( .A1(n829), .A2(n802), .B1(n838), .B2(n814), .C(n565), .ZN(
        n566) );
  AOI221D1 U17 ( .A1(n856), .A2(n816), .B1(n698), .B2(n809), .C(n685), .ZN(
        n722) );
  AOI22D0 U18 ( .A1(n818), .A2(n839), .B1(n821), .B2(n834), .ZN(n770) );
  NR2D0 U19 ( .A1(n818), .A2(n811), .ZN(n454) );
  AOI31D0 U20 ( .A1(n446), .A2(n840), .A3(n818), .B(n700), .ZN(n478) );
  NR2D0 U21 ( .A1(n839), .A2(n818), .ZN(n521) );
  INVD2 U22 ( .I(n778), .ZN(n818) );
  OAI32D1 U23 ( .A1(n591), .A2(n750), .A3(n691), .B1(n590), .B2(n771), .ZN(
        n592) );
  NR3D2 U24 ( .A1(n434), .A2(n435), .A3(n598), .ZN(n631) );
  AOI221D2 U25 ( .A1(n443), .A2(n571), .B1(n848), .B2(n570), .C(n569), .ZN(
        n587) );
  NR2XD1 U26 ( .A1(n784), .A2(n783), .ZN(n785) );
  OAI222D1 U27 ( .A1(n448), .A2(n777), .B1(n776), .B2(n775), .C1(n786), .C2(
        n774), .ZN(n784) );
  CKBD1 U29 ( .I(n755), .Z(n31) );
  BUFFD2 U30 ( .I(n755), .Z(n70) );
  CKND2D1 U31 ( .A1(n445), .A2(n452), .ZN(n682) );
  ND2D1 U32 ( .A1(n445), .A2(n805), .ZN(n778) );
  INVD1 U33 ( .I(n758), .ZN(n807) );
  INVD1 U34 ( .I(n791), .ZN(n809) );
  INVD1 U36 ( .I(n724), .ZN(n801) );
  INVD1 U37 ( .I(n775), .ZN(n835) );
  BUFFD4 U38 ( .I(a[4]), .Z(n446) );
  ND2D0 U39 ( .A1(n445), .A2(n826), .ZN(n755) );
  ND2D2 U40 ( .A1(n432), .A2(n449), .ZN(n744) );
  ND2D1 U41 ( .A1(n445), .A2(n444), .ZN(n649) );
  ND2D1 U42 ( .A1(n432), .A2(n805), .ZN(n791) );
  INVD2 U43 ( .I(n443), .ZN(n800) );
  OAI31D1 U44 ( .A1(n677), .A2(n806), .A3(n825), .B(n676), .ZN(n678) );
  AOI21D1 U45 ( .A1(n821), .A2(n450), .B(n810), .ZN(n590) );
  INVD1 U46 ( .I(n779), .ZN(n843) );
  INVD1 U47 ( .I(a[1]), .ZN(n452) );
  OAI222D0 U48 ( .A1(n782), .A2(n791), .B1(n781), .B2(n780), .C1(n779), .C2(
        n778), .ZN(n783) );
  ND2D1 U49 ( .A1(n444), .A2(n820), .ZN(n781) );
  INVD1 U50 ( .I(n661), .ZN(n842) );
  IND2D1 U51 ( .A1(n443), .B1(n451), .ZN(n750) );
  INVD2 U52 ( .I(n445), .ZN(n820) );
  ND4D1 U53 ( .A1(n722), .A2(n721), .A3(n720), .A4(n719), .ZN(d[1]) );
  AOI221D0 U54 ( .A1(n706), .A2(n864), .B1(n823), .B2(n705), .C(n704), .ZN(
        n720) );
  AOI221D0 U55 ( .A1(n477), .A2(n451), .B1(n828), .B2(n476), .C(n475), .ZN(
        n484) );
  ND4D2 U56 ( .A1(n668), .A2(n667), .A3(n666), .A4(n665), .ZN(d[2]) );
  OAI221D0 U57 ( .A1(n744), .A2(n690), .B1(n752), .B2(n709), .C(n689), .ZN(
        n697) );
  OAI222D1 U58 ( .A1(n443), .A2(n684), .B1(n757), .B2(n683), .C1(n682), .C2(
        n681), .ZN(n685) );
  AOI211XD0 U59 ( .A1(n836), .A2(n594), .B(n592), .C(n593), .ZN(n595) );
  INVD1 U60 ( .I(n710), .ZN(n854) );
  ND2D1 U61 ( .A1(n837), .A2(n854), .ZN(n736) );
  ND2D1 U62 ( .A1(n445), .A2(n834), .ZN(n752) );
  ND2D1 U63 ( .A1(n807), .A2(n443), .ZN(n563) );
  ND2D1 U64 ( .A1(n443), .A2(n444), .ZN(n766) );
  AOI21D1 U65 ( .A1(n867), .A2(n823), .B(n861), .ZN(n573) );
  AN2XD1 U66 ( .A1(n822), .A2(n608), .Z(n427) );
  OAI222D0 U67 ( .A1(n769), .A2(n768), .B1(n767), .B2(n766), .C1(n433), .C2(
        n765), .ZN(n794) );
  OAI222D0 U68 ( .A1(n711), .A2(n737), .B1(n443), .B2(n544), .C1(n791), .C2(
        n780), .ZN(n545) );
  MAOI22D1 U69 ( .A1(n863), .A2(n820), .B1(n633), .B2(n779), .ZN(n519) );
  OAI222D0 U70 ( .A1(n789), .A2(n589), .B1(n781), .B2(n644), .C1(n501), .C2(
        n769), .ZN(n502) );
  INVD1 U71 ( .I(n711), .ZN(n815) );
  OAI222D0 U72 ( .A1(n649), .A2(n728), .B1(n597), .B2(n737), .C1(n643), .C2(
        n670), .ZN(n487) );
  INVD1 U73 ( .I(n736), .ZN(n858) );
  OAI22D1 U74 ( .A1(n474), .A2(n715), .B1(n473), .B2(n766), .ZN(n475) );
  INVD2 U75 ( .I(a[1]), .ZN(n451) );
  INVD2 U76 ( .I(n451), .ZN(n432) );
  ND2D1 U77 ( .A1(n447), .A2(n820), .ZN(n774) );
  INVD2 U78 ( .I(n444), .ZN(n805) );
  BUFFD4 U79 ( .I(n800), .Z(n449) );
  AN2D1 U80 ( .A1(n463), .A2(n449), .Z(n426) );
  ND2D1 U81 ( .A1(n443), .A2(n805), .ZN(n730) );
  CKND2D2 U82 ( .A1(n444), .A2(n452), .ZN(n670) );
  CKND2D0 U83 ( .A1(n443), .A2(n812), .ZN(n734) );
  OAI22D1 U84 ( .A1(n750), .A2(n712), .B1(n646), .B2(n744), .ZN(n647) );
  BUFFD1 U85 ( .I(n730), .Z(n440) );
  ND2D2 U86 ( .A1(n452), .A2(n805), .ZN(n758) );
  CKND2D1 U87 ( .A1(n445), .A2(n447), .ZN(n691) );
  AOI221D1 U88 ( .A1(n803), .A2(n688), .B1(n687), .B2(n812), .C(n686), .ZN(
        n689) );
  ND4D2 U89 ( .A1(n514), .A2(n513), .A3(n512), .A4(n511), .ZN(d[6]) );
  OA221D1 U90 ( .A1(n763), .A2(n192), .B1(n642), .B2(n791), .C(n223), .Z(n667)
         );
  OA221D0 U91 ( .A1(n756), .A2(n758), .B1(n715), .B2(n791), .C(n641), .Z(n192)
         );
  OA222D1 U92 ( .A1(n650), .A2(n649), .B1(n766), .B2(n768), .C1(n648), .C2(
        n778), .Z(n223) );
  INVD2 U93 ( .I(n763), .ZN(n865) );
  OR3D1 U94 ( .A1(n677), .A2(n818), .A3(n452), .Z(n640) );
  ND2D1 U95 ( .A1(n446), .A2(n445), .ZN(n756) );
  AOI22D1 U96 ( .A1(n844), .A2(n812), .B1(n815), .B2(n843), .ZN(n474) );
  CKAN2D1 U97 ( .A1(n540), .A2(n737), .Z(n473) );
  INVD2 U98 ( .I(n771), .ZN(n839) );
  ND2D2 U99 ( .A1(n448), .A2(a[6]), .ZN(n710) );
  OAI22D1 U100 ( .A1(n728), .A2(n758), .B1(n805), .B2(n735), .ZN(n669) );
  CKND2D0 U101 ( .A1(n433), .A2(n445), .ZN(n788) );
  INVD1 U102 ( .I(n451), .ZN(n433) );
  AOI221D1 U103 ( .A1(n829), .A2(n865), .B1(n818), .B2(n839), .C(n533), .ZN(
        n534) );
  AOI221D1 U104 ( .A1(n842), .A2(n831), .B1(n829), .B2(n578), .C(n857), .ZN(
        n501) );
  CKND2D1 U105 ( .A1(a[6]), .A2(n834), .ZN(n779) );
  CKND2D1 U106 ( .A1(n443), .A2(n451), .ZN(n749) );
  NR2D1 U107 ( .A1(n632), .A2(n749), .ZN(n773) );
  OA222D0 U108 ( .A1(n753), .A2(n752), .B1(n751), .B2(n750), .C1(n70), .C2(
        n749), .Z(n764) );
  OAI22D1 U109 ( .A1(n452), .A2(n638), .B1(n637), .B2(n749), .ZN(n639) );
  ND4D4 U110 ( .A1(n631), .A2(n630), .A3(n629), .A4(n628), .ZN(d[3]) );
  ND2D2 U111 ( .A1(n809), .A2(n449), .ZN(n560) );
  AOI221D1 U112 ( .A1(n819), .A2(n578), .B1(n577), .B2(n829), .C(n576), .ZN(
        n586) );
  OA21D0 U113 ( .A1(n690), .A2(n449), .B(n621), .Z(n625) );
  ND2D1 U114 ( .A1(n805), .A2(n820), .ZN(n690) );
  NR4D1 U115 ( .A1(n674), .A2(n442), .A3(n673), .A4(n861), .ZN(n684) );
  CKND2D0 U116 ( .A1(n822), .A2(n433), .ZN(n725) );
  AOI221D4 U117 ( .A1(n851), .A2(n616), .B1(n615), .B2(n449), .C(n614), .ZN(
        n629) );
  ND2D1 U118 ( .A1(n837), .A2(n848), .ZN(n728) );
  AOI221D1 U119 ( .A1(n848), .A2(n659), .B1(n851), .B2(n658), .C(n657), .ZN(
        n666) );
  OA221D1 U120 ( .A1(n752), .A2(n744), .B1(n761), .B2(n670), .C(n224), .Z(n683) );
  OA221D1 U121 ( .A1(n690), .A2(n680), .B1(n679), .B2(n791), .C(n678), .Z(n224) );
  INVD2 U122 ( .I(n752), .ZN(n836) );
  INVD2 U123 ( .I(n670), .ZN(n812) );
  OAI222D1 U124 ( .A1(n440), .A2(n540), .B1(n494), .B2(n757), .C1(n493), .C2(
        n761), .ZN(n498) );
  OAI222D1 U125 ( .A1(n575), .A2(n715), .B1(n574), .B2(n749), .C1(n432), .C2(
        n573), .ZN(n576) );
  OAI222D1 U126 ( .A1(n535), .A2(n781), .B1(n440), .B2(n632), .C1(n534), .C2(
        n724), .ZN(n547) );
  OAI222D1 U127 ( .A1(n469), .A2(n70), .B1(n691), .B2(n520), .C1(n468), .C2(
        n449), .ZN(n470) );
  AOI221D1 U128 ( .A1(n848), .A2(n503), .B1(n808), .B2(n516), .C(n502), .ZN(
        n512) );
  AOI211XD0 U129 ( .A1(n869), .A2(n815), .B(n487), .C(n669), .ZN(n514) );
  ND4D2 U130 ( .A1(n587), .A2(n588), .A3(n586), .A4(n585), .ZN(d[4]) );
  NR4D1 U131 ( .A1(n548), .A2(n547), .A3(n546), .A4(n545), .ZN(n549) );
  ND3D2 U132 ( .A1(n551), .A2(n550), .A3(n549), .ZN(d[5]) );
  AOI221D1 U133 ( .A1(n698), .A2(n750), .B1(n450), .B2(n860), .C(n562), .ZN(
        n567) );
  OAI221D1 U134 ( .A1(n672), .A2(n682), .B1(n671), .B2(n670), .C(n852), .ZN(
        n674) );
  AOI222D1 U135 ( .A1(n814), .A2(n837), .B1(n812), .B2(n489), .C1(n808), .C2(
        n439), .ZN(n494) );
  ND2D2 U136 ( .A1(n848), .A2(n835), .ZN(n726) );
  NR2D0 U137 ( .A1(n757), .A2(n775), .ZN(n698) );
  CKND2D1 U138 ( .A1(n826), .A2(n834), .ZN(n775) );
  ND2D1 U139 ( .A1(n848), .A2(n676), .ZN(n737) );
  INVD6 U140 ( .I(n446), .ZN(n826) );
  OAI32D0 U141 ( .A1(n774), .A2(n479), .A3(n710), .B1(n478), .B2(n744), .ZN(
        n482) );
  AOI221D1 U142 ( .A1(n804), .A2(n693), .B1(n439), .B2(n806), .C(n692), .ZN(
        n694) );
  AOI221D1 U143 ( .A1(n862), .A2(n801), .B1(n865), .B2(n697), .C(n696), .ZN(
        n721) );
  CKND2D1 U144 ( .A1(n448), .A2(n834), .ZN(n733) );
  INVD0 U145 ( .I(n733), .ZN(n864) );
  ND2D0 U146 ( .A1(n444), .A2(n447), .ZN(n751) );
  NR2D0 U147 ( .A1(n445), .A2(n447), .ZN(n687) );
  ND2D0 U148 ( .A1(n447), .A2(n448), .ZN(n708) );
  BUFFD6 U149 ( .I(a[5]), .Z(n447) );
  AOI221D1 U150 ( .A1(n853), .A2(n449), .B1(n863), .B2(n450), .C(n647), .ZN(
        n648) );
  AOI211XD0 U151 ( .A1(n849), .A2(n443), .B(n645), .C(n859), .ZN(n650) );
  OAI222D1 U152 ( .A1(n568), .A2(n763), .B1(n690), .B2(n567), .C1(n757), .C2(
        n566), .ZN(n569) );
  OAI222D1 U153 ( .A1(n817), .A2(n638), .B1(n560), .B2(n540), .C1(n539), .C2(
        n786), .ZN(n546) );
  NR4D1 U154 ( .A1(n538), .A2(n537), .A3(n536), .A4(n601), .ZN(n539) );
  NR2XD1 U155 ( .A1(n806), .A2(n803), .ZN(n695) );
  ND2D2 U156 ( .A1(n433), .A2(n443), .ZN(n724) );
  AOI32D0 U157 ( .A1(n447), .A2(n449), .A3(n824), .B1(n835), .B2(n640), .ZN(
        n641) );
  OAI33D0 U158 ( .A1(n661), .A2(n443), .A3(n805), .B1(n490), .B2(n733), .B3(
        n766), .ZN(n491) );
  CKND2D1 U159 ( .A1(n779), .A2(n733), .ZN(n578) );
  ND2D0 U160 ( .A1(n447), .A2(n845), .ZN(n712) );
  CKAN2D1 U161 ( .A1(n450), .A2(n471), .Z(n410) );
  CKAN2D1 U162 ( .A1(n833), .A2(n842), .Z(n424) );
  NR3D0 U163 ( .A1(n410), .A2(n424), .A3(n470), .ZN(n485) );
  CKND0 U164 ( .I(n451), .ZN(n450) );
  CKAN2D1 U165 ( .A1(n851), .A2(n464), .Z(n425) );
  NR3D0 U166 ( .A1(n425), .A2(n426), .A3(n462), .ZN(n486) );
  INVD2 U167 ( .I(n757), .ZN(n851) );
  OAI22D0 U168 ( .A1(n461), .A2(n786), .B1(n753), .B2(n642), .ZN(n462) );
  CKAN2D1 U169 ( .A1(n848), .A2(n607), .Z(n428) );
  NR3D2 U170 ( .A1(n427), .A2(n428), .A3(n606), .ZN(n630) );
  INVD2 U171 ( .I(n786), .ZN(n848) );
  CKAN2D1 U172 ( .A1(n807), .A2(n831), .Z(n429) );
  CKAN2D1 U173 ( .A1(n815), .A2(n838), .Z(n430) );
  NR3D0 U174 ( .A1(n429), .A2(n430), .A3(n772), .ZN(n787) );
  INVD1 U175 ( .I(n715), .ZN(n831) );
  ND2D1 U176 ( .A1(n448), .A2(n840), .ZN(n763) );
  BUFFD4 U177 ( .I(a[7]), .Z(n448) );
  OAI222D1 U178 ( .A1(n787), .A2(n786), .B1(n445), .B2(n846), .C1(n785), .C2(
        n449), .ZN(n793) );
  NR2D0 U179 ( .A1(n712), .A2(n715), .ZN(n723) );
  ND2D2 U180 ( .A1(n446), .A2(n820), .ZN(n715) );
  NR4D1 U181 ( .A1(n795), .A2(n793), .A3(n794), .A4(n792), .ZN(n796) );
  INVD6 U182 ( .I(n447), .ZN(n834) );
  OR2D0 U183 ( .A1(n708), .A2(a[1]), .Z(n431) );
  ND2D0 U184 ( .A1(n835), .A2(n854), .ZN(n642) );
  CKAN2D1 U185 ( .A1(n808), .A2(n856), .Z(n434) );
  CKAN2D1 U186 ( .A1(n801), .A2(n869), .Z(n435) );
  NR2D0 U187 ( .A1(n649), .A2(n642), .ZN(n436) );
  NR2D0 U188 ( .A1(n597), .A2(n596), .ZN(n437) );
  NR2D0 U189 ( .A1(n595), .A2(n763), .ZN(n438) );
  OR3D1 U190 ( .A1(n436), .A2(n437), .A3(n438), .Z(n598) );
  CKND0 U191 ( .I(n563), .ZN(n808) );
  CKND0 U192 ( .I(n790), .ZN(n869) );
  AOI22D0 U193 ( .A1(n449), .A2(n824), .B1(n820), .B2(n811), .ZN(n597) );
  NR2XD0 U194 ( .A1(n814), .A2(n801), .ZN(n621) );
  ND2D0 U195 ( .A1(n804), .A2(n865), .ZN(n520) );
  ND2D0 U196 ( .A1(n818), .A2(n860), .ZN(n572) );
  CKND2D1 U197 ( .A1(n851), .A2(n839), .ZN(n789) );
  AOI21D0 U198 ( .A1(n801), .A2(n653), .B(n652), .ZN(n656) );
  ND2D0 U200 ( .A1(n450), .A2(a[6]), .ZN(n490) );
  CKND0 U201 ( .I(n675), .ZN(n442) );
  ND3D0 U202 ( .A1(n823), .A2(n676), .A3(n851), .ZN(n765) );
  INVD1 U203 ( .I(n761), .ZN(n828) );
  NR2D0 U204 ( .A1(n643), .A2(n727), .ZN(n746) );
  NR2D0 U205 ( .A1(n823), .A2(n830), .ZN(n660) );
  NR2D0 U206 ( .A1(n806), .A2(n802), .ZN(n622) );
  NR2D0 U207 ( .A1(n816), .A2(n814), .ZN(n472) );
  AOI21D1 U208 ( .A1(n827), .A2(n868), .B(n855), .ZN(n574) );
  AOI21D1 U209 ( .A1(n439), .A2(n848), .B(n857), .ZN(n671) );
  NR2XD0 U210 ( .A1(n849), .A2(n860), .ZN(n672) );
  NR2XD0 U211 ( .A1(n439), .A2(n836), .ZN(n679) );
  CKND2D0 U212 ( .A1(n734), .A2(n744), .ZN(n594) );
  INVD1 U213 ( .I(n691), .ZN(n838) );
  CKND2D0 U214 ( .A1(n829), .A2(n854), .ZN(n613) );
  NR2D0 U216 ( .A1(n515), .A2(n670), .ZN(n577) );
  OAI22D0 U217 ( .A1(n752), .A2(n758), .B1(n771), .B2(n791), .ZN(n692) );
  ND2D0 U218 ( .A1(n444), .A2(n826), .ZN(n633) );
  CKND2D0 U219 ( .A1(n446), .A2(n444), .ZN(n709) );
  NR2XD0 U220 ( .A1(n866), .A2(n516), .ZN(n517) );
  NR2D0 U221 ( .A1(n811), .A2(n807), .ZN(n479) );
  CKND0 U222 ( .I(n780), .ZN(n866) );
  CKND0 U223 ( .I(n589), .ZN(n819) );
  OAI22D0 U224 ( .A1(n761), .A2(n758), .B1(n660), .B2(n744), .ZN(n524) );
  CKND0 U225 ( .I(n744), .ZN(n804) );
  AOI22D0 U226 ( .A1(n867), .A2(n809), .B1(n824), .B2(n853), .ZN(n554) );
  CKND2D0 U227 ( .A1(n868), .A2(n831), .ZN(n790) );
  ND2D0 U228 ( .A1(n837), .A2(n865), .ZN(n681) );
  ND2D0 U229 ( .A1(n829), .A2(n868), .ZN(n767) );
  CKND2D0 U230 ( .A1(n828), .A2(n851), .ZN(n675) );
  CKND2D0 U231 ( .A1(n841), .A2(n831), .ZN(n540) );
  NR2D0 U232 ( .A1(n723), .A2(n863), .ZN(n731) );
  CKND0 U233 ( .I(n726), .ZN(n850) );
  CKND2D0 U234 ( .A1(n806), .A2(n839), .ZN(n651) );
  AOI22D0 U235 ( .A1(n815), .A2(n864), .B1(n807), .B2(n843), .ZN(n575) );
  OAI22D0 U236 ( .A1(n449), .A2(n726), .B1(n452), .B2(n737), .ZN(n532) );
  CKND2D1 U237 ( .A1(n496), .A2(n495), .ZN(n497) );
  OAI33D0 U238 ( .A1(n761), .A2(n805), .A3(n733), .B1(n661), .B2(n433), .B3(
        n660), .ZN(n664) );
  NR2D0 U239 ( .A1(n826), .A2(n834), .ZN(n676) );
  NR2D0 U240 ( .A1(n867), .A2(n853), .ZN(n465) );
  CKND2D0 U241 ( .A1(n837), .A2(n451), .ZN(n680) );
  ND2D0 U242 ( .A1(n788), .A2(n690), .ZN(n529) );
  AOI22D0 U243 ( .A1(n858), .A2(n530), .B1(n698), .B2(n529), .ZN(n531) );
  CKND1 U244 ( .I(n669), .ZN(n852) );
  OAI32D0 U245 ( .A1(n563), .A2(n763), .A3(n752), .B1(n521), .B2(n520), .ZN(
        n522) );
  OAI31D0 U246 ( .A1(n744), .A2(n830), .A3(n757), .B(n743), .ZN(n748) );
  AOI31D0 U247 ( .A1(n854), .A2(n742), .A3(n830), .B(n741), .ZN(n743) );
  ND2D0 U248 ( .A1(n834), .A2(n845), .ZN(n617) );
  AOI32D0 U249 ( .A1(n807), .A2(n449), .A3(n439), .B1(n804), .B2(n556), .ZN(
        n558) );
  CKND2D0 U250 ( .A1(n756), .A2(n751), .ZN(n556) );
  OAI21D0 U251 ( .A1(n756), .A2(n617), .B(n642), .ZN(n516) );
  OAI22D0 U252 ( .A1(n749), .A2(n761), .B1(n609), .B2(n750), .ZN(n616) );
  NR2D0 U253 ( .A1(n832), .A2(n837), .ZN(n609) );
  OAI22D0 U254 ( .A1(n771), .A2(n781), .B1(n433), .B2(n770), .ZN(n772) );
  AOI21D0 U255 ( .A1(n618), .A2(n661), .B(n690), .ZN(n505) );
  AOI31D0 U256 ( .A1(n737), .A2(n736), .A3(n735), .B(n734), .ZN(n738) );
  AOI22D0 U257 ( .A1(n842), .A2(n754), .B1(n844), .B2(n812), .ZN(n762) );
  CKND2D0 U258 ( .A1(n769), .A2(n766), .ZN(n754) );
  INR2D0 U259 ( .A1(n527), .B1(n670), .ZN(n716) );
  ND2D0 U260 ( .A1(n676), .A2(n854), .ZN(n596) );
  CKND2D0 U261 ( .A1(n802), .A2(n820), .ZN(n727) );
  CKND0 U262 ( .I(n708), .ZN(n868) );
  CKND2D0 U263 ( .A1(n788), .A2(n560), .ZN(n561) );
  CKND0 U264 ( .I(n617), .ZN(n847) );
  AOI211XD0 U265 ( .A1(n847), .A2(n815), .B(n492), .C(n491), .ZN(n493) );
  CKND2D1 U266 ( .A1(n603), .A2(n602), .ZN(n607) );
  AOI21D0 U267 ( .A1(n813), .A2(n851), .B(n577), .ZN(n518) );
  AOI21D0 U268 ( .A1(n829), .A2(n864), .B(n700), .ZN(n508) );
  ND2D0 U269 ( .A1(n448), .A2(n504), .ZN(n507) );
  OAI21D0 U270 ( .A1(n661), .A2(n70), .B(n735), .ZN(n543) );
  OAI33D0 U271 ( .A1(n649), .A2(n448), .A3(n775), .B1(n708), .B2(n805), .B3(
        n756), .ZN(n541) );
  CKND0 U272 ( .I(n742), .ZN(n817) );
  ND2D0 U273 ( .A1(n823), .A2(n826), .ZN(n610) );
  AOI21D0 U274 ( .A1(n863), .A2(n824), .B(n700), .ZN(n703) );
  CKND2D0 U275 ( .A1(n691), .A2(n70), .ZN(n693) );
  NR2D0 U276 ( .A1(n863), .A2(n698), .ZN(n457) );
  AOI32D0 U277 ( .A1(n448), .A2(n826), .A3(n807), .B1(n812), .B2(n455), .ZN(
        n456) );
  OAI22D0 U278 ( .A1(n448), .A2(n661), .B1(n756), .B2(n733), .ZN(n455) );
  OAI21D0 U279 ( .A1(n649), .A2(n736), .B(n790), .ZN(n477) );
  AOI21D0 U280 ( .A1(n862), .A2(n450), .B(n698), .ZN(n699) );
  ND4D0 U281 ( .A1(n803), .A2(n842), .A3(n446), .A4(n448), .ZN(n732) );
  OAI21D0 U282 ( .A1(n757), .A2(n618), .B(n726), .ZN(n599) );
  OAI211D0 U283 ( .A1(n559), .A2(n724), .B(n558), .C(n557), .ZN(n570) );
  OAI22D0 U284 ( .A1(n791), .A2(n790), .B1(n789), .B2(n788), .ZN(n792) );
  AOI211D0 U285 ( .A1(n782), .A2(n661), .B(n591), .C(n749), .ZN(n480) );
  OAI31D0 U287 ( .A1(n753), .A2(n782), .A3(n70), .B(n620), .ZN(n627) );
  AOI33D0 U288 ( .A1(n619), .A2(n840), .A3(n809), .B1(n860), .B2(n820), .B3(
        n804), .ZN(n620) );
  OAI22D0 U289 ( .A1(n445), .A2(n618), .B1(n449), .B2(n617), .ZN(n619) );
  AOI21D0 U290 ( .A1(n445), .A2(n865), .B(n825), .ZN(n776) );
  CKND2D0 U291 ( .A1(n724), .A2(n820), .ZN(n580) );
  NR2D0 U292 ( .A1(n736), .A2(n445), .ZN(n700) );
  AOI21D0 U293 ( .A1(n781), .A2(n751), .B(n786), .ZN(n634) );
  AOI21D0 U294 ( .A1(n690), .A2(n591), .B(n749), .ZN(n458) );
  CKND0 U295 ( .I(n644), .ZN(n859) );
  OAI22D0 U296 ( .A1(n452), .A2(n726), .B1(n432), .B2(n643), .ZN(n645) );
  ND2D0 U297 ( .A1(n446), .A2(n805), .ZN(n591) );
  OAI21D0 U298 ( .A1(n714), .A2(n744), .B(n713), .ZN(n718) );
  CKND2D1 U299 ( .A1(n447), .A2(n826), .ZN(n771) );
  OAI211D0 U300 ( .A1(n447), .A2(n788), .B(n633), .C(n70), .ZN(n542) );
  ND2D1 U301 ( .A1(n840), .A2(n845), .ZN(n757) );
  CKND2D0 U302 ( .A1(n444), .A2(n744), .ZN(n742) );
  AOI21D0 U303 ( .A1(n853), .A2(n823), .B(n759), .ZN(n760) );
  OAI33D0 U304 ( .A1(n758), .A2(n757), .A3(n756), .B1(n779), .B2(n805), .B3(
        n31), .ZN(n759) );
  CKND2D0 U305 ( .A1(n447), .A2(n840), .ZN(n515) );
  NR2D0 U306 ( .A1(n802), .A2(n812), .ZN(n655) );
  NR2D0 U307 ( .A1(n446), .A2(n840), .ZN(n467) );
  NR2XD0 U308 ( .A1(n652), .A2(n773), .ZN(n612) );
  NR2D0 U309 ( .A1(n816), .A2(n445), .ZN(n624) );
  CKND2D0 U310 ( .A1(n447), .A2(a[6]), .ZN(n782) );
  AOI32D0 U311 ( .A1(n446), .A2(n845), .A3(n822), .B1(n823), .B2(n553), .ZN(
        n555) );
  INVD1 U312 ( .I(n789), .ZN(n853) );
  INVD1 U313 ( .I(n681), .ZN(n867) );
  INVD1 U314 ( .I(n605), .ZN(n833) );
  INVD1 U315 ( .I(n572), .ZN(n861) );
  AOI222D0 U316 ( .A1(n814), .A2(n831), .B1(n829), .B2(n806), .C1(n838), .C2(
        n812), .ZN(n557) );
  ND2D1 U317 ( .A1(n676), .A2(n865), .ZN(n780) );
  INVD1 U318 ( .I(n596), .ZN(n863) );
  AO221D0 U319 ( .A1(n807), .A2(n439), .B1(n804), .B2(n822), .C(n706), .Z(n658) );
  INVD1 U320 ( .I(n750), .ZN(n802) );
  INVD1 U321 ( .I(n643), .ZN(n860) );
  INVD1 U322 ( .I(n769), .ZN(n811) );
  INVD1 U323 ( .I(n642), .ZN(n862) );
  INVD1 U324 ( .I(n560), .ZN(n810) );
  INVD1 U325 ( .I(n638), .ZN(n856) );
  ND2D1 U326 ( .A1(n818), .A2(n450), .ZN(n589) );
  INVD1 U327 ( .I(n728), .ZN(n849) );
  INVD1 U328 ( .I(n690), .ZN(n821) );
  INVD1 U329 ( .I(n604), .ZN(n857) );
  ND2D1 U330 ( .A1(n801), .A2(n832), .ZN(n605) );
  ND2D1 U331 ( .A1(n827), .A2(n842), .ZN(n707) );
  INVD1 U332 ( .I(n559), .ZN(n827) );
  INVD1 U333 ( .I(n613), .ZN(n855) );
  OAI221D0 U334 ( .A1(n454), .A2(n618), .B1(n781), .B2(n724), .C(n453), .ZN(
        n464) );
  OAI222D0 U335 ( .A1(n766), .A2(n774), .B1(n788), .B2(n651), .C1(n70), .C2(
        n711), .ZN(n659) );
  AOI221D0 U336 ( .A1(n867), .A2(n451), .B1(n849), .B2(n724), .C(n532), .ZN(
        n535) );
  NR4D0 U337 ( .A1(n718), .A2(n741), .A3(n717), .A4(n716), .ZN(n719) );
  OAI222D0 U338 ( .A1(n751), .A2(n724), .B1(n775), .B2(n589), .C1(n756), .C2(
        n766), .ZN(n593) );
  IND4D1 U339 ( .A1(n799), .B1(n798), .B2(n797), .B3(n796), .ZN(d[0]) );
  AOI221D0 U340 ( .A1(n740), .A2(n822), .B1(n821), .B2(n739), .C(n738), .ZN(
        n798) );
  NR4D0 U341 ( .A1(n748), .A2(n747), .A3(n746), .A4(n745), .ZN(n797) );
  OAI221D0 U342 ( .A1(n465), .A2(n781), .B1(n726), .B2(n778), .C(n572), .ZN(
        n471) );
  INVD1 U343 ( .I(n70), .ZN(n829) );
  ND4D1 U344 ( .A1(n484), .A2(n486), .A3(n485), .A4(n483), .ZN(d[7]) );
  NR4D0 U345 ( .A1(n482), .A2(n481), .A3(n717), .A4(n480), .ZN(n483) );
  NR4D0 U346 ( .A1(n584), .A2(n583), .A3(n582), .A4(n745), .ZN(n585) );
  AOI221D0 U347 ( .A1(n818), .A2(n850), .B1(n858), .B2(n824), .C(n552), .ZN(
        n588) );
  NR4D0 U348 ( .A1(n664), .A2(n663), .A3(n662), .A4(n747), .ZN(n665) );
  NR2D1 U349 ( .A1(n843), .A2(n854), .ZN(n646) );
  NR2D1 U350 ( .A1(n627), .A2(n626), .ZN(n628) );
  AOI211D1 U351 ( .A1(n868), .A2(n524), .B(n523), .C(n522), .ZN(n551) );
  INR4D0 U352 ( .A1(n765), .B1(n528), .B2(n746), .B3(n716), .ZN(n550) );
  OAI221D0 U353 ( .A1(n432), .A2(n675), .B1(n727), .B2(n681), .C(n531), .ZN(
        n548) );
  ND2D1 U354 ( .A1(n449), .A2(n805), .ZN(n769) );
  NR3D0 U355 ( .A1(n724), .A2(n826), .A3(n735), .ZN(n582) );
  ND2D1 U356 ( .A1(n854), .A2(n839), .ZN(n643) );
  ND2D1 U357 ( .A1(n687), .A2(n851), .ZN(n735) );
  INVD1 U358 ( .I(n781), .ZN(n822) );
  NR3D0 U359 ( .A1(n515), .A2(n756), .A3(n791), .ZN(n481) );
  INVD1 U360 ( .I(n788), .ZN(n824) );
  NR2D1 U361 ( .A1(n443), .A2(n431), .ZN(n740) );
  INVD1 U362 ( .I(n749), .ZN(n803) );
  ND2D1 U363 ( .A1(n687), .A2(n854), .ZN(n638) );
  INVD1 U364 ( .I(n756), .ZN(n830) );
  NR2D1 U365 ( .A1(n633), .A2(n724), .ZN(n706) );
  NR2D1 U366 ( .A1(n449), .A2(n765), .ZN(n747) );
  INVD1 U367 ( .I(n753), .ZN(n814) );
  ND2D1 U368 ( .A1(n814), .A2(n449), .ZN(n711) );
  INVD1 U369 ( .I(n682), .ZN(n825) );
  ND2D1 U370 ( .A1(n820), .A2(n826), .ZN(n761) );
  ND2D1 U371 ( .A1(n838), .A2(n854), .ZN(n768) );
  ND2D1 U372 ( .A1(n805), .A2(n826), .ZN(n559) );
  INVD1 U373 ( .I(n734), .ZN(n813) );
  INVD1 U374 ( .I(n515), .ZN(n841) );
  AOI221D0 U375 ( .A1(n810), .A2(n439), .B1(n835), .B2(n561), .C(n706), .ZN(
        n568) );
  INVD1 U376 ( .I(n709), .ZN(n832) );
  INVD1 U377 ( .I(n618), .ZN(n837) );
  OAI222D0 U378 ( .A1(n444), .A2(n656), .B1(n655), .B2(n790), .C1(n654), .C2(
        n789), .ZN(n657) );
  OAI222D0 U379 ( .A1(n758), .A2(n691), .B1(n488), .B2(n771), .C1(n432), .C2(
        n756), .ZN(n499) );
  OAI222D0 U380 ( .A1(n581), .A2(n780), .B1(n789), .B2(n580), .C1(n579), .C2(
        n782), .ZN(n584) );
  OA221D0 U381 ( .A1(n758), .A2(n733), .B1(n766), .B2(n779), .C(n441), .Z(n469) );
  OAI221D0 U382 ( .A1(n622), .A2(n771), .B1(n756), .B2(n766), .C(n500), .ZN(
        n503) );
  OAI222D0 U383 ( .A1(n758), .A2(n767), .B1(n695), .B2(n726), .C1(n694), .C2(
        n786), .ZN(n696) );
  OAI222D0 U384 ( .A1(n758), .A2(n613), .B1(n612), .B2(n805), .C1(n611), .C2(
        n681), .ZN(n614) );
  OAI222D0 U385 ( .A1(n643), .A2(n805), .B1(n617), .B2(n610), .C1(n445), .C2(
        n726), .ZN(n615) );
  OAI222D0 U386 ( .A1(n736), .A2(n725), .B1(n703), .B2(n449), .C1(n702), .C2(
        n779), .ZN(n704) );
  NR4D0 U387 ( .A1(n432), .A2(n845), .A3(n769), .A4(n761), .ZN(n701) );
  OAI222D0 U388 ( .A1(n432), .A2(n782), .B1(n750), .B2(n763), .C1(n757), .C2(
        n753), .ZN(n492) );
  OAI222D0 U389 ( .A1(n519), .A2(n749), .B1(n518), .B2(n756), .C1(n517), .C2(
        n769), .ZN(n523) );
  ND2D1 U390 ( .A1(n432), .A2(n444), .ZN(n753) );
  OAI211D1 U391 ( .A1(n708), .A2(n682), .B(n555), .C(n554), .ZN(n571) );
  INVD1 U392 ( .I(n773), .ZN(n846) );
  NR3D0 U393 ( .A1(n744), .A2(n445), .A3(n771), .ZN(n537) );
  OAI222D0 U394 ( .A1(n479), .A2(n712), .B1(n472), .B2(n710), .C1(n733), .C2(
        n734), .ZN(n476) );
  NR4D0 U395 ( .A1(n775), .A2(n763), .A3(n670), .A4(n445), .ZN(n745) );
  NR4D0 U396 ( .A1(n691), .A2(n758), .A3(n786), .A4(n826), .ZN(n662) );
  NR4D0 U397 ( .A1(n510), .A2(n509), .A3(n525), .A4(n526), .ZN(n511) );
  AOI211XD0 U398 ( .A1(n865), .A2(n499), .B(n498), .C(n497), .ZN(n513) );
  NR4D0 U399 ( .A1(n460), .A2(n459), .A3(n536), .A4(n458), .ZN(n461) );
  OAI222D0 U400 ( .A1(n752), .A2(n560), .B1(n649), .B2(n724), .C1(n753), .C2(
        n691), .ZN(n460) );
  AOI221D0 U401 ( .A1(n812), .A2(n543), .B1(n851), .B2(n542), .C(n541), .ZN(
        n544) );
  OAI222D0 U402 ( .A1(n764), .A2(n763), .B1(n762), .B2(n761), .C1(n443), .C2(
        n760), .ZN(n795) );
  NR3D0 U403 ( .A1(n744), .A2(n446), .A3(n617), .ZN(n652) );
  OAI221D0 U404 ( .A1(n744), .A2(n733), .B1(n450), .B2(n789), .C(n732), .ZN(
        n739) );
  OAI221D0 U405 ( .A1(n617), .A2(n591), .B1(n445), .B2(n780), .C(n707), .ZN(
        n533) );
  NR4D0 U406 ( .A1(n636), .A2(n635), .A3(n855), .A4(n634), .ZN(n637) );
  OAI222D0 U407 ( .A1(n763), .A2(n633), .B1(n445), .B2(n632), .C1(n757), .C2(
        n774), .ZN(n636) );
  NR3D0 U408 ( .A1(n449), .A2(n446), .A3(n691), .ZN(n601) );
  AOI222D0 U409 ( .A1(n809), .A2(n828), .B1(n830), .B2(n811), .C1(n813), .C2(
        n447), .ZN(n603) );
  NR3D0 U410 ( .A1(n781), .A2(n448), .A3(n446), .ZN(n673) );
  NR3D0 U411 ( .A1(n725), .A2(n446), .A3(n845), .ZN(n663) );
  OAI221D0 U412 ( .A1(n744), .A2(n737), .B1(n710), .B2(n750), .C(n600), .ZN(
        n608) );
  AOI221D0 U413 ( .A1(n841), .A2(n801), .B1(n599), .B2(n451), .C(n740), .ZN(
        n600) );
  OAI222D0 U414 ( .A1(n625), .A2(n780), .B1(n624), .B2(n728), .C1(n623), .C2(
        n761), .ZN(n626) );
  OA22D0 U415 ( .A1(n782), .A2(n749), .B1(n733), .B2(n622), .Z(n623) );
  ND2D1 U416 ( .A1(n446), .A2(n834), .ZN(n618) );
  OAI222D0 U417 ( .A1(n508), .A2(n750), .B1(n826), .B2(n507), .C1(n506), .C2(
        n724), .ZN(n510) );
  INR2D1 U418 ( .A1(n767), .B1(n505), .ZN(n506) );
  INVD1 U419 ( .I(n782), .ZN(n844) );
  CKBD4 U420 ( .I(a[0]), .Z(n443) );
  AOI221D0 U421 ( .A1(n801), .A2(n821), .B1(n808), .B2(n836), .C(n601), .ZN(
        n602) );
  ND2D1 U422 ( .A1(n836), .A2(n854), .ZN(n604) );
  AOI22D0 U423 ( .A1(n836), .A2(n812), .B1(n809), .B2(n838), .ZN(n453) );
  INVD1 U424 ( .I(n774), .ZN(n439) );
  OAI31D0 U425 ( .A1(n807), .A2(n803), .A3(n818), .B(n866), .ZN(n495) );
  OAI22D0 U426 ( .A1(n649), .A2(n749), .B1(n750), .B2(n778), .ZN(n504) );
  OAI211D0 U427 ( .A1(n834), .A2(n761), .B(n778), .C(n756), .ZN(n688) );
  AOI22D0 U428 ( .A1(n809), .A2(n842), .B1(n818), .B2(n826), .ZN(n777) );
  OAI221D0 U429 ( .A1(n449), .A2(n737), .B1(n710), .B2(n724), .C(n699), .ZN(
        n705) );
  AOI211XD0 U430 ( .A1(n810), .A2(n830), .B(n833), .C(n701), .ZN(n702) );
  NR3D0 U431 ( .A1(n677), .A2(n807), .A3(n822), .ZN(n654) );
  AOI21D1 U432 ( .A1(n803), .A2(n841), .B(n740), .ZN(n441) );
  INVD1 U433 ( .I(n766), .ZN(n816) );
  NR2D1 U434 ( .A1(n810), .A2(n813), .ZN(n581) );
  OAI31D0 U435 ( .A1(n820), .A2(n810), .A3(n816), .B(n698), .ZN(n496) );
  AOI22D0 U436 ( .A1(n832), .A2(n802), .B1(n830), .B2(n444), .ZN(n579) );
  AOI31D0 U437 ( .A1(n444), .A2(n834), .A3(n803), .B(n833), .ZN(n500) );
  AOI21D0 U438 ( .A1(n736), .A2(n675), .B(n444), .ZN(n635) );
  NR4D0 U439 ( .A1(n715), .A2(n769), .A3(n763), .A4(n834), .ZN(n741) );
  OAI22D0 U440 ( .A1(n840), .A2(n715), .B1(n826), .B2(n661), .ZN(n653) );
  OAI22D0 U441 ( .A1(n771), .A2(n690), .B1(n695), .B2(n715), .ZN(n459) );
  OAI222D0 U442 ( .A1(n731), .A2(n440), .B1(n729), .B2(n728), .C1(n727), .C2(
        n726), .ZN(n799) );
  AOI21D0 U443 ( .A1(n691), .A2(n771), .B(n440), .ZN(n686) );
  OAI222D0 U444 ( .A1(n733), .A2(n605), .B1(n440), .B2(n768), .C1(n621), .C2(
        n604), .ZN(n606) );
  OAI222D0 U445 ( .A1(n440), .A2(n604), .B1(n737), .B2(n682), .C1(n643), .C2(
        n766), .ZN(n552) );
  OAI222D0 U446 ( .A1(n440), .A2(n70), .B1(n695), .B2(n691), .C1(n761), .C2(
        n560), .ZN(n538) );
  CKND2D0 U447 ( .A1(n440), .A2(n758), .ZN(n530) );
  NR3D0 U448 ( .A1(n834), .A2(n433), .A3(n440), .ZN(n536) );
  NR4D0 U449 ( .A1(n443), .A2(n840), .A3(n775), .A4(n781), .ZN(n583) );
  NR2D1 U450 ( .A1(n765), .A2(n443), .ZN(n717) );
  AOI22D0 U451 ( .A1(n814), .A2(n443), .B1(n450), .B2(n823), .ZN(n488) );
  AN4D1 U452 ( .A1(n676), .A2(n824), .A3(n443), .A4(n851), .Z(n525) );
  AOI211D1 U453 ( .A1(n825), .A2(n443), .B(n823), .C(n816), .ZN(n611) );
  OAI21D0 U454 ( .A1(n443), .A2(n691), .B(n70), .ZN(n489) );
  AOI221D1 U455 ( .A1(n467), .A2(n814), .B1(n858), .B2(n824), .C(n466), .ZN(
        n468) );
  INVD2 U456 ( .I(a[6]), .ZN(n840) );
  NR4D0 U457 ( .A1(a[6]), .A2(n820), .A3(n733), .A4(n766), .ZN(n509) );
  OA33D0 U458 ( .A1(n712), .A2(n756), .A3(n749), .B1(n711), .B2(n710), .B3(
        n774), .Z(n713) );
  NR3D0 U459 ( .A1(n710), .A2(n834), .A3(n715), .ZN(n527) );
  OAI22D0 U460 ( .A1(a[6]), .A2(n446), .B1(n447), .B2(n763), .ZN(n553) );
endmodule


module aes_sbox_11 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n70, n187, n192, n287, n310, n314, n404, n405, n408, n409, n410, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863;

  OA21D1 U35 ( .A1(n702), .A2(n701), .B(n700), .Z(n707) );
  OR4D1 U199 ( .A1(n656), .A2(n575), .A3(n521), .A4(n520), .Z(n523) );
  AN2XD1 U215 ( .A1(n522), .A2(n809), .Z(n521) );
  AN2XD1 U271 ( .A1(n535), .A2(n730), .Z(n468) );
  INVD2 U1 ( .I(n751), .ZN(n800) );
  ND4D3 U2 ( .A1(n192), .A2(n580), .A3(n579), .A4(n578), .ZN(d[4]) );
  ND2D1 U3 ( .A1(n450), .A2(n437), .ZN(n746) );
  AOI32D0 U4 ( .A1(n446), .A2(n819), .A3(n800), .B1(n805), .B2(n454), .ZN(n455) );
  INVD2 U5 ( .I(n446), .ZN(n839) );
  AOI21D1 U6 ( .A1(n847), .A2(n816), .B(n752), .ZN(n753) );
  OAI221D1 U7 ( .A1(n666), .A2(n676), .B1(n665), .B2(n664), .C(n846), .ZN(n668) );
  OAI222D1 U8 ( .A1(n446), .A2(n770), .B1(n769), .B2(n768), .C1(n779), .C2(
        n767), .ZN(n777) );
  INVD4 U9 ( .I(n664), .ZN(n805) );
  OAI22D0 U10 ( .A1(n429), .A2(n705), .B1(n638), .B2(n737), .ZN(n639) );
  AOI221D1 U11 ( .A1(n822), .A2(n859), .B1(n811), .B2(n832), .C(n528), .ZN(
        n529) );
  CKND2D1 U12 ( .A1(n813), .A2(n819), .ZN(n754) );
  CKND6 U13 ( .I(n444), .ZN(n819) );
  CKND2D2 U14 ( .A1(n842), .A2(n828), .ZN(n719) );
  INVD3 U15 ( .I(n779), .ZN(n842) );
  AOI221D1 U16 ( .A1(n835), .A2(n794), .B1(n591), .B2(n448), .C(n733), .ZN(
        n592) );
  CKND2D2 U17 ( .A1(n450), .A2(n442), .ZN(n717) );
  CKAN2D1 U18 ( .A1(n718), .A2(n717), .Z(n722) );
  OAI221D1 U19 ( .A1(n614), .A2(n764), .B1(n749), .B2(n759), .C(n495), .ZN(
        n498) );
  CKND2 U20 ( .I(n663), .ZN(n846) );
  OAI22D2 U21 ( .A1(n721), .A2(n751), .B1(n798), .B2(n728), .ZN(n663) );
  OAI21D2 U22 ( .A1(n750), .A2(n610), .B(n719), .ZN(n591) );
  NR2D1 U23 ( .A1(n705), .A2(n708), .ZN(n716) );
  AOI221D1 U24 ( .A1(n861), .A2(n448), .B1(n843), .B2(n717), .C(n527), .ZN(
        n530) );
  OAI221D1 U25 ( .A1(n737), .A2(n730), .B1(n703), .B2(n429), .C(n592), .ZN(
        n600) );
  INVD3 U26 ( .I(n448), .ZN(n450) );
  BUFFD6 U27 ( .I(a[4]), .Z(n444) );
  INVD1 U28 ( .I(n768), .ZN(n828) );
  ND2D1 U29 ( .A1(a[6]), .A2(n839), .ZN(n779) );
  BUFFD4 U30 ( .I(a[7]), .Z(n446) );
  ND2D3 U31 ( .A1(a[2]), .A2(n451), .ZN(n664) );
  BUFFD6 U32 ( .I(a[0]), .Z(n442) );
  INVD1 U33 ( .I(n784), .ZN(n802) );
  CKND2D1 U34 ( .A1(n443), .A2(n819), .ZN(n748) );
  ND2D0 U36 ( .A1(n793), .A2(n798), .ZN(n762) );
  CKND2D2 U37 ( .A1(n442), .A2(n448), .ZN(n742) );
  INVD1 U38 ( .I(n771), .ZN(n811) );
  AOI221D2 U39 ( .A1(n442), .A2(n564), .B1(n842), .B2(n563), .C(n562), .ZN(
        n580) );
  IND4D1 U40 ( .A1(n792), .B1(n791), .B2(n790), .B3(n789), .ZN(d[0]) );
  INVD1 U41 ( .I(n708), .ZN(n824) );
  INVD1 U42 ( .I(n655), .ZN(n836) );
  OAI221D0 U43 ( .A1(n609), .A2(n583), .B1(n443), .B2(n773), .C(n700), .ZN(
        n528) );
  ND2D1 U44 ( .A1(n827), .A2(n834), .ZN(n655) );
  INVD1 U45 ( .I(n767), .ZN(n833) );
  INVD1 U46 ( .I(n742), .ZN(n796) );
  INVD1 U47 ( .I(n772), .ZN(n837) );
  AOI211D1 U48 ( .A1(n803), .A2(n823), .B(n826), .C(n694), .ZN(n695) );
  AOI221D1 U49 ( .A1(n859), .A2(n644), .B1(n856), .B2(n802), .C(n643), .ZN(
        n661) );
  OAI221D0 U50 ( .A1(n749), .A2(n751), .B1(n708), .B2(n432), .C(n633), .ZN(
        n644) );
  INVD1 U51 ( .I(n704), .ZN(n808) );
  INVD1 U52 ( .I(n717), .ZN(n794) );
  ND3D1 U53 ( .A1(n546), .A2(n545), .A3(n544), .ZN(d[5]) );
  AOI221D0 U54 ( .A1(n811), .A2(n844), .B1(n852), .B2(n817), .C(n547), .ZN(
        n192) );
  AN2XD1 U55 ( .A1(n781), .A2(n555), .Z(n431) );
  NR2D1 U56 ( .A1(n561), .A2(n756), .ZN(n405) );
  NR2D1 U57 ( .A1(n750), .A2(n559), .ZN(n409) );
  INVD2 U58 ( .I(n442), .ZN(n793) );
  ND2D2 U59 ( .A1(n442), .A2(n798), .ZN(n723) );
  ND2D1 U60 ( .A1(n798), .A2(n813), .ZN(n683) );
  ND2D1 U61 ( .A1(n450), .A2(n793), .ZN(n737) );
  AN3XD1 U62 ( .A1(n622), .A2(n620), .A3(n621), .Z(n70) );
  INVD2 U63 ( .I(a[2]), .ZN(n798) );
  AOI221D1 U64 ( .A1(n860), .A2(n793), .B1(n852), .B2(n807), .C(n631), .ZN(
        n662) );
  AOI21D1 U65 ( .A1(n684), .A2(n764), .B(n723), .ZN(n679) );
  AOI221D1 U66 ( .A1(n699), .A2(n858), .B1(n816), .B2(n698), .C(n697), .ZN(
        n713) );
  OAI22D1 U67 ( .A1(n764), .A2(n774), .B1(n449), .B2(n763), .ZN(n765) );
  ND2D2 U68 ( .A1(n451), .A2(n798), .ZN(n751) );
  INVD1 U69 ( .I(n782), .ZN(n847) );
  AOI221D1 U70 ( .A1(n815), .A2(n600), .B1(n842), .B2(n599), .C(n598), .ZN(
        n622) );
  OAI222D0 U71 ( .A1(n726), .A2(n597), .B1(n723), .B2(n761), .C1(n613), .C2(
        n596), .ZN(n598) );
  AOI211XD0 U72 ( .A1(n863), .A2(n808), .B(n482), .C(n663), .ZN(n509) );
  AOI221D1 U73 ( .A1(n797), .A2(n686), .B1(n833), .B2(n433), .C(n685), .ZN(
        n687) );
  OAI222D0 U74 ( .A1(n751), .A2(n760), .B1(n688), .B2(n719), .C1(n687), .C2(
        n779), .ZN(n689) );
  INVD1 U75 ( .I(n691), .ZN(n287) );
  AOI221D1 U76 ( .A1(n691), .A2(n429), .B1(n449), .B2(n854), .C(n556), .ZN(
        n560) );
  AOI21D1 U77 ( .A1(n856), .A2(n449), .B(n691), .ZN(n692) );
  NR2XD0 U78 ( .A1(n750), .A2(n768), .ZN(n691) );
  ND4D2 U79 ( .A1(n661), .A2(n662), .A3(n660), .A4(n659), .ZN(d[2]) );
  OAI31D1 U80 ( .A1(n818), .A2(n799), .A3(n671), .B(n670), .ZN(n672) );
  OA221D1 U81 ( .A1(n683), .A2(n674), .B1(n673), .B2(n432), .C(n672), .Z(n441)
         );
  ND2D2 U82 ( .A1(n830), .A2(n848), .ZN(n729) );
  INVD2 U83 ( .I(n610), .ZN(n830) );
  ND2D1 U84 ( .A1(n450), .A2(n798), .ZN(n784) );
  AOI31D1 U85 ( .A1(n802), .A2(n859), .A3(n680), .B(n716), .ZN(n439) );
  AOI22D1 U86 ( .A1(n811), .A2(n832), .B1(n814), .B2(n827), .ZN(n763) );
  OA221D1 U87 ( .A1(n751), .A2(n726), .B1(n759), .B2(n772), .C(n187), .Z(n466)
         );
  AOI21D1 U88 ( .A1(n796), .A2(n835), .B(n733), .ZN(n187) );
  AOI211XD1 U89 ( .A1(n859), .A2(n494), .B(n493), .C(n492), .ZN(n508) );
  OAI222D1 U90 ( .A1(n723), .A2(n535), .B1(n489), .B2(n750), .C1(n488), .C2(
        n754), .ZN(n493) );
  OAI222D1 U91 ( .A1(n568), .A2(n708), .B1(n567), .B2(n742), .C1(n449), .C2(
        n566), .ZN(n569) );
  OAI222D1 U92 ( .A1(n641), .A2(n634), .B1(n589), .B2(n588), .C1(n587), .C2(
        n756), .ZN(n590) );
  AOI221D1 U93 ( .A1(n845), .A2(n463), .B1(n462), .B2(n793), .C(n461), .ZN(
        n481) );
  OAI221D0 U94 ( .A1(n456), .A2(n641), .B1(n771), .B2(n730), .C(n455), .ZN(
        n462) );
  ND4D3 U95 ( .A1(n481), .A2(n480), .A3(n479), .A4(n478), .ZN(d[7]) );
  OA221D1 U96 ( .A1(n745), .A2(n737), .B1(n754), .B2(n664), .C(n441), .Z(n677)
         );
  OA221D1 U97 ( .A1(n630), .A2(n759), .B1(n287), .B2(n784), .C(n310), .Z(n715)
         );
  AN3XD1 U98 ( .A1(n410), .A2(n424), .A3(n425), .Z(n310) );
  OA221D1 U99 ( .A1(n748), .A2(n429), .B1(n684), .B2(n746), .C(n440), .Z(n559)
         );
  ND2D1 U100 ( .A1(n852), .A2(n793), .ZN(n636) );
  INVD2 U101 ( .I(n729), .ZN(n852) );
  NR2D1 U102 ( .A1(n560), .A2(n683), .ZN(n408) );
  CKND2D1 U103 ( .A1(n446), .A2(n827), .ZN(n726) );
  ND2D0 U104 ( .A1(n772), .A2(n726), .ZN(n571) );
  OAI22D0 U105 ( .A1(n446), .A2(n655), .B1(n749), .B2(n726), .ZN(n454) );
  INVD1 U106 ( .I(n726), .ZN(n858) );
  AOI211XD0 U107 ( .A1(n841), .A2(n808), .B(n487), .C(n486), .ZN(n488) );
  OAI31D1 U108 ( .A1(n703), .A2(n445), .A3(n450), .B(n636), .ZN(n556) );
  AOI221D1 U109 ( .A1(n801), .A2(n850), .B1(n794), .B2(n863), .C(n590), .ZN(
        n623) );
  NR4D1 U110 ( .A1(n543), .A2(n542), .A3(n541), .A4(n540), .ZN(n544) );
  OAI222D1 U111 ( .A1(n530), .A2(n774), .B1(n723), .B2(n624), .C1(n529), .C2(
        n717), .ZN(n542) );
  ND2D2 U112 ( .A1(n800), .A2(n442), .ZN(n557) );
  OAI222D1 U113 ( .A1(n642), .A2(n641), .B1(n759), .B2(n761), .C1(n640), .C2(
        n771), .ZN(n643) );
  AOI221D1 U114 ( .A1(n472), .A2(n448), .B1(n821), .B2(n471), .C(n470), .ZN(
        n479) );
  INVD3 U115 ( .I(n641), .ZN(n816) );
  ND2D2 U116 ( .A1(n443), .A2(a[2]), .ZN(n641) );
  AOI22D1 U117 ( .A1(n830), .A2(n816), .B1(n805), .B2(n827), .ZN(n558) );
  AOI221D1 U118 ( .A1(n847), .A2(n793), .B1(n857), .B2(n450), .C(n639), .ZN(
        n640) );
  CKND2D1 U119 ( .A1(n445), .A2(n834), .ZN(n510) );
  CKND2D1 U120 ( .A1(n445), .A2(n446), .ZN(n701) );
  CKND2D2 U121 ( .A1(n819), .A2(n827), .ZN(n768) );
  CKND2D2 U122 ( .A1(n445), .A2(n819), .ZN(n764) );
  CKND2D1 U123 ( .A1(n443), .A2(n445), .ZN(n684) );
  NR2XD0 U124 ( .A1(n819), .A2(n827), .ZN(n670) );
  CKND2D2 U125 ( .A1(n443), .A2(n827), .ZN(n745) );
  ND2D2 U126 ( .A1(n444), .A2(n827), .ZN(n610) );
  INVD6 U127 ( .I(n445), .ZN(n827) );
  NR4D1 U128 ( .A1(n788), .A2(n787), .A3(n786), .A4(n785), .ZN(n789) );
  AOI221D1 U129 ( .A1(n800), .A2(n824), .B1(n808), .B2(n831), .C(n765), .ZN(
        n780) );
  INVD6 U130 ( .I(n443), .ZN(n813) );
  BUFFD8 U131 ( .I(a[3]), .Z(n443) );
  OAI222D1 U132 ( .A1(n780), .A2(n779), .B1(n443), .B2(n840), .C1(n778), .C2(
        n793), .ZN(n786) );
  ND2D1 U133 ( .A1(n443), .A2(n451), .ZN(n676) );
  AN2XD1 U134 ( .A1(n442), .A2(n813), .Z(n671) );
  ND2D4 U135 ( .A1(n442), .A2(a[2]), .ZN(n759) );
  CKND2D1 U136 ( .A1(a[6]), .A2(n827), .ZN(n772) );
  OA221D1 U137 ( .A1(n448), .A2(n314), .B1(n597), .B2(n655), .C(n404), .Z(n480) );
  OA221D0 U138 ( .A1(n464), .A2(n774), .B1(n719), .B2(n771), .C(n565), .Z(n314) );
  OA222D0 U139 ( .A1(n466), .A2(n748), .B1(n684), .B2(n515), .C1(n465), .C2(
        n793), .Z(n404) );
  ND2D1 U140 ( .A1(n830), .A2(n842), .ZN(n721) );
  ND4D2 U141 ( .A1(n715), .A2(n714), .A3(n713), .A4(n712), .ZN(d[1]) );
  INVD2 U142 ( .I(n447), .ZN(n451) );
  AOI221D1 U143 ( .A1(n856), .A2(n794), .B1(n859), .B2(n690), .C(n689), .ZN(
        n714) );
  ND2D3 U144 ( .A1(n446), .A2(a[6]), .ZN(n703) );
  ND2D2 U145 ( .A1(n834), .A2(n839), .ZN(n750) );
  ND2D2 U146 ( .A1(n446), .A2(n834), .ZN(n756) );
  OR2D0 U147 ( .A1(n444), .A2(n834), .Z(n438) );
  INVD4 U148 ( .I(a[6]), .ZN(n834) );
  OR3D1 U149 ( .A1(n405), .A2(n408), .A3(n409), .Z(n562) );
  OA221D0 U150 ( .A1(n555), .A2(n767), .B1(n768), .B2(n431), .C(n430), .Z(n561) );
  OR2XD1 U151 ( .A1(n678), .A2(n442), .Z(n410) );
  OR2D0 U152 ( .A1(n677), .A2(n750), .Z(n424) );
  OR2D0 U153 ( .A1(n435), .A2(n675), .Z(n425) );
  ND2D1 U154 ( .A1(n830), .A2(n859), .ZN(n675) );
  CKAN2D1 U155 ( .A1(n842), .A2(n498), .Z(n426) );
  CKAN2D1 U156 ( .A1(n801), .A2(n511), .Z(n427) );
  NR3D0 U157 ( .A1(n426), .A2(n427), .A3(n497), .ZN(n507) );
  INVD1 U158 ( .I(n557), .ZN(n801) );
  OAI21D0 U159 ( .A1(n749), .A2(n609), .B(n634), .ZN(n511) );
  ND4D2 U160 ( .A1(n509), .A2(n508), .A3(n507), .A4(n506), .ZN(d[6]) );
  INR4D1 U161 ( .A1(n669), .B1(n855), .B2(n667), .B3(n668), .ZN(n678) );
  ND2D2 U162 ( .A1(n444), .A2(n813), .ZN(n708) );
  NR2D1 U163 ( .A1(n624), .A2(n742), .ZN(n766) );
  INVD2 U164 ( .I(n764), .ZN(n832) );
  OAI22D0 U165 ( .A1(n745), .A2(n751), .B1(n764), .B2(n432), .ZN(n685) );
  OAI32D0 U166 ( .A1(n583), .A2(n429), .A3(n684), .B1(n582), .B2(n764), .ZN(
        n584) );
  ND2D0 U167 ( .A1(n793), .A2(n448), .ZN(n743) );
  ND2D2 U168 ( .A1(n802), .A2(n793), .ZN(n555) );
  ND2D1 U169 ( .A1(n807), .A2(n793), .ZN(n704) );
  BUFFD6 U170 ( .I(a[5]), .Z(n445) );
  INVD1 U171 ( .I(n743), .ZN(n428) );
  CKND3 U172 ( .I(n428), .ZN(n429) );
  INVD4 U173 ( .I(a[1]), .ZN(n448) );
  CKND1 U174 ( .I(n699), .ZN(n430) );
  INVD2 U175 ( .I(n555), .ZN(n803) );
  ND2D0 U176 ( .A1(n450), .A2(n798), .ZN(n432) );
  CKND2D2 U177 ( .A1(n623), .A2(n70), .ZN(d[3]) );
  CKND0 U178 ( .I(n448), .ZN(n449) );
  ND2D0 U179 ( .A1(n829), .A2(n848), .ZN(n596) );
  CKND1 U180 ( .I(n774), .ZN(n815) );
  AOI221D1 U181 ( .A1(n812), .A2(n571), .B1(n570), .B2(n822), .C(n569), .ZN(
        n579) );
  CKND0 U182 ( .I(n581), .ZN(n812) );
  NR2D0 U183 ( .A1(n807), .A2(n794), .ZN(n613) );
  NR2D0 U184 ( .A1(n837), .A2(n848), .ZN(n638) );
  CKND2D0 U185 ( .A1(n828), .A2(n848), .ZN(n634) );
  ND2D0 U186 ( .A1(n832), .A2(n839), .ZN(n624) );
  CKND2D0 U187 ( .A1(n831), .A2(n848), .ZN(n761) );
  CKND2D0 U188 ( .A1(n822), .A2(n848), .ZN(n605) );
  OAI211D1 U189 ( .A1(n701), .A2(n435), .B(n550), .C(n549), .ZN(n564) );
  ND2D0 U190 ( .A1(n445), .A2(n839), .ZN(n705) );
  NR2D0 U191 ( .A1(n758), .A2(n442), .ZN(n710) );
  ND2D0 U192 ( .A1(n445), .A2(a[6]), .ZN(n775) );
  CKND0 U193 ( .I(n773), .ZN(n860) );
  ND2D0 U194 ( .A1(n845), .A2(n832), .ZN(n782) );
  AOI22D0 U195 ( .A1(n861), .A2(n802), .B1(n817), .B2(n847), .ZN(n549) );
  NR2D0 U196 ( .A1(n804), .A2(n800), .ZN(n474) );
  CKND2D0 U197 ( .A1(n862), .A2(n824), .ZN(n783) );
  CKND2D0 U198 ( .A1(n811), .A2(n854), .ZN(n565) );
  ND2D0 U200 ( .A1(n822), .A2(n862), .ZN(n760) );
  CKND2D0 U201 ( .A1(n821), .A2(n845), .ZN(n669) );
  ND2D0 U202 ( .A1(n835), .A2(n824), .ZN(n535) );
  ND2D0 U203 ( .A1(n797), .A2(n859), .ZN(n515) );
  NR2D0 U204 ( .A1(n716), .A2(n857), .ZN(n724) );
  CKND0 U205 ( .I(n719), .ZN(n844) );
  NR2D0 U206 ( .A1(n825), .A2(n830), .ZN(n601) );
  OAI31D0 U207 ( .A1(n737), .A2(n823), .A3(n750), .B(n736), .ZN(n741) );
  AOI31D0 U208 ( .A1(n848), .A2(n735), .A3(n823), .B(n734), .ZN(n736) );
  OAI22D0 U209 ( .A1(n754), .A2(n751), .B1(n654), .B2(n737), .ZN(n519) );
  CKND2D0 U210 ( .A1(n781), .A2(n683), .ZN(n524) );
  CKND2D0 U211 ( .A1(n723), .A2(n751), .ZN(n525) );
  OAI31D0 U212 ( .A1(n800), .A2(n796), .A3(n811), .B(n860), .ZN(n490) );
  ND2D0 U213 ( .A1(n827), .A2(n839), .ZN(n609) );
  AOI32D0 U214 ( .A1(n800), .A2(n793), .A3(n833), .B1(n797), .B2(n551), .ZN(
        n553) );
  CKND2D0 U216 ( .A1(n749), .A2(n744), .ZN(n551) );
  AOI21D0 U217 ( .A1(n610), .A2(n655), .B(n683), .ZN(n500) );
  NR2D0 U218 ( .A1(n816), .A2(n823), .ZN(n654) );
  CKND2D0 U219 ( .A1(n815), .A2(n449), .ZN(n718) );
  AOI22D0 U220 ( .A1(n808), .A2(n858), .B1(n800), .B2(n837), .ZN(n568) );
  CKND2D0 U221 ( .A1(n795), .A2(n813), .ZN(n720) );
  CKND0 U222 ( .I(n701), .ZN(n862) );
  MAOI22D0 U223 ( .A1(n857), .A2(n813), .B1(n625), .B2(n772), .ZN(n514) );
  AOI21D0 U224 ( .A1(n806), .A2(n845), .B(n570), .ZN(n513) );
  AOI22D0 U225 ( .A1(n802), .A2(n836), .B1(n811), .B2(n819), .ZN(n770) );
  AOI22D0 U226 ( .A1(n807), .A2(n442), .B1(n449), .B2(n816), .ZN(n483) );
  NR2XD0 U227 ( .A1(n777), .A2(n776), .ZN(n778) );
  NR2D0 U228 ( .A1(n809), .A2(n807), .ZN(n467) );
  CKND0 U229 ( .I(n609), .ZN(n841) );
  CKND0 U230 ( .I(n735), .ZN(n810) );
  CKND2D0 U231 ( .A1(n816), .A2(n819), .ZN(n602) );
  NR2XD0 U232 ( .A1(n646), .A2(n766), .ZN(n604) );
  AOI211D0 U233 ( .A1(n818), .A2(n442), .B(n816), .C(n809), .ZN(n603) );
  OAI33D0 U234 ( .A1(n754), .A2(n798), .A3(n726), .B1(n655), .B2(n449), .B3(
        n654), .ZN(n658) );
  AOI21D0 U235 ( .A1(n833), .A2(n842), .B(n851), .ZN(n665) );
  NR2D0 U236 ( .A1(n861), .A2(n847), .ZN(n464) );
  NR2D0 U237 ( .A1(n857), .A2(n691), .ZN(n456) );
  INVD2 U238 ( .I(n703), .ZN(n848) );
  OAI22D0 U239 ( .A1(n764), .A2(n683), .B1(n688), .B2(n708), .ZN(n458) );
  AOI21D0 U240 ( .A1(n683), .A2(n583), .B(n742), .ZN(n457) );
  ND2D0 U241 ( .A1(n450), .A2(n443), .ZN(n781) );
  AOI211D0 U242 ( .A1(n775), .A2(n655), .B(n583), .C(n742), .ZN(n475) );
  CKND0 U243 ( .I(n636), .ZN(n853) );
  AOI211XD0 U244 ( .A1(n843), .A2(n442), .B(n637), .C(n853), .ZN(n642) );
  NR2D0 U245 ( .A1(n803), .A2(n806), .ZN(n574) );
  CKND2D0 U246 ( .A1(n717), .A2(n813), .ZN(n573) );
  OAI22D0 U247 ( .A1(n834), .A2(n708), .B1(n819), .B2(n655), .ZN(n647) );
  OAI22D0 U248 ( .A1(n451), .A2(n630), .B1(n629), .B2(n742), .ZN(n631) );
  AOI22D0 U249 ( .A1(n838), .A2(n805), .B1(n808), .B2(n837), .ZN(n469) );
  OAI22D0 U250 ( .A1(n469), .A2(n708), .B1(n468), .B2(n759), .ZN(n470) );
  CKND2D0 U251 ( .A1(n727), .A2(n737), .ZN(n586) );
  NR2D0 U252 ( .A1(n625), .A2(n717), .ZN(n699) );
  OAI32D0 U253 ( .A1(n767), .A2(n474), .A3(n703), .B1(n473), .B2(n737), .ZN(
        n477) );
  OAI21D0 U254 ( .A1(n707), .A2(n737), .B(n706), .ZN(n711) );
  AOI22D0 U255 ( .A1(n836), .A2(n747), .B1(n838), .B2(n805), .ZN(n755) );
  CKND2D0 U256 ( .A1(n762), .A2(n759), .ZN(n747) );
  NR2D0 U257 ( .A1(n811), .A2(n804), .ZN(n453) );
  AOI22D0 U258 ( .A1(n829), .A2(n805), .B1(n802), .B2(n831), .ZN(n452) );
  CKND2D1 U259 ( .A1(n595), .A2(n594), .ZN(n599) );
  CKND2D0 U260 ( .A1(n798), .A2(n819), .ZN(n554) );
  AOI21D0 U261 ( .A1(n794), .A2(n647), .B(n646), .ZN(n650) );
  NR2D0 U262 ( .A1(n795), .A2(n805), .ZN(n649) );
  OAI33D0 U263 ( .A1(n655), .A2(n442), .A3(n798), .B1(n485), .B2(n726), .B3(
        n759), .ZN(n486) );
  ND2D0 U264 ( .A1(n450), .A2(a[6]), .ZN(n485) );
  AOI32D0 U265 ( .A1(n444), .A2(n839), .A3(n815), .B1(n816), .B2(n548), .ZN(
        n550) );
  INVD1 U266 ( .I(n448), .ZN(n447) );
  INVD1 U267 ( .I(n675), .ZN(n861) );
  INVD1 U268 ( .I(n783), .ZN(n863) );
  INVD1 U269 ( .I(n597), .ZN(n826) );
  INVD1 U270 ( .I(n565), .ZN(n855) );
  INVD1 U272 ( .I(n630), .ZN(n850) );
  INVD1 U273 ( .I(n588), .ZN(n857) );
  INVD1 U274 ( .I(n634), .ZN(n856) );
  ND2D1 U275 ( .A1(n794), .A2(n825), .ZN(n597) );
  INVD1 U276 ( .I(n635), .ZN(n854) );
  ND2D1 U277 ( .A1(n811), .A2(n450), .ZN(n581) );
  INVD1 U278 ( .I(n596), .ZN(n851) );
  ND2D1 U279 ( .A1(n820), .A2(n836), .ZN(n700) );
  INVD1 U280 ( .I(n721), .ZN(n843) );
  INVD1 U281 ( .I(n605), .ZN(n849) );
  AOI221D0 U282 ( .A1(n796), .A2(n681), .B1(n680), .B2(n805), .C(n679), .ZN(
        n682) );
  OAI221D0 U283 ( .A1(n449), .A2(n669), .B1(n720), .B2(n675), .C(n526), .ZN(
        n543) );
  AOI21D1 U284 ( .A1(n820), .A2(n862), .B(n849), .ZN(n567) );
  AOI21D1 U285 ( .A1(n861), .A2(n816), .B(n855), .ZN(n566) );
  OAI222D0 U286 ( .A1(n723), .A2(n748), .B1(n688), .B2(n684), .C1(n754), .C2(
        n555), .ZN(n533) );
  AOI21D1 U287 ( .A1(n814), .A2(n450), .B(n803), .ZN(n582) );
  NR4D0 U288 ( .A1(n708), .A2(n762), .A3(n756), .A4(n827), .ZN(n734) );
  ND2D1 U289 ( .A1(n491), .A2(n490), .ZN(n492) );
  NR4D0 U290 ( .A1(n741), .A2(n740), .A3(n739), .A4(n738), .ZN(n790) );
  AOI221D0 U291 ( .A1(n733), .A2(n815), .B1(n814), .B2(n732), .C(n731), .ZN(
        n791) );
  OAI222D0 U292 ( .A1(n724), .A2(n723), .B1(n722), .B2(n721), .C1(n720), .C2(
        n719), .ZN(n792) );
  NR4D0 U293 ( .A1(n658), .A2(n657), .A3(n656), .A4(n740), .ZN(n659) );
  NR2D1 U294 ( .A1(n619), .A2(n618), .ZN(n620) );
  AOI221D0 U295 ( .A1(n845), .A2(n608), .B1(n607), .B2(n793), .C(n606), .ZN(
        n621) );
  NR2D1 U296 ( .A1(n701), .A2(n429), .ZN(n733) );
  NR4D0 U297 ( .A1(n477), .A2(n476), .A3(n710), .A4(n475), .ZN(n478) );
  INR4D0 U298 ( .A1(n758), .B1(n523), .B2(n739), .B3(n709), .ZN(n545) );
  AOI211D1 U299 ( .A1(n862), .A2(n519), .B(n518), .C(n517), .ZN(n546) );
  NR4D0 U300 ( .A1(n711), .A2(n734), .A3(n710), .A4(n709), .ZN(n712) );
  ND2D1 U301 ( .A1(n680), .A2(n845), .ZN(n728) );
  NR3D0 U302 ( .A1(n717), .A2(n819), .A3(n728), .ZN(n575) );
  NR4D0 U303 ( .A1(n577), .A2(n576), .A3(n575), .A4(n738), .ZN(n578) );
  INVD1 U304 ( .I(n746), .ZN(n807) );
  INVD1 U305 ( .I(n683), .ZN(n814) );
  ND2D1 U306 ( .A1(n848), .A2(n832), .ZN(n635) );
  INVD1 U307 ( .I(n702), .ZN(n825) );
  INVD1 U308 ( .I(n762), .ZN(n804) );
  INVD1 U309 ( .I(n510), .ZN(n835) );
  INVD1 U310 ( .I(n756), .ZN(n859) );
  INVD1 U311 ( .I(n745), .ZN(n829) );
  INVD1 U312 ( .I(n727), .ZN(n806) );
  INVD1 U313 ( .I(n676), .ZN(n818) );
  INVD1 U314 ( .I(n554), .ZN(n820) );
  INVD1 U315 ( .I(n750), .ZN(n845) );
  INVD1 U316 ( .I(n723), .ZN(n799) );
  NR2D1 U317 ( .A1(n860), .A2(n511), .ZN(n512) );
  OA22D0 U318 ( .A1(n775), .A2(n742), .B1(n726), .B2(n614), .Z(n615) );
  INVD1 U319 ( .I(n766), .ZN(n840) );
  OAI222D0 U320 ( .A1(n729), .A2(n718), .B1(n696), .B2(n793), .C1(n695), .C2(
        n772), .ZN(n697) );
  NR4D0 U321 ( .A1(n450), .A2(n839), .A3(n762), .A4(n754), .ZN(n694) );
  OAI222D0 U322 ( .A1(n704), .A2(n730), .B1(n442), .B2(n539), .C1(n432), .C2(
        n773), .ZN(n540) );
  AOI221D0 U323 ( .A1(n794), .A2(n814), .B1(n801), .B2(n829), .C(n593), .ZN(
        n594) );
  AOI222D0 U324 ( .A1(n802), .A2(n821), .B1(n823), .B2(n804), .C1(n806), .C2(
        n445), .ZN(n595) );
  OAI222D0 U325 ( .A1(n574), .A2(n773), .B1(n782), .B2(n573), .C1(n572), .C2(
        n775), .ZN(n577) );
  OAI222D0 U326 ( .A1(n450), .A2(n775), .B1(n429), .B2(n756), .C1(n750), .C2(
        n746), .ZN(n487) );
  OAI222D0 U327 ( .A1(n474), .A2(n705), .B1(n467), .B2(n703), .C1(n726), .C2(
        n727), .ZN(n471) );
  OAI222D0 U328 ( .A1(n775), .A2(n432), .B1(n774), .B2(n773), .C1(n772), .C2(
        n771), .ZN(n776) );
  NR2XD0 U329 ( .A1(n843), .A2(n854), .ZN(n666) );
  OAI222D0 U330 ( .A1(n751), .A2(n605), .B1(n604), .B2(n798), .C1(n603), .C2(
        n675), .ZN(n606) );
  AOI211XD0 U331 ( .A1(n829), .A2(n586), .B(n585), .C(n584), .ZN(n587) );
  OAI211D1 U332 ( .A1(n554), .A2(n717), .B(n553), .C(n552), .ZN(n563) );
  OAI221D0 U333 ( .A1(n737), .A2(n726), .B1(n450), .B2(n782), .C(n725), .ZN(
        n732) );
  OAI222D0 U334 ( .A1(n782), .A2(n581), .B1(n774), .B2(n636), .C1(n496), .C2(
        n762), .ZN(n497) );
  AOI221D0 U335 ( .A1(n836), .A2(n824), .B1(n822), .B2(n571), .C(n851), .ZN(
        n496) );
  NR4D0 U336 ( .A1(n505), .A2(n504), .A3(n520), .A4(n521), .ZN(n506) );
  INVD1 U337 ( .I(n759), .ZN(n809) );
  OAI222D0 U338 ( .A1(n762), .A2(n761), .B1(n760), .B2(n759), .C1(n449), .C2(
        n758), .ZN(n787) );
  OAI222D0 U339 ( .A1(n757), .A2(n756), .B1(n755), .B2(n754), .C1(n442), .C2(
        n753), .ZN(n788) );
  OAI221D0 U340 ( .A1(n453), .A2(n610), .B1(n774), .B2(n717), .C(n452), .ZN(
        n463) );
  NR3D0 U341 ( .A1(n737), .A2(n444), .A3(n609), .ZN(n646) );
  NR4D0 U342 ( .A1(n442), .A2(n834), .A3(n768), .A4(n774), .ZN(n576) );
  OAI222D0 U343 ( .A1(n810), .A2(n630), .B1(n555), .B2(n535), .C1(n534), .C2(
        n779), .ZN(n541) );
  NR4D0 U344 ( .A1(n533), .A2(n532), .A3(n531), .A4(n593), .ZN(n534) );
  NR4D0 U345 ( .A1(n459), .A2(n458), .A3(n531), .A4(n457), .ZN(n460) );
  ND2D1 U346 ( .A1(n444), .A2(n443), .ZN(n749) );
  NR4D0 U347 ( .A1(n628), .A2(n627), .A3(n849), .A4(n626), .ZN(n629) );
  ND2D1 U348 ( .A1(n443), .A2(n798), .ZN(n771) );
  NR3D0 U349 ( .A1(n703), .A2(n827), .A3(n708), .ZN(n522) );
  NR3D0 U350 ( .A1(n718), .A2(n444), .A3(n839), .ZN(n657) );
  OAI222D0 U351 ( .A1(n751), .A2(n684), .B1(n483), .B2(n764), .C1(n449), .C2(
        n749), .ZN(n494) );
  ND2D1 U352 ( .A1(n442), .A2(n805), .ZN(n727) );
  ND2D1 U353 ( .A1(n445), .A2(n813), .ZN(n767) );
  ND2D1 U354 ( .A1(n444), .A2(n798), .ZN(n583) );
  OA221D0 U355 ( .A1(n438), .A2(n746), .B1(n729), .B2(n781), .C(n439), .Z(n465) );
  INVD1 U356 ( .I(n775), .ZN(n838) );
  OAI222D0 U357 ( .A1(n744), .A2(n717), .B1(n768), .B2(n581), .C1(n749), .C2(
        n759), .ZN(n585) );
  OAI222D0 U358 ( .A1(n503), .A2(n429), .B1(n819), .B2(n502), .C1(n501), .C2(
        n717), .ZN(n505) );
  ND2D1 U359 ( .A1(n446), .A2(n499), .ZN(n502) );
  INR2D1 U360 ( .A1(n760), .B1(n500), .ZN(n501) );
  OAI222D0 U361 ( .A1(n759), .A2(n767), .B1(n781), .B2(n645), .C1(n748), .C2(
        n704), .ZN(n653) );
  OAI222D0 U362 ( .A1(n635), .A2(n798), .B1(n609), .B2(n602), .C1(n443), .C2(
        n719), .ZN(n607) );
  CKND0 U363 ( .I(n723), .ZN(n433) );
  CKBD0 U364 ( .I(n745), .Z(n434) );
  NR2D0 U365 ( .A1(n443), .A2(n445), .ZN(n680) );
  AOI21D0 U366 ( .A1(n443), .A2(n859), .B(n818), .ZN(n769) );
  OAI222D0 U367 ( .A1(n756), .A2(n625), .B1(n443), .B2(n624), .C1(n750), .C2(
        n767), .ZN(n628) );
  NR2D0 U368 ( .A1(n729), .A2(n443), .ZN(n693) );
  NR3D0 U369 ( .A1(n737), .A2(n443), .A3(n764), .ZN(n532) );
  NR2D0 U370 ( .A1(n809), .A2(n443), .ZN(n616) );
  OAI211D0 U371 ( .A1(n827), .A2(n754), .B(n771), .C(n749), .ZN(n681) );
  AOI33D0 U372 ( .A1(n611), .A2(n834), .A3(n802), .B1(n854), .B2(n813), .B3(
        n797), .ZN(n612) );
  NR4D0 U373 ( .A1(a[6]), .A2(n813), .A3(n726), .A4(n759), .ZN(n504) );
  OAI31D1 U374 ( .A1(n813), .A2(n803), .A3(n809), .B(n691), .ZN(n491) );
  CKND2D1 U375 ( .A1(a[2]), .A2(n813), .ZN(n774) );
  OAI33D0 U376 ( .A1(n641), .A2(n446), .A3(n768), .B1(n701), .B2(n798), .B3(
        n749), .ZN(n536) );
  ND2D1 U377 ( .A1(n684), .A2(n748), .ZN(n686) );
  OAI31D1 U378 ( .A1(n746), .A2(n775), .A3(n748), .B(n612), .ZN(n619) );
  OAI21D1 U379 ( .A1(n655), .A2(n748), .B(n728), .ZN(n538) );
  OAI21D0 U380 ( .A1(n442), .A2(n684), .B(n748), .ZN(n484) );
  OAI33D0 U381 ( .A1(n751), .A2(n750), .A3(n749), .B1(n772), .B2(n798), .B3(
        n748), .ZN(n752) );
  INVD1 U382 ( .I(n749), .ZN(n823) );
  OA33D0 U383 ( .A1(n705), .A2(n749), .A3(n742), .B1(n704), .B2(n703), .B3(
        n767), .Z(n706) );
  OAI222D0 U384 ( .A1(n514), .A2(n742), .B1(n513), .B2(n749), .C1(n512), .C2(
        n762), .ZN(n518) );
  NR3D0 U385 ( .A1(n510), .A2(n749), .A3(n432), .ZN(n476) );
  ND2D1 U386 ( .A1(n680), .A2(n848), .ZN(n630) );
  OAI22D0 U387 ( .A1(n432), .A2(n783), .B1(n782), .B2(n781), .ZN(n785) );
  AOI21D1 U388 ( .A1(n857), .A2(n817), .B(n693), .ZN(n696) );
  AOI21D1 U389 ( .A1(n822), .A2(n858), .B(n693), .ZN(n503) );
  AOI31D1 U390 ( .A1(n444), .A2(n834), .A3(n811), .B(n693), .ZN(n473) );
  OAI222D0 U391 ( .A1(n617), .A2(n773), .B1(n616), .B2(n721), .C1(n615), .C2(
        n754), .ZN(n618) );
  AOI221D0 U392 ( .A1(n805), .A2(n538), .B1(n845), .B2(n537), .C(n536), .ZN(
        n539) );
  ND2D0 U393 ( .A1(a[2]), .A2(n819), .ZN(n625) );
  AOI222D0 U394 ( .A1(n807), .A2(n824), .B1(n822), .B2(n433), .C1(n831), .C2(
        n805), .ZN(n552) );
  NR2D0 U395 ( .A1(n799), .A2(n795), .ZN(n614) );
  NR2XD0 U396 ( .A1(n433), .A2(n796), .ZN(n688) );
  CKND2D0 U397 ( .A1(n433), .A2(n832), .ZN(n645) );
  ND4D1 U398 ( .A1(n796), .A2(n836), .A3(n444), .A4(n446), .ZN(n725) );
  OAI221D0 U399 ( .A1(n793), .A2(n730), .B1(n703), .B2(n717), .C(n692), .ZN(
        n698) );
  NR3D0 U400 ( .A1(n774), .A2(n446), .A3(n444), .ZN(n667) );
  CKBD0 U401 ( .I(n676), .Z(n435) );
  CKND0 U402 ( .I(a[2]), .ZN(n436) );
  INVD1 U403 ( .I(n436), .ZN(n437) );
  INVD1 U404 ( .I(n781), .ZN(n817) );
  OA222D1 U405 ( .A1(n664), .A2(n767), .B1(n442), .B2(n558), .C1(n749), .C2(
        n557), .Z(n440) );
  INVD1 U406 ( .I(n748), .ZN(n822) );
  CKND1 U407 ( .I(n429), .ZN(n795) );
  INVD1 U408 ( .I(n684), .ZN(n831) );
  NR2D0 U409 ( .A1(n510), .A2(n664), .ZN(n570) );
  CKND2D0 U410 ( .A1(n830), .A2(n448), .ZN(n674) );
  AOI222D0 U411 ( .A1(n807), .A2(n830), .B1(n805), .B2(n484), .C1(n801), .C2(
        n833), .ZN(n489) );
  OR3D0 U412 ( .A1(n671), .A2(n811), .A3(n451), .Z(n632) );
  AN4D1 U413 ( .A1(n670), .A2(n817), .A3(n442), .A4(n845), .Z(n520) );
  ND2D1 U414 ( .A1(n670), .A2(n859), .ZN(n773) );
  ND3D0 U415 ( .A1(n816), .A2(n670), .A3(n845), .ZN(n758) );
  ND2D0 U416 ( .A1(n670), .A2(n848), .ZN(n588) );
  CKND2D1 U417 ( .A1(n842), .A2(n670), .ZN(n730) );
  OAI32D0 U418 ( .A1(n557), .A2(n756), .A3(n434), .B1(n516), .B2(n515), .ZN(
        n517) );
  OAI221D0 U419 ( .A1(n737), .A2(n683), .B1(n745), .B2(n702), .C(n682), .ZN(
        n690) );
  OAI222D0 U420 ( .A1(n745), .A2(n555), .B1(n641), .B2(n717), .C1(n746), .C2(
        n684), .ZN(n459) );
  OAI22D0 U421 ( .A1(n742), .A2(n754), .B1(n601), .B2(n429), .ZN(n608) );
  NR2D1 U422 ( .A1(n793), .A2(n758), .ZN(n740) );
  OA21D0 U423 ( .A1(n683), .A2(n793), .B(n613), .Z(n617) );
  OAI22D0 U424 ( .A1(n443), .A2(n610), .B1(n793), .B2(n609), .ZN(n611) );
  OAI22D0 U425 ( .A1(n641), .A2(n742), .B1(n429), .B2(n771), .ZN(n499) );
  OA222D0 U426 ( .A1(n746), .A2(n434), .B1(n744), .B2(n429), .C1(n748), .C2(
        n742), .Z(n757) );
  AOI32D0 U427 ( .A1(n445), .A2(n793), .A3(n817), .B1(n828), .B2(n632), .ZN(
        n633) );
  AOI22D0 U428 ( .A1(n793), .A2(n817), .B1(n813), .B2(n804), .ZN(n589) );
  OAI22D0 U429 ( .A1(n793), .A2(n719), .B1(n451), .B2(n730), .ZN(n527) );
  NR3D0 U430 ( .A1(n793), .A2(n444), .A3(n684), .ZN(n593) );
  OAI222D0 U431 ( .A1(n437), .A2(n650), .B1(n649), .B2(n783), .C1(n648), .C2(
        n782), .ZN(n651) );
  AOI22D0 U432 ( .A1(n825), .A2(n795), .B1(n823), .B2(n437), .ZN(n572) );
  CKND2D0 U433 ( .A1(n437), .A2(n737), .ZN(n735) );
  AOI31D0 U434 ( .A1(n437), .A2(n827), .A3(n796), .B(n826), .ZN(n495) );
  CKND2D0 U435 ( .A1(n444), .A2(n437), .ZN(n702) );
  CKND2D0 U436 ( .A1(n437), .A2(n445), .ZN(n744) );
  NR3D0 U437 ( .A1(n815), .A2(n800), .A3(n671), .ZN(n648) );
  AO221D0 U438 ( .A1(n800), .A2(n833), .B1(n797), .B2(n815), .C(n699), .Z(n652) );
  OAI222D0 U439 ( .A1(n641), .A2(n721), .B1(n589), .B2(n730), .C1(n635), .C2(
        n664), .ZN(n482) );
  INR2D1 U440 ( .A1(n522), .B1(n664), .ZN(n709) );
  NR4D0 U441 ( .A1(n768), .A2(n756), .A3(n664), .A4(n443), .ZN(n738) );
  OAI222D0 U442 ( .A1(n723), .A2(n596), .B1(n730), .B2(n435), .C1(n635), .C2(
        n759), .ZN(n547) );
  NR3D0 U443 ( .A1(n827), .A2(n450), .A3(n723), .ZN(n531) );
  NR2D1 U444 ( .A1(n832), .A2(n811), .ZN(n516) );
  NR2D1 U445 ( .A1(n635), .A2(n720), .ZN(n739) );
  OAI22D0 U446 ( .A1(n451), .A2(n719), .B1(n449), .B2(n635), .ZN(n637) );
  OAI21D0 U447 ( .A1(n641), .A2(n729), .B(n783), .ZN(n472) );
  AOI31D0 U448 ( .A1(n730), .A2(n729), .A3(n728), .B(n727), .ZN(n731) );
  AOI22D0 U449 ( .A1(n852), .A2(n525), .B1(n691), .B2(n524), .ZN(n526) );
  AOI21D0 U450 ( .A1(n729), .A2(n669), .B(n437), .ZN(n627) );
  OAI22D0 U451 ( .A1(a[6]), .A2(n444), .B1(n445), .B2(n756), .ZN(n548) );
  OAI211D0 U452 ( .A1(n445), .A2(n781), .B(n625), .C(n748), .ZN(n537) );
  INVD1 U453 ( .I(n737), .ZN(n797) );
  INVD1 U454 ( .I(n754), .ZN(n821) );
  NR2D0 U455 ( .A1(n833), .A2(n829), .ZN(n673) );
  AOI221D1 U456 ( .A1(n842), .A2(n653), .B1(n845), .B2(n652), .C(n651), .ZN(
        n660) );
  OAI22D0 U457 ( .A1(n460), .A2(n779), .B1(n746), .B2(n634), .ZN(n461) );
  NR4D0 U458 ( .A1(n684), .A2(n751), .A3(n779), .A4(n819), .ZN(n656) );
  AOI21D0 U459 ( .A1(n774), .A2(n744), .B(n779), .ZN(n626) );
endmodule


module aes_sbox_10 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n65, n70, n71, n142, n148, n175, n176, n192, n342, n405, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865;

  AN2XD1 U28 ( .A1(n723), .A2(n425), .Z(n727) );
  OA21D1 U35 ( .A1(n708), .A2(n707), .B(n706), .Z(n713) );
  OR3D1 U88 ( .A1(n678), .A2(n813), .A3(n452), .Z(n639) );
  OR4D1 U199 ( .A1(n663), .A2(n581), .A3(n526), .A4(n525), .Z(n528) );
  AN2XD1 U215 ( .A1(n527), .A2(n811), .Z(n526) );
  AN2XD1 U271 ( .A1(n539), .A2(n734), .Z(n473) );
  AO21D1 U297 ( .A1(n799), .A2(n837), .B(n737), .Z(n466) );
  OAI222D1 U1 ( .A1(n786), .A2(n588), .B1(n778), .B2(n643), .C1(n501), .C2(
        n766), .ZN(n502) );
  INVD2 U2 ( .I(n709), .ZN(n850) );
  NR2XD1 U3 ( .A1(n839), .A2(n850), .ZN(n645) );
  CKND2D1 U4 ( .A1(n831), .A2(n850), .ZN(n603) );
  CKND2D0 U5 ( .A1(n830), .A2(n850), .ZN(n641) );
  CKND2D0 U6 ( .A1(n677), .A2(n850), .ZN(n595) );
  CKND2D2 U7 ( .A1(n854), .A2(n448), .ZN(n643) );
  ND2D1 U8 ( .A1(n442), .A2(n807), .ZN(n731) );
  AOI221D1 U9 ( .A1(n862), .A2(n448), .B1(n854), .B2(n809), .C(n638), .ZN(n669) );
  IND4D2 U10 ( .A1(n796), .B1(n795), .B2(n794), .B3(n793), .ZN(d[0]) );
  BUFFD6 U11 ( .I(a[3]), .Z(n444) );
  CKND2D1 U12 ( .A1(n829), .A2(n836), .ZN(n662) );
  INVD1 U13 ( .I(n750), .ZN(n809) );
  AOI221D1 U14 ( .A1(n861), .A2(n651), .B1(n858), .B2(n804), .C(n650), .ZN(
        n668) );
  AOI221D1 U15 ( .A1(n803), .A2(n852), .B1(n71), .B2(n865), .C(n597), .ZN(n630) );
  INVD1 U16 ( .I(n772), .ZN(n830) );
  INVD1 U17 ( .I(n671), .ZN(n807) );
  ND4D2 U18 ( .A1(n630), .A2(n629), .A3(n628), .A4(n627), .ZN(d[3]) );
  AOI221D1 U19 ( .A1(n817), .A2(n607), .B1(n844), .B2(n606), .C(n605), .ZN(
        n629) );
  ND2D1 U20 ( .A1(n802), .A2(n442), .ZN(n562) );
  ND2D1 U21 ( .A1(n801), .A2(n815), .ZN(n691) );
  ND2D1 U22 ( .A1(n815), .A2(n821), .ZN(n758) );
  INVD1 U23 ( .I(n788), .ZN(n804) );
  INVD3 U24 ( .I(n444), .ZN(n815) );
  INVD1 U25 ( .I(n691), .ZN(n816) );
  NR3D0 U26 ( .A1(n148), .A2(n175), .A3(n693), .ZN(n695) );
  OAI222D0 U27 ( .A1(n710), .A2(n734), .B1(n442), .B2(n543), .C1(n788), .C2(
        n777), .ZN(n544) );
  OAI221D0 U29 ( .A1(n741), .A2(n734), .B1(n709), .B2(n747), .C(n599), .ZN(
        n607) );
  INVD1 U30 ( .I(n778), .ZN(n817) );
  INVD2 U31 ( .I(n783), .ZN(n844) );
  ND2D1 U32 ( .A1(n688), .A2(n847), .ZN(n732) );
  INVD2 U33 ( .I(n754), .ZN(n847) );
  NR2D0 U34 ( .A1(n692), .A2(n520), .ZN(n440) );
  OAI222D0 U36 ( .A1(n433), .A2(n752), .B1(n696), .B2(n692), .C1(n758), .C2(
        n559), .ZN(n537) );
  AN4D1 U37 ( .A1(n677), .A2(n819), .A3(n442), .A4(n847), .Z(n525) );
  ND3D0 U38 ( .A1(n818), .A2(n677), .A3(n847), .ZN(n762) );
  INVD2 U39 ( .I(n71), .ZN(n425) );
  AN2XD1 U40 ( .A1(n442), .A2(n801), .Z(n65) );
  OA221D0 U41 ( .A1(n691), .A2(n681), .B1(n680), .B2(n788), .C(n679), .Z(n70)
         );
  AN2D1 U42 ( .A1(n450), .A2(n442), .Z(n71) );
  ND2D1 U43 ( .A1(n832), .A2(n844), .ZN(n726) );
  NR2D1 U44 ( .A1(n806), .A2(n802), .ZN(n479) );
  CKND2D2 U45 ( .A1(n804), .A2(n448), .ZN(n559) );
  NR2XD0 U46 ( .A1(n781), .A2(n780), .ZN(n782) );
  OAI22D1 U47 ( .A1(n474), .A2(n714), .B1(n473), .B2(n763), .ZN(n475) );
  AOI221D2 U48 ( .A1(n697), .A2(n747), .B1(n449), .B2(n856), .C(n561), .ZN(
        n566) );
  AOI211XD1 U49 ( .A1(n805), .A2(n825), .B(n828), .C(n700), .ZN(n701) );
  AOI211XD1 U50 ( .A1(n861), .A2(n499), .B(n498), .C(n497), .ZN(n513) );
  CKND2D1 U51 ( .A1(n447), .A2(n829), .ZN(n730) );
  OA221D0 U52 ( .A1(n741), .A2(n691), .B1(n749), .B2(n708), .C(n690), .Z(n437)
         );
  AOI221D1 U53 ( .A1(n799), .A2(n689), .B1(n688), .B2(n807), .C(n687), .ZN(
        n690) );
  INVD1 U54 ( .I(n760), .ZN(n861) );
  OA221D1 U55 ( .A1(n752), .A2(n760), .B1(n775), .B2(n768), .C(n142), .Z(n533)
         );
  ND2D2 U56 ( .A1(n447), .A2(n836), .ZN(n760) );
  OAI22D1 U57 ( .A1(n726), .A2(n755), .B1(n801), .B2(n732), .ZN(n670) );
  OAI222D1 U58 ( .A1(n671), .A2(n771), .B1(n442), .B2(n563), .C1(n753), .C2(
        n562), .ZN(n564) );
  AOI221D1 U59 ( .A1(n847), .A2(n615), .B1(n614), .B2(n448), .C(n613), .ZN(
        n628) );
  INVD1 U60 ( .I(n746), .ZN(n799) );
  CKND2D1 U61 ( .A1(n442), .A2(n451), .ZN(n746) );
  ND2D3 U62 ( .A1(n836), .A2(n841), .ZN(n754) );
  INVD2 U63 ( .I(n447), .ZN(n841) );
  ND2D0 U64 ( .A1(n446), .A2(n841), .ZN(n711) );
  ND2D2 U65 ( .A1(a[6]), .A2(n841), .ZN(n783) );
  CKND2D1 U66 ( .A1(n834), .A2(n841), .ZN(n631) );
  CKND2D0 U67 ( .A1(n829), .A2(n841), .ZN(n616) );
  AOI21D1 U68 ( .A1(n444), .A2(n861), .B(n820), .ZN(n773) );
  ND2D2 U69 ( .A1(n448), .A2(n451), .ZN(n747) );
  OAI22D0 U70 ( .A1(n747), .A2(n711), .B1(n645), .B2(n741), .ZN(n646) );
  CKND0 U71 ( .I(n747), .ZN(n798) );
  OA221D0 U72 ( .A1(n616), .A2(n590), .B1(n444), .B2(n777), .C(n706), .Z(n142)
         );
  INVD2 U73 ( .I(n775), .ZN(n813) );
  INVD2 U74 ( .I(n768), .ZN(n834) );
  INVD2 U75 ( .I(n451), .ZN(n450) );
  ND2D1 U76 ( .A1(n450), .A2(n443), .ZN(n750) );
  INVD2 U77 ( .I(n559), .ZN(n805) );
  AOI221D1 U78 ( .A1(n844), .A2(n660), .B1(n847), .B2(n659), .C(n658), .ZN(
        n667) );
  CKND2D1 U79 ( .A1(n449), .A2(n444), .ZN(n785) );
  OAI222D0 U80 ( .A1(n574), .A2(n714), .B1(n573), .B2(n746), .C1(n449), .C2(
        n572), .ZN(n575) );
  NR4D1 U81 ( .A1(n537), .A2(n536), .A3(n535), .A4(n600), .ZN(n538) );
  AOI21D0 U82 ( .A1(n778), .A2(n748), .B(n783), .ZN(n633) );
  CKND1 U83 ( .I(n785), .ZN(n819) );
  OAI222D0 U84 ( .A1(n749), .A2(n559), .B1(n648), .B2(n425), .C1(n750), .C2(
        n692), .ZN(n460) );
  ND2D1 U85 ( .A1(n444), .A2(n829), .ZN(n749) );
  AOI221D1 U86 ( .A1(n468), .A2(n809), .B1(n854), .B2(n819), .C(n467), .ZN(
        n469) );
  CKND0 U87 ( .I(n730), .ZN(n860) );
  OAI222D1 U89 ( .A1(n649), .A2(n648), .B1(n763), .B2(n765), .C1(n647), .C2(
        n775), .ZN(n650) );
  OAI222D1 U90 ( .A1(n534), .A2(n778), .B1(n433), .B2(n631), .C1(n533), .C2(
        n425), .ZN(n546) );
  AOI221D1 U91 ( .A1(n477), .A2(n451), .B1(n823), .B2(n476), .C(n475), .ZN(
        n484) );
  AOI221D1 U92 ( .A1(n705), .A2(n860), .B1(n818), .B2(n704), .C(n703), .ZN(
        n719) );
  ND2D2 U93 ( .A1(n450), .A2(n801), .ZN(n788) );
  INR4D0 U94 ( .A1(n676), .B1(n675), .B2(n674), .B3(n857), .ZN(n685) );
  AOI221D1 U95 ( .A1(n802), .A2(n860), .B1(n811), .B2(n839), .C(n466), .ZN(
        n470) );
  AOI21D2 U96 ( .A1(n816), .A2(n449), .B(n805), .ZN(n589) );
  CKND2D2 U97 ( .A1(n444), .A2(n821), .ZN(n752) );
  OAI211D0 U98 ( .A1(n446), .A2(n785), .B(n632), .C(n752), .ZN(n541) );
  OAI21D0 U99 ( .A1(n662), .A2(n752), .B(n732), .ZN(n542) );
  AOI221D2 U100 ( .A1(n442), .A2(n570), .B1(n844), .B2(n569), .C(n568), .ZN(
        n586) );
  AOI211XD1 U101 ( .A1(n831), .A2(n593), .B(n591), .C(n592), .ZN(n594) );
  AOI222D1 U102 ( .A1(n809), .A2(n832), .B1(n807), .B2(n489), .C1(n803), .C2(
        n835), .ZN(n494) );
  OAI222D1 U103 ( .A1(n433), .A2(n539), .B1(n494), .B2(n754), .C1(n493), .C2(
        n758), .ZN(n498) );
  AOI221D1 U104 ( .A1(n838), .A2(n826), .B1(n824), .B2(n577), .C(n853), .ZN(
        n501) );
  INVD6 U105 ( .I(n445), .ZN(n821) );
  AOI211XD0 U106 ( .A1(n865), .A2(n810), .B(n487), .C(n670), .ZN(n514) );
  OAI221D1 U107 ( .A1(n673), .A2(n683), .B1(n672), .B2(n671), .C(n848), .ZN(
        n675) );
  ND2D2 U108 ( .A1(n821), .A2(n829), .ZN(n772) );
  OAI22D0 U109 ( .A1(n461), .A2(n783), .B1(n750), .B2(n641), .ZN(n462) );
  ND4D2 U110 ( .A1(n514), .A2(n513), .A3(n512), .A4(n511), .ZN(d[6]) );
  INVD6 U111 ( .I(n446), .ZN(n829) );
  OAI32D1 U112 ( .A1(n590), .A2(n747), .A3(n692), .B1(n589), .B2(n768), .ZN(
        n591) );
  ND2D2 U113 ( .A1(n832), .A2(n850), .ZN(n733) );
  INVD2 U114 ( .I(n617), .ZN(n832) );
  ND2D2 U115 ( .A1(n447), .A2(a[6]), .ZN(n709) );
  BUFFD4 U116 ( .I(a[7]), .Z(n447) );
  OAI222D1 U117 ( .A1(n567), .A2(n760), .B1(n691), .B2(n566), .C1(n565), .C2(
        n754), .ZN(n568) );
  ND2D2 U118 ( .A1(n444), .A2(n801), .ZN(n775) );
  NR3D1 U119 ( .A1(n429), .A2(n430), .A3(n686), .ZN(n721) );
  ND2D2 U120 ( .A1(n446), .A2(n821), .ZN(n768) );
  INVD2 U121 ( .I(a[6]), .ZN(n836) );
  AOI221D1 U122 ( .A1(n863), .A2(n451), .B1(n845), .B2(n425), .C(n532), .ZN(
        n534) );
  NR2XD1 U123 ( .A1(n65), .A2(n799), .ZN(n696) );
  ND4D2 U124 ( .A1(n486), .A2(n485), .A3(n484), .A4(n483), .ZN(d[7]) );
  AOI21D1 U125 ( .A1(n863), .A2(n818), .B(n857), .ZN(n572) );
  ND2D3 U126 ( .A1(n449), .A2(n448), .ZN(n741) );
  CKND2 U127 ( .I(n451), .ZN(n449) );
  AOI221D1 U128 ( .A1(n849), .A2(n448), .B1(n859), .B2(n449), .C(n646), .ZN(
        n647) );
  CKND1 U129 ( .I(n786), .ZN(n849) );
  CKND3 U130 ( .I(a[1]), .ZN(n451) );
  NR4D1 U131 ( .A1(n790), .A2(n791), .A3(n792), .A4(n789), .ZN(n793) );
  OAI222D1 U132 ( .A1(n784), .A2(n783), .B1(n444), .B2(n842), .C1(n782), .C2(
        n448), .ZN(n790) );
  OA222D0 U133 ( .A1(n750), .A2(n749), .B1(n748), .B2(n747), .C1(n752), .C2(
        n746), .Z(n761) );
  ND2D1 U134 ( .A1(n445), .A2(n815), .ZN(n714) );
  ND4D2 U135 ( .A1(n721), .A2(n720), .A3(n719), .A4(n718), .ZN(d[1]) );
  AN2XD1 U136 ( .A1(n800), .A2(n694), .Z(n148) );
  CKAN2D1 U137 ( .A1(n835), .A2(n65), .Z(n175) );
  INVD1 U138 ( .I(n741), .ZN(n800) );
  CKAN2D1 U139 ( .A1(n824), .A2(n798), .Z(n176) );
  CKAN2D1 U140 ( .A1(n833), .A2(n809), .Z(n192) );
  NR3D0 U141 ( .A1(n176), .A2(n192), .A3(n564), .ZN(n565) );
  NR2D1 U142 ( .A1(n812), .A2(n637), .ZN(n342) );
  NR2D0 U143 ( .A1(n559), .A2(n539), .ZN(n405) );
  NR2D0 U144 ( .A1(n538), .A2(n783), .ZN(n424) );
  OR3D1 U145 ( .A1(n342), .A2(n405), .A3(n424), .Z(n545) );
  ND2D1 U146 ( .A1(n837), .A2(n826), .ZN(n539) );
  NR4D1 U147 ( .A1(n547), .A2(n546), .A3(n545), .A4(n544), .ZN(n548) );
  CKBD4 U148 ( .I(n797), .Z(n448) );
  CKND0 U149 ( .I(n442), .ZN(n797) );
  AOI221D1 U150 ( .A1(n844), .A2(n503), .B1(n803), .B2(n516), .C(n502), .ZN(
        n512) );
  AOI221D1 U151 ( .A1(n802), .A2(n826), .B1(n810), .B2(n833), .C(n769), .ZN(
        n784) );
  ND4D2 U152 ( .A1(n586), .A2(n587), .A3(n585), .A4(n584), .ZN(d[4]) );
  AOI221D1 U153 ( .A1(n814), .A2(n577), .B1(n576), .B2(n824), .C(n575), .ZN(
        n585) );
  OAI222D1 U154 ( .A1(n648), .A2(n641), .B1(n596), .B2(n595), .C1(n594), .C2(
        n760), .ZN(n597) );
  ND4D2 U155 ( .A1(n669), .A2(n668), .A3(n667), .A4(n666), .ZN(d[2]) );
  NR2D1 U156 ( .A1(n707), .A2(n747), .ZN(n737) );
  NR2D0 U157 ( .A1(n845), .A2(n856), .ZN(n673) );
  ND2D0 U158 ( .A1(n832), .A2(n861), .ZN(n682) );
  ND2D0 U159 ( .A1(n444), .A2(n452), .ZN(n683) );
  NR2D0 U160 ( .A1(n442), .A2(n685), .ZN(n426) );
  NR2D0 U161 ( .A1(n684), .A2(n754), .ZN(n427) );
  NR2D0 U162 ( .A1(n683), .A2(n682), .ZN(n428) );
  OR3D1 U163 ( .A1(n426), .A2(n427), .A3(n428), .Z(n686) );
  CKAN2D1 U164 ( .A1(n852), .A2(n811), .Z(n429) );
  CKAN2D1 U165 ( .A1(n697), .A2(n804), .Z(n430) );
  CKND2D0 U166 ( .A1(n831), .A2(n800), .ZN(n431) );
  CKND2D0 U167 ( .A1(n823), .A2(n807), .ZN(n432) );
  AN3XD1 U168 ( .A1(n431), .A2(n432), .A3(n70), .Z(n684) );
  INVD1 U169 ( .I(n763), .ZN(n811) );
  CKND2D0 U170 ( .A1(n442), .A2(n801), .ZN(n433) );
  INVD4 U171 ( .I(n443), .ZN(n801) );
  INR2D1 U172 ( .A1(n764), .B1(n505), .ZN(n506) );
  BUFFD6 U173 ( .I(a[0]), .Z(n442) );
  ND2D0 U174 ( .A1(n813), .A2(n856), .ZN(n571) );
  NR2D0 U175 ( .A1(n809), .A2(n71), .ZN(n620) );
  CKND0 U176 ( .I(n724), .ZN(n846) );
  OAI31D1 U177 ( .A1(n678), .A2(n65), .A3(n820), .B(n677), .ZN(n679) );
  NR2XD0 U178 ( .A1(n835), .A2(n831), .ZN(n680) );
  NR2D0 U179 ( .A1(n631), .A2(n746), .ZN(n770) );
  AOI21D1 U180 ( .A1(n822), .A2(n864), .B(n851), .ZN(n573) );
  CKND2D0 U181 ( .A1(n688), .A2(n850), .ZN(n637) );
  CKND2D0 U182 ( .A1(n833), .A2(n850), .ZN(n765) );
  CKND2D0 U183 ( .A1(n824), .A2(n850), .ZN(n612) );
  CKND2D0 U184 ( .A1(n785), .A2(n691), .ZN(n529) );
  ND2D0 U185 ( .A1(n443), .A2(n815), .ZN(n778) );
  NR2D0 U186 ( .A1(n445), .A2(n836), .ZN(n468) );
  AOI22D1 U187 ( .A1(n832), .A2(n818), .B1(n807), .B2(n829), .ZN(n563) );
  ND2D0 U188 ( .A1(n443), .A2(n821), .ZN(n632) );
  CKND2D1 U189 ( .A1(n776), .A2(n730), .ZN(n577) );
  BUFFD4 U190 ( .I(a[5]), .Z(n446) );
  CKND0 U191 ( .I(n777), .ZN(n862) );
  CKND0 U192 ( .I(n588), .ZN(n814) );
  OAI22D0 U193 ( .A1(n758), .A2(n755), .B1(n661), .B2(n741), .ZN(n524) );
  OAI31D0 U194 ( .A1(n802), .A2(n799), .A3(n813), .B(n862), .ZN(n495) );
  ND2D0 U195 ( .A1(n847), .A2(n834), .ZN(n786) );
  AOI22D0 U196 ( .A1(n863), .A2(n804), .B1(n819), .B2(n849), .ZN(n553) );
  ND2D0 U197 ( .A1(n817), .A2(n449), .ZN(n723) );
  NR2D0 U198 ( .A1(n642), .A2(n725), .ZN(n743) );
  CKND2D0 U200 ( .A1(n864), .A2(n826), .ZN(n787) );
  NR2D0 U201 ( .A1(n65), .A2(n798), .ZN(n621) );
  ND2D0 U202 ( .A1(n824), .A2(n864), .ZN(n764) );
  CKND2D0 U203 ( .A1(n823), .A2(n847), .ZN(n676) );
  NR2D0 U204 ( .A1(n722), .A2(n859), .ZN(n728) );
  CKND0 U205 ( .I(n643), .ZN(n855) );
  CKND2D0 U206 ( .A1(n731), .A2(n741), .ZN(n593) );
  CKND2D0 U207 ( .A1(n65), .A2(n834), .ZN(n652) );
  OAI22D0 U208 ( .A1(n448), .A2(n724), .B1(n452), .B2(n734), .ZN(n532) );
  CKND2D0 U209 ( .A1(n785), .A2(n559), .ZN(n560) );
  NR2D0 U210 ( .A1(n754), .A2(n772), .ZN(n697) );
  AOI22D0 U211 ( .A1(n831), .A2(n807), .B1(n804), .B2(n833), .ZN(n453) );
  NR2D0 U212 ( .A1(n813), .A2(n806), .ZN(n454) );
  NR2D0 U213 ( .A1(n863), .A2(n849), .ZN(n465) );
  CKND2D0 U214 ( .A1(n832), .A2(n451), .ZN(n681) );
  AOI22D0 U216 ( .A1(n854), .A2(n530), .B1(n697), .B2(n529), .ZN(n531) );
  OAI32D0 U217 ( .A1(n562), .A2(n760), .A3(n749), .B1(n521), .B2(n520), .ZN(
        n522) );
  NR2D0 U218 ( .A1(n834), .A2(n813), .ZN(n521) );
  CKND2D1 U219 ( .A1(n496), .A2(n495), .ZN(n497) );
  OAI22D0 U220 ( .A1(n648), .A2(n746), .B1(n747), .B2(n775), .ZN(n504) );
  OAI31D0 U221 ( .A1(n741), .A2(n825), .A3(n754), .B(n740), .ZN(n745) );
  AOI22D0 U222 ( .A1(n448), .A2(n819), .B1(n815), .B2(n806), .ZN(n596) );
  AOI32D0 U223 ( .A1(n802), .A2(n448), .A3(n835), .B1(n800), .B2(n555), .ZN(
        n557) );
  CKND2D0 U224 ( .A1(n753), .A2(n748), .ZN(n555) );
  OAI21D0 U225 ( .A1(n753), .A2(n616), .B(n641), .ZN(n516) );
  OAI22D0 U226 ( .A1(n746), .A2(n758), .B1(n608), .B2(n747), .ZN(n615) );
  NR2D0 U227 ( .A1(n827), .A2(n832), .ZN(n608) );
  CKND0 U228 ( .I(n753), .ZN(n825) );
  OAI22D0 U229 ( .A1(n768), .A2(n778), .B1(n449), .B2(n767), .ZN(n769) );
  AOI22D0 U230 ( .A1(n813), .A2(n834), .B1(n816), .B2(n829), .ZN(n767) );
  NR2D0 U231 ( .A1(n448), .A2(n762), .ZN(n744) );
  CKND2D0 U232 ( .A1(n809), .A2(n448), .ZN(n710) );
  AOI31D0 U233 ( .A1(n734), .A2(n733), .A3(n732), .B(n731), .ZN(n735) );
  NR2D0 U234 ( .A1(n515), .A2(n671), .ZN(n576) );
  INR2D0 U235 ( .A1(n527), .B1(n671), .ZN(n715) );
  AOI22D0 U236 ( .A1(n838), .A2(n751), .B1(n840), .B2(n807), .ZN(n759) );
  CKND2D0 U237 ( .A1(n798), .A2(n815), .ZN(n725) );
  OAI21D0 U238 ( .A1(n648), .A2(n733), .B(n787), .ZN(n477) );
  CKND0 U239 ( .I(n707), .ZN(n864) );
  OAI211D0 U240 ( .A1(n829), .A2(n758), .B(n775), .C(n753), .ZN(n689) );
  CKND0 U241 ( .I(n562), .ZN(n803) );
  ND2D0 U242 ( .A1(n449), .A2(n471), .ZN(n434) );
  CKND2D0 U243 ( .A1(n828), .A2(n838), .ZN(n435) );
  AOI21D0 U244 ( .A1(n849), .A2(n818), .B(n756), .ZN(n757) );
  OAI21D0 U245 ( .A1(n442), .A2(n692), .B(n752), .ZN(n489) );
  OAI22D0 U246 ( .A1(n452), .A2(n637), .B1(n636), .B2(n746), .ZN(n638) );
  AOI211XD0 U247 ( .A1(n843), .A2(n810), .B(n492), .C(n491), .ZN(n493) );
  CKND0 U248 ( .I(n616), .ZN(n843) );
  AOI22D0 U249 ( .A1(n804), .A2(n838), .B1(n813), .B2(n821), .ZN(n774) );
  AOI21D0 U250 ( .A1(n808), .A2(n847), .B(n576), .ZN(n518) );
  MAOI22D0 U251 ( .A1(n859), .A2(n815), .B1(n632), .B2(n776), .ZN(n519) );
  NR2D0 U252 ( .A1(n811), .A2(n809), .ZN(n472) );
  CKND2D0 U253 ( .A1(n818), .A2(n821), .ZN(n609) );
  NR2XD0 U254 ( .A1(n653), .A2(n770), .ZN(n611) );
  AOI211D0 U255 ( .A1(n820), .A2(n442), .B(n818), .C(n811), .ZN(n610) );
  NR2D0 U256 ( .A1(n798), .A2(n807), .ZN(n656) );
  AOI211XD0 U257 ( .A1(n845), .A2(n442), .B(n644), .C(n855), .ZN(n649) );
  OAI22D0 U258 ( .A1(n452), .A2(n724), .B1(n449), .B2(n642), .ZN(n644) );
  AOI32D0 U259 ( .A1(n447), .A2(n821), .A3(n802), .B1(n807), .B2(n455), .ZN(
        n456) );
  NR2D0 U260 ( .A1(n859), .A2(n697), .ZN(n457) );
  OAI22D0 U261 ( .A1(n447), .A2(n662), .B1(n753), .B2(n730), .ZN(n455) );
  AOI21D0 U262 ( .A1(n858), .A2(n449), .B(n697), .ZN(n698) );
  ND4D0 U263 ( .A1(n799), .A2(n838), .A3(n445), .A4(n447), .ZN(n729) );
  OAI21D0 U264 ( .A1(n754), .A2(n617), .B(n724), .ZN(n598) );
  AOI31D0 U265 ( .A1(n445), .A2(n836), .A3(n813), .B(n699), .ZN(n478) );
  AOI211D0 U266 ( .A1(n779), .A2(n662), .B(n590), .C(n746), .ZN(n480) );
  OAI31D0 U267 ( .A1(n750), .A2(n779), .A3(n752), .B(n619), .ZN(n626) );
  AOI33D0 U268 ( .A1(n618), .A2(n836), .A3(n804), .B1(n856), .B2(n815), .B3(
        n800), .ZN(n619) );
  OAI22D0 U269 ( .A1(n444), .A2(n617), .B1(n448), .B2(n616), .ZN(n618) );
  CKND0 U270 ( .I(n739), .ZN(n812) );
  AOI21D0 U272 ( .A1(n859), .A2(n819), .B(n699), .ZN(n702) );
  CKND2D0 U273 ( .A1(n425), .A2(n815), .ZN(n579) );
  NR2D0 U274 ( .A1(n733), .A2(n444), .ZN(n699) );
  OAI22D0 U275 ( .A1(n836), .A2(n714), .B1(n821), .B2(n662), .ZN(n654) );
  AOI21D0 U276 ( .A1(n691), .A2(n590), .B(n746), .ZN(n458) );
  AO31D0 U277 ( .A1(n804), .A2(n861), .A3(n688), .B(n722), .Z(n467) );
  AOI22D0 U278 ( .A1(n809), .A2(n442), .B1(n449), .B2(n818), .ZN(n488) );
  OAI21D0 U279 ( .A1(n713), .A2(n741), .B(n712), .ZN(n717) );
  CKND2D0 U280 ( .A1(n443), .A2(n741), .ZN(n739) );
  CKND2D1 U281 ( .A1(n601), .A2(n602), .ZN(n606) );
  CKND0 U282 ( .I(n779), .ZN(n840) );
  CKND2D0 U283 ( .A1(n692), .A2(n752), .ZN(n694) );
  AOI32D0 U284 ( .A1(n446), .A2(n448), .A3(n819), .B1(n830), .B2(n639), .ZN(
        n640) );
  AOI21D0 U285 ( .A1(n824), .A2(n860), .B(n699), .ZN(n508) );
  AOI32D0 U286 ( .A1(n445), .A2(n841), .A3(n817), .B1(n818), .B2(n552), .ZN(
        n554) );
  BUFFD4 U287 ( .I(a[4]), .Z(n445) );
  BUFFD4 U288 ( .I(a[2]), .Z(n443) );
  INVD1 U289 ( .I(n682), .ZN(n863) );
  INVD1 U290 ( .I(n787), .ZN(n865) );
  INVD1 U291 ( .I(n571), .ZN(n857) );
  AOI222D0 U292 ( .A1(n809), .A2(n826), .B1(n824), .B2(n65), .C1(n833), .C2(
        n807), .ZN(n556) );
  INVD1 U293 ( .I(n758), .ZN(n823) );
  INVD1 U294 ( .I(n595), .ZN(n859) );
  AO221D0 U295 ( .A1(n802), .A2(n835), .B1(n800), .B2(n817), .C(n705), .Z(n659) );
  ND2D1 U296 ( .A1(n813), .A2(n449), .ZN(n588) );
  INVD1 U298 ( .I(n642), .ZN(n856) );
  INVD1 U299 ( .I(n710), .ZN(n810) );
  INVD1 U300 ( .I(n558), .ZN(n822) );
  INVD1 U301 ( .I(n637), .ZN(n852) );
  ND2D1 U302 ( .A1(n822), .A2(n838), .ZN(n706) );
  NR2D1 U303 ( .A1(n818), .A2(n825), .ZN(n661) );
  INVD1 U304 ( .I(n726), .ZN(n845) );
  INVD1 U305 ( .I(n755), .ZN(n802) );
  ND2D1 U306 ( .A1(n71), .A2(n827), .ZN(n604) );
  INVD1 U307 ( .I(n733), .ZN(n854) );
  INVD1 U308 ( .I(n603), .ZN(n853) );
  INVD1 U309 ( .I(n612), .ZN(n851) );
  OAI222D0 U310 ( .A1(n755), .A2(n692), .B1(n488), .B2(n768), .C1(n449), .C2(
        n753), .ZN(n499) );
  OAI222D0 U311 ( .A1(n763), .A2(n771), .B1(n785), .B2(n652), .C1(n752), .C2(
        n710), .ZN(n660) );
  OAI222D0 U312 ( .A1(n748), .A2(n425), .B1(n772), .B2(n588), .C1(n753), .C2(
        n763), .ZN(n592) );
  AOI221D0 U313 ( .A1(n805), .A2(n835), .B1(n830), .B2(n560), .C(n705), .ZN(
        n567) );
  OAI222D0 U314 ( .A1(n648), .A2(n726), .B1(n596), .B2(n734), .C1(n642), .C2(
        n671), .ZN(n487) );
  NR4D0 U315 ( .A1(n665), .A2(n664), .A3(n663), .A4(n744), .ZN(n666) );
  AOI221D0 U316 ( .A1(n737), .A2(n817), .B1(n816), .B2(n736), .C(n735), .ZN(
        n795) );
  NR4D0 U317 ( .A1(n745), .A2(n744), .A3(n743), .A4(n742), .ZN(n794) );
  INVD1 U318 ( .I(n752), .ZN(n824) );
  NR4D0 U319 ( .A1(n482), .A2(n481), .A3(n716), .A4(n480), .ZN(n483) );
  NR4D0 U320 ( .A1(n583), .A2(n582), .A3(n581), .A4(n742), .ZN(n584) );
  AOI221D0 U321 ( .A1(n813), .A2(n846), .B1(n854), .B2(n819), .C(n551), .ZN(
        n587) );
  NR2D1 U322 ( .A1(n626), .A2(n625), .ZN(n627) );
  OAI221D0 U323 ( .A1(n449), .A2(n676), .B1(n725), .B2(n682), .C(n531), .ZN(
        n547) );
  ND3D1 U324 ( .A1(n550), .A2(n549), .A3(n548), .ZN(d[5]) );
  AOI211D1 U325 ( .A1(n864), .A2(n524), .B(n523), .C(n522), .ZN(n550) );
  INR4D0 U326 ( .A1(n762), .B1(n528), .B2(n743), .B3(n715), .ZN(n549) );
  AN3XD1 U327 ( .A1(n434), .A2(n435), .A3(n436), .Z(n485) );
  NR3D0 U328 ( .A1(n439), .A2(n440), .A3(n441), .ZN(n436) );
  OAI221D0 U329 ( .A1(n454), .A2(n617), .B1(n778), .B2(n425), .C(n453), .ZN(
        n464) );
  ND2D1 U330 ( .A1(n452), .A2(n801), .ZN(n755) );
  AOI31D1 U331 ( .A1(n850), .A2(n739), .A3(n825), .B(n738), .ZN(n740) );
  ND2D1 U332 ( .A1(n844), .A2(n830), .ZN(n724) );
  NR2D1 U333 ( .A1(n632), .A2(n425), .ZN(n705) );
  NR4D0 U334 ( .A1(n717), .A2(n738), .A3(n716), .A4(n715), .ZN(n718) );
  OA221D0 U335 ( .A1(n641), .A2(n425), .B1(n760), .B2(n437), .C(n438), .Z(n720) );
  INVD1 U336 ( .I(n714), .ZN(n826) );
  NR3D0 U337 ( .A1(n425), .A2(n821), .A3(n732), .ZN(n581) );
  INVD1 U338 ( .I(n749), .ZN(n831) );
  ND2D1 U339 ( .A1(n850), .A2(n834), .ZN(n642) );
  INVD1 U340 ( .I(n692), .ZN(n833) );
  NR2D1 U341 ( .A1(n711), .A2(n714), .ZN(n722) );
  INVD1 U342 ( .I(n683), .ZN(n820) );
  INVD1 U343 ( .I(n515), .ZN(n837) );
  INVD1 U344 ( .I(n648), .ZN(n818) );
  INVD1 U345 ( .I(n731), .ZN(n808) );
  INVD1 U346 ( .I(n708), .ZN(n827) );
  NR4D0 U347 ( .A1(n635), .A2(n634), .A3(n851), .A4(n633), .ZN(n636) );
  OAI222D0 U348 ( .A1(n443), .A2(n657), .B1(n656), .B2(n787), .C1(n655), .C2(
        n786), .ZN(n658) );
  AOI21D1 U349 ( .A1(n71), .A2(n654), .B(n653), .ZN(n657) );
  OAI222D0 U350 ( .A1(n779), .A2(n788), .B1(n778), .B2(n777), .C1(n776), .C2(
        n775), .ZN(n780) );
  OAI222D0 U351 ( .A1(n580), .A2(n777), .B1(n786), .B2(n579), .C1(n578), .C2(
        n779), .ZN(n583) );
  OAI211D1 U352 ( .A1(n707), .A2(n683), .B(n554), .C(n553), .ZN(n570) );
  OAI211D1 U353 ( .A1(n558), .A2(n425), .B(n557), .C(n556), .ZN(n569) );
  AOI221D0 U354 ( .A1(n807), .A2(n542), .B1(n847), .B2(n541), .C(n540), .ZN(
        n543) );
  INVD1 U355 ( .I(n770), .ZN(n842) );
  NR3D0 U356 ( .A1(n741), .A2(n444), .A3(n768), .ZN(n536) );
  OAI222D0 U357 ( .A1(n519), .A2(n746), .B1(n518), .B2(n753), .C1(n517), .C2(
        n766), .ZN(n523) );
  NR2D1 U358 ( .A1(n862), .A2(n516), .ZN(n517) );
  OAI31D1 U359 ( .A1(n709), .A2(n446), .A3(n449), .B(n643), .ZN(n561) );
  OAI222D0 U360 ( .A1(n624), .A2(n777), .B1(n623), .B2(n726), .C1(n622), .C2(
        n758), .ZN(n625) );
  NR2D1 U361 ( .A1(n811), .A2(n444), .ZN(n623) );
  OA22D0 U362 ( .A1(n779), .A2(n746), .B1(n730), .B2(n621), .Z(n622) );
  OAI222D0 U363 ( .A1(n760), .A2(n632), .B1(n444), .B2(n631), .C1(n754), .C2(
        n771), .ZN(n635) );
  NR2D1 U364 ( .A1(n444), .A2(n446), .ZN(n688) );
  OAI222D0 U365 ( .A1(n733), .A2(n723), .B1(n702), .B2(n448), .C1(n701), .C2(
        n776), .ZN(n703) );
  OAI221D0 U366 ( .A1(n621), .A2(n768), .B1(n753), .B2(n763), .C(n500), .ZN(
        n503) );
  NR4D0 U367 ( .A1(n772), .A2(n760), .A3(n671), .A4(n444), .ZN(n742) );
  ND2D1 U368 ( .A1(n444), .A2(n446), .ZN(n692) );
  CKND1 U369 ( .I(n670), .ZN(n848) );
  OAI221D0 U370 ( .A1(n457), .A2(n648), .B1(n775), .B2(n734), .C(n456), .ZN(
        n463) );
  NR4D0 U371 ( .A1(n510), .A2(n509), .A3(n525), .A4(n526), .ZN(n511) );
  OAI222D0 U372 ( .A1(n766), .A2(n765), .B1(n764), .B2(n763), .C1(n449), .C2(
        n762), .ZN(n791) );
  OAI222D0 U373 ( .A1(n761), .A2(n760), .B1(n759), .B2(n758), .C1(n442), .C2(
        n757), .ZN(n792) );
  NR3D0 U374 ( .A1(n741), .A2(n445), .A3(n616), .ZN(n653) );
  NR4D0 U375 ( .A1(n460), .A2(n459), .A3(n535), .A4(n458), .ZN(n461) );
  ND2D1 U376 ( .A1(n444), .A2(n443), .ZN(n648) );
  OAI222D0 U377 ( .A1(n449), .A2(n779), .B1(n747), .B2(n760), .C1(n754), .C2(
        n750), .ZN(n492) );
  NR4D0 U378 ( .A1(n442), .A2(n836), .A3(n772), .A4(n778), .ZN(n582) );
  NR3D0 U379 ( .A1(n778), .A2(n447), .A3(n445), .ZN(n674) );
  NR3D0 U380 ( .A1(n448), .A2(n445), .A3(n692), .ZN(n600) );
  ND2D1 U381 ( .A1(n442), .A2(n443), .ZN(n763) );
  ND2D1 U382 ( .A1(n445), .A2(n829), .ZN(n617) );
  OAI221D0 U383 ( .A1(n741), .A2(n730), .B1(n450), .B2(n786), .C(n729), .ZN(
        n736) );
  ND2D1 U384 ( .A1(n446), .A2(n815), .ZN(n771) );
  NR2D1 U385 ( .A1(n762), .A2(n442), .ZN(n716) );
  ND2D1 U386 ( .A1(n443), .A2(n452), .ZN(n671) );
  OAI222D0 U387 ( .A1(n508), .A2(n747), .B1(n821), .B2(n507), .C1(n506), .C2(
        n425), .ZN(n510) );
  ND2D1 U388 ( .A1(n447), .A2(n504), .ZN(n507) );
  ND2D1 U389 ( .A1(n443), .A2(n446), .ZN(n748) );
  NR3D0 U390 ( .A1(n723), .A2(n445), .A3(n841), .ZN(n664) );
  ND2D1 U391 ( .A1(n445), .A2(n444), .ZN(n753) );
  ND2D1 U392 ( .A1(n446), .A2(n447), .ZN(n707) );
  AOI221D0 U393 ( .A1(n71), .A2(n816), .B1(n803), .B2(n831), .C(n600), .ZN(
        n601) );
  AOI222D0 U394 ( .A1(n804), .A2(n823), .B1(n825), .B2(n806), .C1(n808), .C2(
        n446), .ZN(n602) );
  INVD1 U395 ( .I(n776), .ZN(n839) );
  ND2D1 U396 ( .A1(n446), .A2(n836), .ZN(n515) );
  ND2D1 U397 ( .A1(n445), .A2(n443), .ZN(n708) );
  OAI221D0 U398 ( .A1(n753), .A2(n755), .B1(n714), .B2(n788), .C(n640), .ZN(
        n651) );
  OAI222D0 U399 ( .A1(n479), .A2(n711), .B1(n472), .B2(n709), .C1(n730), .C2(
        n731), .ZN(n476) );
  AOI221D0 U400 ( .A1(n837), .A2(n71), .B1(n598), .B2(n451), .C(n737), .ZN(
        n599) );
  OAI221D0 U401 ( .A1(n448), .A2(n734), .B1(n709), .B2(n425), .C(n698), .ZN(
        n704) );
  INVD1 U402 ( .I(a[1]), .ZN(n452) );
  IAO21D1 U403 ( .A1(n771), .A2(n783), .B(n853), .ZN(n672) );
  INVD1 U404 ( .I(n771), .ZN(n835) );
  ND2D1 U405 ( .A1(n677), .A2(n861), .ZN(n777) );
  ND2D1 U406 ( .A1(n844), .A2(n677), .ZN(n734) );
  NR2D1 U407 ( .A1(n821), .A2(n829), .ZN(n677) );
  OAI222D0 U408 ( .A1(n447), .A2(n774), .B1(n773), .B2(n772), .C1(n783), .C2(
        n771), .ZN(n781) );
  NR4D0 U409 ( .A1(n692), .A2(n755), .A3(n783), .A4(n821), .ZN(n663) );
  OA222D0 U410 ( .A1(n755), .A2(n764), .B1(n696), .B2(n724), .C1(n695), .C2(
        n783), .Z(n438) );
  INVD1 U411 ( .I(n641), .ZN(n858) );
  NR4D0 U412 ( .A1(n450), .A2(n841), .A3(n766), .A4(n758), .ZN(n700) );
  CKND2D1 U413 ( .A1(n448), .A2(n801), .ZN(n766) );
  INVD0 U414 ( .I(n766), .ZN(n806) );
  NR4D0 U415 ( .A1(n714), .A2(n766), .A3(n760), .A4(n829), .ZN(n738) );
  ND2D0 U416 ( .A1(n766), .A2(n763), .ZN(n751) );
  OA21D1 U417 ( .A1(n833), .A2(n834), .B(n65), .Z(n687) );
  OAI33D0 U418 ( .A1(n662), .A2(n442), .A3(n801), .B1(n490), .B2(n730), .B3(
        n763), .ZN(n491) );
  OAI33D0 U419 ( .A1(n758), .A2(n801), .A3(n730), .B1(n662), .B2(n449), .B3(
        n661), .ZN(n665) );
  OAI222D0 U420 ( .A1(n642), .A2(n801), .B1(n616), .B2(n609), .C1(n444), .C2(
        n724), .ZN(n614) );
  OAI222D0 U421 ( .A1(n755), .A2(n612), .B1(n611), .B2(n801), .C1(n610), .C2(
        n682), .ZN(n613) );
  OAI33D0 U422 ( .A1(n648), .A2(n447), .A3(n772), .B1(n707), .B2(n801), .B3(
        n753), .ZN(n540) );
  CKND2D0 U423 ( .A1(n445), .A2(n801), .ZN(n590) );
  CKND2D0 U424 ( .A1(n801), .A2(n821), .ZN(n558) );
  NR2D1 U425 ( .A1(n470), .A2(n752), .ZN(n439) );
  NR2D0 U426 ( .A1(n469), .A2(n448), .ZN(n441) );
  OAI221D0 U427 ( .A1(n465), .A2(n778), .B1(n724), .B2(n775), .C(n571), .ZN(
        n471) );
  INVD1 U428 ( .I(n604), .ZN(n828) );
  INVD1 U429 ( .I(n662), .ZN(n838) );
  ND2D1 U430 ( .A1(n800), .A2(n861), .ZN(n520) );
  AN2XD1 U431 ( .A1(n442), .A2(n815), .Z(n678) );
  OA21D0 U432 ( .A1(n691), .A2(n448), .B(n620), .Z(n624) );
  AOI21D0 U433 ( .A1(n617), .A2(n662), .B(n691), .ZN(n505) );
  OAI22D0 U434 ( .A1(n768), .A2(n691), .B1(n696), .B2(n714), .ZN(n459) );
  NR3D0 U435 ( .A1(n515), .A2(n753), .A3(n788), .ZN(n481) );
  OAI22D0 U436 ( .A1(n788), .A2(n787), .B1(n786), .B2(n785), .ZN(n789) );
  OAI22D0 U437 ( .A1(n749), .A2(n755), .B1(n768), .B2(n788), .ZN(n693) );
  AOI22D0 U438 ( .A1(n810), .A2(n860), .B1(n802), .B2(n839), .ZN(n574) );
  AOI22D0 U439 ( .A1(n840), .A2(n807), .B1(n810), .B2(n839), .ZN(n474) );
  OAI33D0 U440 ( .A1(n755), .A2(n754), .A3(n753), .B1(n776), .B2(n801), .B3(
        n752), .ZN(n756) );
  OAI222D0 U441 ( .A1(n728), .A2(n433), .B1(n727), .B2(n726), .C1(n725), .C2(
        n724), .ZN(n796) );
  OAI222D0 U442 ( .A1(n730), .A2(n604), .B1(n433), .B2(n765), .C1(n620), .C2(
        n603), .ZN(n605) );
  OAI222D0 U443 ( .A1(n433), .A2(n603), .B1(n734), .B2(n683), .C1(n642), .C2(
        n763), .ZN(n551) );
  CKND2D0 U444 ( .A1(n433), .A2(n755), .ZN(n530) );
  NR3D0 U445 ( .A1(n829), .A2(n450), .A3(n433), .ZN(n535) );
  NR3D0 U446 ( .A1(n678), .A2(n802), .A3(n817), .ZN(n655) );
  CKND2D0 U447 ( .A1(n449), .A2(a[6]), .ZN(n490) );
  CKND2D0 U448 ( .A1(n446), .A2(a[6]), .ZN(n779) );
  CKND2D1 U449 ( .A1(a[6]), .A2(n829), .ZN(n776) );
  AOI31D0 U450 ( .A1(n443), .A2(n829), .A3(n799), .B(n828), .ZN(n500) );
  AOI22D0 U451 ( .A1(n827), .A2(n798), .B1(n825), .B2(n443), .ZN(n578) );
  AOI21D0 U452 ( .A1(n733), .A2(n676), .B(n443), .ZN(n634) );
  AOI221D1 U453 ( .A1(n847), .A2(n464), .B1(n463), .B2(n448), .C(n462), .ZN(
        n486) );
  NR2D1 U454 ( .A1(n805), .A2(n808), .ZN(n580) );
  OAI31D0 U455 ( .A1(n815), .A2(n805), .A3(n811), .B(n697), .ZN(n496) );
  OAI32D1 U456 ( .A1(n771), .A2(n479), .A3(n709), .B1(n478), .B2(n741), .ZN(
        n482) );
  NR4D0 U457 ( .A1(a[6]), .A2(n815), .A3(n730), .A4(n763), .ZN(n509) );
  OA33D0 U458 ( .A1(n711), .A2(n753), .A3(n746), .B1(n710), .B2(n709), .B3(
        n771), .Z(n712) );
  NR3D0 U459 ( .A1(n709), .A2(n829), .A3(n714), .ZN(n527) );
  OAI22D0 U460 ( .A1(a[6]), .A2(n445), .B1(n446), .B2(n760), .ZN(n552) );
endmodule


module aes_sbox_9 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n14, n53, n64, n65, n70, n142, n187, n223, n224, n235, n244, n245,
         n277, n410, n412, n413, n414, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864;

  AN2XD1 U28 ( .A1(n724), .A2(n723), .Z(n728) );
  OA21D1 U35 ( .A1(n708), .A2(n707), .B(n706), .Z(n713) );
  OR4D1 U199 ( .A1(n661), .A2(n585), .A3(n529), .A4(n528), .Z(n531) );
  AN2XD1 U215 ( .A1(n530), .A2(n812), .Z(n529) );
  AN2XD1 U271 ( .A1(n543), .A2(n735), .Z(n476) );
  INVD1 U1 ( .I(n750), .ZN(n831) );
  ND2D1 U2 ( .A1(n451), .A2(n829), .ZN(n750) );
  NR2XD0 U3 ( .A1(n782), .A2(n781), .ZN(n783) );
  INVD3 U4 ( .I(a[1]), .ZN(n457) );
  NR2D2 U5 ( .A1(n142), .A2(n801), .ZN(n694) );
  NR2D1 U6 ( .A1(n810), .A2(n799), .ZN(n623) );
  OAI222D1 U7 ( .A1(n756), .A2(n765), .B1(n694), .B2(n725), .C1(n693), .C2(
        n784), .ZN(n695) );
  OAI222D0 U8 ( .A1(n441), .A2(n753), .B1(n694), .B2(n690), .C1(n759), .C2(
        n563), .ZN(n541) );
  AOI221D1 U9 ( .A1(n470), .A2(n810), .B1(n853), .B2(n819), .C(n469), .ZN(n471) );
  AO31D0 U10 ( .A1(n805), .A2(n860), .A3(n686), .B(n722), .Z(n469) );
  INVD2 U11 ( .I(n734), .ZN(n853) );
  OAI22D0 U12 ( .A1(n70), .A2(n689), .B1(n694), .B2(n714), .ZN(n465) );
  INVD2 U13 ( .I(n689), .ZN(n816) );
  IAO22D0 U14 ( .B1(n858), .B2(n815), .A1(n633), .A2(n777), .ZN(n522) );
  ND2D1 U15 ( .A1(a[6]), .A2(n829), .ZN(n777) );
  AOI221XD4 U16 ( .A1(n849), .A2(n455), .B1(n858), .B2(n437), .C(n646), .ZN(
        n647) );
  AOI221D2 U17 ( .A1(n438), .A2(n826), .B1(n811), .B2(n833), .C(n770), .ZN(
        n785) );
  IIND4D4 U18 ( .A1(n53), .A2(n14), .B1(n631), .B2(n630), .ZN(d[3]) );
  AO221D1 U19 ( .A1(n817), .A2(n610), .B1(n844), .B2(n609), .C(n608), .Z(n14)
         );
  INVD1 U20 ( .I(n690), .ZN(n833) );
  OA222D1 U21 ( .A1(n648), .A2(n641), .B1(n600), .B2(n599), .C1(n598), .C2(
        n761), .Z(n187) );
  INVD2 U22 ( .I(n755), .ZN(n847) );
  INVD1 U23 ( .I(n787), .ZN(n849) );
  OAI31D2 U24 ( .A1(n676), .A2(n142), .A3(n820), .B(n675), .ZN(n677) );
  AOI221D4 U25 ( .A1(n847), .A2(n618), .B1(n617), .B2(n455), .C(n616), .ZN(
        n631) );
  OAI222D1 U26 ( .A1(n756), .A2(n615), .B1(n614), .B2(n803), .C1(n613), .C2(
        n681), .ZN(n616) );
  OAI221D2 U27 ( .A1(n566), .A2(n638), .B1(n723), .B2(n788), .C(n187), .ZN(n53) );
  INVD4 U29 ( .I(n453), .ZN(n829) );
  OAI22D2 U30 ( .A1(n748), .A2(n711), .B1(n645), .B2(n742), .ZN(n646) );
  AOI221D2 U31 ( .A1(n838), .A2(n826), .B1(n824), .B2(n581), .C(n852), .ZN(
        n504) );
  OAI221D1 U32 ( .A1(n742), .A2(n735), .B1(n709), .B2(n748), .C(n602), .ZN(
        n610) );
  IND4D2 U33 ( .A1(n797), .B1(n796), .B2(n795), .B3(n794), .ZN(d[0]) );
  ND4D3 U34 ( .A1(n721), .A2(n720), .A3(n719), .A4(n718), .ZN(d[1]) );
  INVD2 U36 ( .I(n769), .ZN(n64) );
  CKND2 U37 ( .I(n64), .ZN(n65) );
  CKND2 U38 ( .I(n64), .ZN(n70) );
  AOI211XD2 U39 ( .A1(n831), .A2(n597), .B(n595), .C(n596), .ZN(n598) );
  OAI32D2 U40 ( .A1(n594), .A2(n748), .A3(n690), .B1(n593), .B2(n70), .ZN(n595) );
  AOI21D2 U41 ( .A1(n816), .A2(n436), .B(n442), .ZN(n593) );
  INVD2 U42 ( .I(n65), .ZN(n834) );
  CKND2D1 U43 ( .A1(n453), .A2(n815), .ZN(n772) );
  INVD6 U44 ( .I(n451), .ZN(n815) );
  ND2D1 U45 ( .A1(a[6]), .A2(n841), .ZN(n784) );
  ND2D1 U46 ( .A1(n452), .A2(n815), .ZN(n714) );
  ND2D1 U47 ( .A1(n452), .A2(n451), .ZN(n754) );
  ND2D1 U48 ( .A1(n454), .A2(n836), .ZN(n761) );
  CKND2D1 U49 ( .A1(n803), .A2(n815), .ZN(n689) );
  ND2D0 U50 ( .A1(n815), .A2(n821), .ZN(n759) );
  OAI222D0 U51 ( .A1(n454), .A2(n775), .B1(n774), .B2(n773), .C1(n784), .C2(
        n772), .ZN(n782) );
  INVD1 U52 ( .I(n606), .ZN(n852) );
  BUFFD2 U53 ( .I(a[5]), .Z(n453) );
  ND2D1 U54 ( .A1(n453), .A2(n821), .ZN(n769) );
  ND2D1 U55 ( .A1(n451), .A2(n453), .ZN(n690) );
  CKND2D1 U56 ( .A1(n805), .A2(n455), .ZN(n563) );
  INVD1 U57 ( .I(n669), .ZN(n808) );
  INVD1 U58 ( .I(n751), .ZN(n810) );
  BUFFD2 U59 ( .I(a[4]), .Z(n452) );
  INVD1 U60 ( .I(n660), .ZN(n838) );
  INVD1 U61 ( .I(n777), .ZN(n839) );
  AN2XD1 U62 ( .A1(n458), .A2(n803), .Z(n438) );
  ND2D1 U63 ( .A1(n451), .A2(n821), .ZN(n753) );
  INVD2 U64 ( .I(n789), .ZN(n805) );
  ND2D1 U65 ( .A1(n458), .A2(n803), .ZN(n756) );
  INVD4 U66 ( .I(n452), .ZN(n821) );
  NR3D1 U67 ( .A1(n244), .A2(n245), .A3(n572), .ZN(n590) );
  ND4D2 U68 ( .A1(n489), .A2(n488), .A3(n487), .A4(n486), .ZN(d[7]) );
  ND3D1 U69 ( .A1(n427), .A2(n428), .A3(n429), .ZN(n791) );
  AOI21D1 U70 ( .A1(n835), .A2(n844), .B(n852), .ZN(n670) );
  OAI221D0 U71 ( .A1(n689), .A2(n679), .B1(n678), .B2(n789), .C(n677), .ZN(
        n680) );
  NR2D1 U72 ( .A1(n455), .A2(n451), .ZN(n676) );
  NR2D1 U73 ( .A1(n821), .A2(n829), .ZN(n675) );
  OAI222D0 U74 ( .A1(n441), .A2(n543), .B1(n497), .B2(n755), .C1(n496), .C2(
        n759), .ZN(n501) );
  INVD1 U75 ( .I(n779), .ZN(n817) );
  OAI221D0 U76 ( .A1(n742), .A2(n689), .B1(n750), .B2(n708), .C(n688), .ZN(
        n696) );
  INVD1 U77 ( .I(n784), .ZN(n844) );
  OAI222D0 U78 ( .A1(n813), .A2(n638), .B1(n563), .B2(n543), .C1(n542), .C2(
        n784), .ZN(n549) );
  NR4D0 U79 ( .A1(n541), .A2(n540), .A3(n539), .A4(n603), .ZN(n542) );
  NR4D0 U80 ( .A1(n466), .A2(n465), .A3(n539), .A4(n464), .ZN(n467) );
  ND2D1 U81 ( .A1(n836), .A2(n841), .ZN(n755) );
  NR3D1 U82 ( .A1(n431), .A2(n432), .A3(n473), .ZN(n488) );
  ND3D1 U83 ( .A1(n433), .A2(n434), .A3(n435), .ZN(n473) );
  AOI21D1 U84 ( .A1(n862), .A2(n818), .B(n856), .ZN(n576) );
  ND2D1 U85 ( .A1(n451), .A2(n803), .ZN(n776) );
  AN2XD1 U86 ( .A1(n449), .A2(n803), .Z(n142) );
  INVD3 U87 ( .I(n450), .ZN(n803) );
  CKBD4 U88 ( .I(n798), .Z(n455) );
  AOI221D2 U89 ( .A1(n824), .A2(n800), .B1(n833), .B2(n810), .C(n568), .ZN(
        n569) );
  ND2D1 U90 ( .A1(n449), .A2(n457), .ZN(n747) );
  AOI221D1 U91 ( .A1(n808), .A2(n546), .B1(n847), .B2(n545), .C(n544), .ZN(
        n547) );
  ND2D0 U92 ( .A1(n453), .A2(n841), .ZN(n711) );
  INR4D1 U93 ( .A1(n674), .B1(n856), .B2(n672), .B3(n673), .ZN(n684) );
  OAI221D1 U94 ( .A1(n671), .A2(n682), .B1(n670), .B2(n669), .C(n848), .ZN(
        n673) );
  OA222D1 U95 ( .A1(n449), .A2(n684), .B1(n683), .B2(n755), .C1(n682), .C2(
        n681), .Z(n448) );
  ND2D1 U96 ( .A1(n456), .A2(n449), .ZN(n723) );
  CKND1 U97 ( .I(n457), .ZN(n456) );
  ND2D1 U98 ( .A1(n454), .A2(n829), .ZN(n731) );
  CKND0 U99 ( .I(n731), .ZN(n859) );
  OA221D1 U100 ( .A1(n756), .A2(n731), .B1(n764), .B2(n777), .C(n443), .Z(n472) );
  OR2XD1 U101 ( .A1(n570), .A2(n689), .Z(n410) );
  AOI221D2 U102 ( .A1(n814), .A2(n581), .B1(n580), .B2(n824), .C(n579), .ZN(
        n589) );
  NR2XD1 U103 ( .A1(n839), .A2(n850), .ZN(n645) );
  ND2D0 U104 ( .A1(n777), .A2(n731), .ZN(n581) );
  AOI21D0 U105 ( .A1(n801), .A2(n837), .B(n738), .ZN(n443) );
  ND4D3 U106 ( .A1(n589), .A2(n590), .A3(n591), .A4(n588), .ZN(d[4]) );
  ND4D1 U107 ( .A1(n515), .A2(n516), .A3(n517), .A4(n514), .ZN(d[6]) );
  CKND2D1 U108 ( .A1(n829), .A2(n836), .ZN(n660) );
  OAI211D0 U109 ( .A1(n829), .A2(n759), .B(n776), .C(n754), .ZN(n687) );
  OA222D1 U110 ( .A1(n649), .A2(n648), .B1(n764), .B2(n766), .C1(n647), .C2(
        n776), .Z(n446) );
  ND2D2 U111 ( .A1(n853), .A2(n455), .ZN(n643) );
  OA221D0 U112 ( .A1(n755), .A2(n223), .B1(n224), .B2(n449), .C(n235), .Z(n489) );
  OAI222D1 U113 ( .A1(n578), .A2(n714), .B1(n577), .B2(n747), .C1(n437), .C2(
        n576), .ZN(n579) );
  CKND2D1 U114 ( .A1(n450), .A2(n815), .ZN(n779) );
  NR2D0 U115 ( .A1(n835), .A2(n831), .ZN(n678) );
  ND2D1 U116 ( .A1(n430), .A2(n437), .ZN(n592) );
  INVD1 U117 ( .I(n566), .ZN(n804) );
  CKND1 U118 ( .I(n723), .ZN(n799) );
  OA22D0 U119 ( .A1(n467), .A2(n784), .B1(n751), .B2(n641), .Z(n235) );
  ND2D2 U120 ( .A1(n456), .A2(n803), .ZN(n789) );
  NR2D0 U121 ( .A1(n518), .A2(n669), .ZN(n580) );
  ND2D1 U122 ( .A1(n450), .A2(n458), .ZN(n669) );
  OAI22D1 U123 ( .A1(n70), .A2(n779), .B1(n437), .B2(n768), .ZN(n770) );
  INVD1 U124 ( .I(n668), .ZN(n848) );
  OA221D0 U125 ( .A1(n460), .A2(n620), .B1(n779), .B2(n723), .C(n459), .Z(n223) );
  OA221D0 U126 ( .A1(n463), .A2(n648), .B1(n776), .B2(n735), .C(n462), .Z(n224) );
  OAI222D1 U127 ( .A1(n538), .A2(n779), .B1(n441), .B2(n632), .C1(n537), .C2(
        n723), .ZN(n550) );
  CKND2D1 U128 ( .A1(n451), .A2(n458), .ZN(n682) );
  INVD1 U129 ( .I(a[1]), .ZN(n458) );
  AOI22D1 U130 ( .A1(n430), .A2(n834), .B1(n816), .B2(n829), .ZN(n768) );
  NR4D1 U131 ( .A1(n550), .A2(n551), .A3(n549), .A4(n548), .ZN(n552) );
  ND2D2 U132 ( .A1(n437), .A2(n455), .ZN(n742) );
  CKND1 U133 ( .I(n457), .ZN(n437) );
  CKND0 U134 ( .I(n742), .ZN(n802) );
  AOI21D1 U135 ( .A1(n857), .A2(n437), .B(n697), .ZN(n698) );
  OAI22D1 U136 ( .A1(n727), .A2(n756), .B1(n803), .B2(n733), .ZN(n668) );
  OAI222D1 U137 ( .A1(n749), .A2(n723), .B1(n773), .B2(n592), .C1(n754), .C2(
        n764), .ZN(n596) );
  AOI221D1 U138 ( .A1(n801), .A2(n687), .B1(n686), .B2(n808), .C(n685), .ZN(
        n688) );
  AOI221D1 U139 ( .A1(n802), .A2(n692), .B1(n835), .B2(n142), .C(n691), .ZN(
        n693) );
  AOI211XD0 U140 ( .A1(n845), .A2(n449), .B(n644), .C(n854), .ZN(n649) );
  CKND2D2 U141 ( .A1(n455), .A2(n457), .ZN(n748) );
  AOI221D1 U142 ( .A1(n697), .A2(n748), .B1(a[1]), .B2(n855), .C(n565), .ZN(
        n570) );
  AOI221D1 U143 ( .A1(n837), .A2(n799), .B1(n601), .B2(n457), .C(n738), .ZN(
        n602) );
  OAI222D1 U144 ( .A1(n734), .A2(n724), .B1(n702), .B2(n455), .C1(n701), .C2(
        n777), .ZN(n703) );
  AOI221D1 U145 ( .A1(n480), .A2(n457), .B1(n823), .B2(n479), .C(n478), .ZN(
        n487) );
  AOI222D1 U146 ( .A1(n805), .A2(n823), .B1(n825), .B2(n807), .C1(n809), .C2(
        n453), .ZN(n605) );
  AOI221D1 U147 ( .A1(n844), .A2(n658), .B1(n847), .B2(n657), .C(n656), .ZN(
        n665) );
  OAI22D1 U148 ( .A1(n477), .A2(n714), .B1(n476), .B2(n764), .ZN(n478) );
  AOI221D1 U149 ( .A1(n824), .A2(n860), .B1(n430), .B2(n834), .C(n536), .ZN(
        n537) );
  CKAN2D1 U150 ( .A1(n449), .A2(n574), .Z(n244) );
  CKAN2D1 U151 ( .A1(n844), .A2(n573), .Z(n245) );
  OR2D0 U152 ( .A1(n571), .A2(n761), .Z(n277) );
  OR2XD1 U153 ( .A1(n569), .A2(n755), .Z(n412) );
  ND3D2 U154 ( .A1(n277), .A2(n410), .A3(n412), .ZN(n572) );
  OAI211D0 U155 ( .A1(n562), .A2(n723), .B(n561), .C(n560), .ZN(n573) );
  OA221D1 U156 ( .A1(n638), .A2(n764), .B1(n447), .B2(n789), .C(n448), .Z(n721) );
  INVD3 U157 ( .I(n454), .ZN(n841) );
  ND2D1 U158 ( .A1(n832), .A2(n844), .ZN(n727) );
  AOI221D1 U159 ( .A1(n844), .A2(n506), .B1(n804), .B2(n519), .C(n505), .ZN(
        n515) );
  AOI221D1 U160 ( .A1(n705), .A2(n859), .B1(n818), .B2(n704), .C(n703), .ZN(
        n719) );
  ND2D0 U161 ( .A1(n803), .A2(n821), .ZN(n562) );
  AOI221D1 U162 ( .A1(n857), .A2(n799), .B1(n696), .B2(n860), .C(n695), .ZN(
        n720) );
  OR2D0 U163 ( .A1(n669), .A2(n772), .Z(n413) );
  OR2XD1 U164 ( .A1(n449), .A2(n567), .Z(n414) );
  OR2D0 U165 ( .A1(n754), .A2(n566), .Z(n424) );
  ND3D2 U166 ( .A1(n413), .A2(n414), .A3(n424), .ZN(n568) );
  AOI22D1 U167 ( .A1(n832), .A2(n818), .B1(n808), .B2(n829), .ZN(n567) );
  CKAN2D1 U168 ( .A1(n861), .A2(n455), .Z(n425) );
  CKAN2D1 U169 ( .A1(n853), .A2(n810), .Z(n426) );
  NR3D0 U170 ( .A1(n425), .A2(n426), .A3(n639), .ZN(n667) );
  ND4D2 U171 ( .A1(n667), .A2(n666), .A3(n665), .A4(n664), .ZN(d[2]) );
  OR2XD1 U172 ( .A1(n785), .A2(n784), .Z(n427) );
  OR2D0 U173 ( .A1(n451), .A2(n842), .Z(n428) );
  OR2XD1 U174 ( .A1(n783), .A2(n455), .Z(n429) );
  CKND0 U175 ( .I(n771), .ZN(n842) );
  NR4D1 U176 ( .A1(n793), .A2(n792), .A3(n791), .A4(n790), .ZN(n794) );
  AN4D1 U177 ( .A1(n675), .A2(n819), .A3(n449), .A4(n847), .Z(n528) );
  ND2D0 U178 ( .A1(n675), .A2(n850), .ZN(n599) );
  ND3D0 U179 ( .A1(n818), .A2(n675), .A3(n847), .ZN(n763) );
  ND2D1 U180 ( .A1(n844), .A2(n675), .ZN(n735) );
  OAI22D0 U181 ( .A1(n759), .A2(n756), .B1(n659), .B2(n742), .ZN(n527) );
  CKND2D0 U182 ( .A1(n441), .A2(n756), .ZN(n533) );
  CKND2D2 U183 ( .A1(n821), .A2(n829), .ZN(n773) );
  INVD1 U184 ( .I(n776), .ZN(n430) );
  AN2XD1 U185 ( .A1(n437), .A2(n474), .Z(n431) );
  CKAN2D1 U186 ( .A1(n828), .A2(n838), .Z(n432) );
  OR2D0 U187 ( .A1(n472), .A2(n753), .Z(n433) );
  OR2D0 U188 ( .A1(n690), .A2(n523), .Z(n434) );
  OR2D0 U189 ( .A1(n455), .A2(n471), .Z(n435) );
  CKND0 U190 ( .I(n457), .ZN(n436) );
  ND2D0 U191 ( .A1(n837), .A2(n826), .ZN(n543) );
  ND2D1 U192 ( .A1(n850), .A2(n834), .ZN(n642) );
  ND2D1 U193 ( .A1(n831), .A2(n850), .ZN(n606) );
  ND2D1 U194 ( .A1(n454), .A2(a[6]), .ZN(n709) );
  BUFFD4 U195 ( .I(a[7]), .Z(n454) );
  ND2D0 U196 ( .A1(n449), .A2(n803), .ZN(n441) );
  CKAN2D1 U197 ( .A1(n831), .A2(n802), .Z(n439) );
  CKAN2D1 U198 ( .A1(n823), .A2(n808), .Z(n440) );
  NR3D0 U200 ( .A1(n680), .A2(n439), .A3(n440), .ZN(n683) );
  NR2D0 U201 ( .A1(n633), .A2(n723), .ZN(n705) );
  OAI31D0 U202 ( .A1(n709), .A2(n453), .A3(n436), .B(n643), .ZN(n565) );
  OAI211D0 U203 ( .A1(n707), .A2(n682), .B(n558), .C(n557), .ZN(n574) );
  CKND0 U204 ( .I(n643), .ZN(n854) );
  BUFFD4 U205 ( .I(a[0]), .Z(n449) );
  CKND2D0 U206 ( .A1(n430), .A2(n855), .ZN(n575) );
  ND2D0 U207 ( .A1(n802), .A2(n860), .ZN(n523) );
  AOI21D1 U208 ( .A1(n822), .A2(n863), .B(n851), .ZN(n577) );
  CKND2D0 U209 ( .A1(n786), .A2(n689), .ZN(n532) );
  NR2D0 U210 ( .A1(n632), .A2(n747), .ZN(n771) );
  NR2XD0 U211 ( .A1(n861), .A2(n519), .ZN(n520) );
  CKND2D1 U212 ( .A1(n454), .A2(n507), .ZN(n510) );
  CKND0 U213 ( .I(n740), .ZN(n813) );
  CKND2D0 U214 ( .A1(n690), .A2(n753), .ZN(n692) );
  OAI22D0 U216 ( .A1(n750), .A2(n756), .B1(n70), .B2(n789), .ZN(n691) );
  CKND2D0 U217 ( .A1(n436), .A2(a[6]), .ZN(n493) );
  CKND0 U218 ( .I(n778), .ZN(n861) );
  NR2XD0 U219 ( .A1(n845), .A2(n855), .ZN(n671) );
  CKND0 U220 ( .I(n592), .ZN(n814) );
  ND2D0 U221 ( .A1(n847), .A2(n834), .ZN(n787) );
  AOI22D0 U222 ( .A1(n862), .A2(n805), .B1(n819), .B2(n849), .ZN(n557) );
  ND2D0 U223 ( .A1(n817), .A2(n436), .ZN(n724) );
  CKND2D0 U224 ( .A1(n863), .A2(n826), .ZN(n788) );
  ND2D0 U225 ( .A1(n832), .A2(n860), .ZN(n681) );
  ND2D0 U226 ( .A1(n824), .A2(n863), .ZN(n765) );
  CKND2D0 U227 ( .A1(n823), .A2(n847), .ZN(n674) );
  CKND0 U228 ( .I(n725), .ZN(n846) );
  NR2D0 U229 ( .A1(n722), .A2(n858), .ZN(n729) );
  NR2D0 U230 ( .A1(n862), .A2(n849), .ZN(n468) );
  CKND2D0 U231 ( .A1(n832), .A2(n457), .ZN(n679) );
  OAI33D0 U232 ( .A1(n759), .A2(n803), .A3(n731), .B1(n660), .B2(a[1]), .B3(
        n659), .ZN(n663) );
  AOI221D0 U233 ( .A1(n430), .A2(n846), .B1(n853), .B2(n819), .C(n555), .ZN(
        n591) );
  CKND2D0 U234 ( .A1(n786), .A2(n563), .ZN(n564) );
  AOI21D0 U235 ( .A1(n690), .A2(n70), .B(n441), .ZN(n685) );
  AOI22D0 U236 ( .A1(n853), .A2(n533), .B1(n697), .B2(n532), .ZN(n534) );
  OAI32D0 U237 ( .A1(n566), .A2(n761), .A3(n750), .B1(n524), .B2(n523), .ZN(
        n525) );
  NR2D0 U238 ( .A1(n834), .A2(n430), .ZN(n524) );
  CKND2D0 U239 ( .A1(n754), .A2(n749), .ZN(n559) );
  NR2D0 U240 ( .A1(n827), .A2(n832), .ZN(n611) );
  CKND2D0 U241 ( .A1(n767), .A2(n764), .ZN(n752) );
  OAI31D0 U242 ( .A1(n742), .A2(n825), .A3(n755), .B(n741), .ZN(n746) );
  AOI31D0 U243 ( .A1(n850), .A2(n740), .A3(n825), .B(n739), .ZN(n741) );
  NR2D0 U244 ( .A1(n430), .A2(n807), .ZN(n460) );
  ND2D0 U245 ( .A1(n829), .A2(n841), .ZN(n619) );
  OAI21D0 U246 ( .A1(n754), .A2(n619), .B(n641), .ZN(n519) );
  CKND0 U247 ( .I(n754), .ZN(n825) );
  CKND2D0 U248 ( .A1(n810), .A2(n455), .ZN(n710) );
  CKND2D0 U249 ( .A1(n830), .A2(n850), .ZN(n641) );
  AOI31D0 U250 ( .A1(n735), .A2(n734), .A3(n733), .B(n732), .ZN(n736) );
  INR2D0 U251 ( .A1(n530), .B1(n669), .ZN(n715) );
  CKND2D0 U252 ( .A1(n686), .A2(n850), .ZN(n638) );
  OAI21D0 U253 ( .A1(n648), .A2(n734), .B(n788), .ZN(n480) );
  CKND2D0 U254 ( .A1(n732), .A2(n742), .ZN(n597) );
  CKND2D0 U255 ( .A1(n800), .A2(n815), .ZN(n726) );
  CKND0 U256 ( .I(n707), .ZN(n863) );
  CKND2D0 U257 ( .A1(n833), .A2(n850), .ZN(n766) );
  ND2D0 U258 ( .A1(n834), .A2(n841), .ZN(n632) );
  CKND2D0 U259 ( .A1(n824), .A2(n850), .ZN(n615) );
  OAI31D0 U260 ( .A1(n815), .A2(n806), .A3(n812), .B(n697), .ZN(n499) );
  CKND2D1 U261 ( .A1(n499), .A2(n498), .ZN(n500) );
  ND2D0 U262 ( .A1(n455), .A2(n803), .ZN(n767) );
  AOI21D0 U263 ( .A1(n451), .A2(n860), .B(n820), .ZN(n774) );
  AOI22D0 U264 ( .A1(n805), .A2(n838), .B1(n430), .B2(n821), .ZN(n775) );
  AOI22D0 U265 ( .A1(n810), .A2(n449), .B1(n436), .B2(n818), .ZN(n491) );
  NR2D0 U266 ( .A1(n812), .A2(n810), .ZN(n475) );
  OAI21D0 U267 ( .A1(n660), .A2(n753), .B(n733), .ZN(n546) );
  OAI33D0 U268 ( .A1(n648), .A2(n454), .A3(n773), .B1(n707), .B2(n803), .B3(
        n754), .ZN(n544) );
  AOI21D0 U269 ( .A1(n689), .A2(n594), .B(n747), .ZN(n464) );
  AOI21D0 U270 ( .A1(n824), .A2(n859), .B(n699), .ZN(n511) );
  AOI211XD0 U272 ( .A1(n843), .A2(n811), .B(n495), .C(n494), .ZN(n496) );
  CKND0 U273 ( .I(n619), .ZN(n843) );
  NR2D0 U274 ( .A1(n806), .A2(n809), .ZN(n584) );
  CKND2D0 U275 ( .A1(n723), .A2(n815), .ZN(n583) );
  OAI21D0 U276 ( .A1(n755), .A2(n620), .B(n725), .ZN(n601) );
  CKND2D0 U277 ( .A1(n818), .A2(n821), .ZN(n612) );
  NR2XD0 U278 ( .A1(n651), .A2(n771), .ZN(n614) );
  AOI211D0 U279 ( .A1(n820), .A2(n449), .B(n818), .C(n812), .ZN(n613) );
  ND4D0 U280 ( .A1(n801), .A2(n838), .A3(n452), .A4(n454), .ZN(n730) );
  OAI22D0 U281 ( .A1(n789), .A2(n788), .B1(n787), .B2(n786), .ZN(n790) );
  OAI32D0 U282 ( .A1(n772), .A2(n482), .A3(n709), .B1(n481), .B2(n742), .ZN(
        n485) );
  AOI31D0 U283 ( .A1(n452), .A2(n836), .A3(n430), .B(n699), .ZN(n481) );
  OAI22D0 U284 ( .A1(n454), .A2(n660), .B1(n754), .B2(n731), .ZN(n461) );
  NR2D0 U285 ( .A1(n858), .A2(n697), .ZN(n463) );
  OAI22D0 U286 ( .A1(n458), .A2(n725), .B1(n437), .B2(n642), .ZN(n644) );
  AOI211D0 U287 ( .A1(n780), .A2(n660), .B(n594), .C(n747), .ZN(n483) );
  AOI33D0 U288 ( .A1(n621), .A2(n836), .A3(n805), .B1(n855), .B2(n815), .B3(
        n802), .ZN(n622) );
  OAI31D0 U289 ( .A1(n751), .A2(n780), .A3(n753), .B(n622), .ZN(n629) );
  NR2D0 U290 ( .A1(n734), .A2(n451), .ZN(n699) );
  OAI22D0 U291 ( .A1(n458), .A2(n638), .B1(n637), .B2(n747), .ZN(n639) );
  AOI21D0 U292 ( .A1(n858), .A2(n819), .B(n699), .ZN(n702) );
  OAI211D0 U293 ( .A1(n453), .A2(n786), .B(n633), .C(n753), .ZN(n545) );
  CKND2D0 U294 ( .A1(n449), .A2(n808), .ZN(n732) );
  CKND2D1 U295 ( .A1(n605), .A2(n604), .ZN(n609) );
  OAI21D0 U296 ( .A1(n449), .A2(n690), .B(n753), .ZN(n492) );
  AOI21D0 U297 ( .A1(n849), .A2(n818), .B(n757), .ZN(n758) );
  OAI33D0 U298 ( .A1(n756), .A2(n755), .A3(n754), .B1(n777), .B2(n803), .B3(
        n753), .ZN(n757) );
  CKND2D0 U299 ( .A1(n453), .A2(n836), .ZN(n518) );
  OAI21D0 U300 ( .A1(n713), .A2(n742), .B(n712), .ZN(n717) );
  OA33D0 U301 ( .A1(n711), .A2(n754), .A3(n747), .B1(n710), .B2(n709), .B3(
        n772), .Z(n712) );
  AOI21D0 U302 ( .A1(n809), .A2(n847), .B(n580), .ZN(n521) );
  CKND0 U303 ( .I(n697), .ZN(n447) );
  NR2D0 U304 ( .A1(n452), .A2(n836), .ZN(n470) );
  OAI33D0 U305 ( .A1(n660), .A2(n449), .A3(n803), .B1(n493), .B2(n731), .B3(
        n764), .ZN(n494) );
  CKND2D0 U306 ( .A1(n453), .A2(a[6]), .ZN(n780) );
  AOI32D0 U307 ( .A1(n452), .A2(n841), .A3(n817), .B1(n818), .B2(n556), .ZN(
        n558) );
  OAI22D0 U308 ( .A1(a[6]), .A2(n452), .B1(n453), .B2(n761), .ZN(n556) );
  CKBD4 U309 ( .I(a[3]), .Z(n451) );
  BUFFD4 U310 ( .I(a[2]), .Z(n450) );
  INVD1 U311 ( .I(n681), .ZN(n862) );
  INVD1 U312 ( .I(n788), .ZN(n864) );
  INVD1 U313 ( .I(n575), .ZN(n856) );
  INVD1 U314 ( .I(n607), .ZN(n828) );
  NR2D1 U315 ( .A1(n642), .A2(n726), .ZN(n744) );
  NR2D1 U316 ( .A1(n818), .A2(n825), .ZN(n659) );
  INVD1 U317 ( .I(n599), .ZN(n858) );
  ND2D1 U318 ( .A1(n799), .A2(n827), .ZN(n607) );
  INVD1 U319 ( .I(n642), .ZN(n855) );
  INVD1 U320 ( .I(n727), .ZN(n845) );
  INVD1 U321 ( .I(n767), .ZN(n807) );
  INVD1 U322 ( .I(n759), .ZN(n823) );
  INVD1 U323 ( .I(n710), .ZN(n811) );
  ND2D1 U324 ( .A1(n822), .A2(n838), .ZN(n706) );
  INVD1 U325 ( .I(n562), .ZN(n822) );
  INVD1 U326 ( .I(n615), .ZN(n851) );
  NR2D1 U327 ( .A1(n755), .A2(n773), .ZN(n697) );
  OAI222D0 U328 ( .A1(n441), .A2(n606), .B1(n735), .B2(n682), .C1(n642), .C2(
        n764), .ZN(n555) );
  OAI221D0 U329 ( .A1(n468), .A2(n779), .B1(n725), .B2(n776), .C(n575), .ZN(
        n474) );
  OAI222D0 U330 ( .A1(n764), .A2(n772), .B1(n786), .B2(n650), .C1(n753), .C2(
        n710), .ZN(n658) );
  OAI222D0 U331 ( .A1(n731), .A2(n607), .B1(n441), .B2(n766), .C1(n623), .C2(
        n606), .ZN(n608) );
  OAI222D0 U332 ( .A1(n787), .A2(n592), .B1(n779), .B2(n643), .C1(n504), .C2(
        n767), .ZN(n505) );
  NR4D0 U333 ( .A1(n485), .A2(n484), .A3(n716), .A4(n483), .ZN(n486) );
  OAI222D0 U334 ( .A1(n729), .A2(n441), .B1(n728), .B2(n727), .C1(n726), .C2(
        n725), .ZN(n797) );
  AOI221D0 U335 ( .A1(n738), .A2(n817), .B1(n816), .B2(n737), .C(n736), .ZN(
        n796) );
  NR4D0 U336 ( .A1(n746), .A2(n745), .A3(n744), .A4(n743), .ZN(n795) );
  NR4D0 U337 ( .A1(n587), .A2(n586), .A3(n585), .A4(n743), .ZN(n588) );
  AOI221D0 U338 ( .A1(n806), .A2(n835), .B1(n830), .B2(n564), .C(n705), .ZN(
        n571) );
  INVD1 U339 ( .I(n753), .ZN(n824) );
  NR4D0 U340 ( .A1(n663), .A2(n662), .A3(n661), .A4(n745), .ZN(n664) );
  NR2D1 U341 ( .A1(n629), .A2(n628), .ZN(n630) );
  OAI221D0 U342 ( .A1(n436), .A2(n674), .B1(n726), .B2(n681), .C(n534), .ZN(
        n551) );
  NR3D0 U343 ( .A1(n829), .A2(n437), .A3(n441), .ZN(n539) );
  NR2D1 U344 ( .A1(n707), .A2(n748), .ZN(n738) );
  NR4D0 U345 ( .A1(n717), .A2(n739), .A3(n716), .A4(n715), .ZN(n718) );
  ND3D1 U346 ( .A1(n554), .A2(n553), .A3(n552), .ZN(d[5]) );
  AOI211D1 U347 ( .A1(n863), .A2(n527), .B(n526), .C(n525), .ZN(n554) );
  INR4D0 U348 ( .A1(n763), .B1(n531), .B2(n744), .B3(n715), .ZN(n553) );
  NR3D0 U349 ( .A1(n723), .A2(n821), .A3(n733), .ZN(n585) );
  INVD1 U350 ( .I(n772), .ZN(n835) );
  INVD1 U351 ( .I(n786), .ZN(n819) );
  ND2D1 U352 ( .A1(n686), .A2(n847), .ZN(n733) );
  NR3D0 U353 ( .A1(n518), .A2(n754), .A3(n789), .ZN(n484) );
  ND2D1 U354 ( .A1(n844), .A2(n830), .ZN(n725) );
  ND2D1 U355 ( .A1(n832), .A2(n850), .ZN(n734) );
  INVD1 U356 ( .I(n682), .ZN(n820) );
  NR2D1 U357 ( .A1(n711), .A2(n714), .ZN(n722) );
  NR3D0 U358 ( .A1(n676), .A2(n430), .A3(n458), .ZN(n444) );
  INVD1 U359 ( .I(n620), .ZN(n832) );
  INVD1 U360 ( .I(n648), .ZN(n818) );
  INVD1 U361 ( .I(n518), .ZN(n837) );
  INVD1 U362 ( .I(n761), .ZN(n860) );
  INVD1 U363 ( .I(n708), .ZN(n827) );
  INVD1 U364 ( .I(n747), .ZN(n801) );
  INVD1 U365 ( .I(n732), .ZN(n809) );
  OAI221D0 U366 ( .A1(n455), .A2(n735), .B1(n709), .B2(n723), .C(n698), .ZN(
        n704) );
  OAI222D0 U367 ( .A1(n780), .A2(n789), .B1(n779), .B2(n778), .C1(n777), .C2(
        n776), .ZN(n781) );
  AOI221D0 U368 ( .A1(n799), .A2(n816), .B1(n804), .B2(n831), .C(n603), .ZN(
        n604) );
  OAI222D0 U369 ( .A1(n750), .A2(n563), .B1(n648), .B2(n723), .C1(n751), .C2(
        n690), .ZN(n466) );
  OAI222D0 U370 ( .A1(n710), .A2(n735), .B1(n449), .B2(n547), .C1(n789), .C2(
        n778), .ZN(n548) );
  OAI222D0 U371 ( .A1(n522), .A2(n747), .B1(n521), .B2(n754), .C1(n520), .C2(
        n767), .ZN(n526) );
  AOI222D0 U372 ( .A1(n810), .A2(n832), .B1(n808), .B2(n492), .C1(n804), .C2(
        n835), .ZN(n497) );
  OAI222D0 U373 ( .A1(n627), .A2(n778), .B1(n626), .B2(n727), .C1(n625), .C2(
        n759), .ZN(n628) );
  NR2D1 U374 ( .A1(n812), .A2(n451), .ZN(n626) );
  OA22D0 U375 ( .A1(n780), .A2(n747), .B1(n731), .B2(n624), .Z(n625) );
  AOI221D0 U376 ( .A1(n862), .A2(n457), .B1(n845), .B2(n723), .C(n535), .ZN(
        n538) );
  OAI221D0 U377 ( .A1(n619), .A2(n594), .B1(n451), .B2(n778), .C(n706), .ZN(
        n536) );
  OAI222D0 U378 ( .A1(n584), .A2(n778), .B1(n787), .B2(n583), .C1(n582), .C2(
        n780), .ZN(n587) );
  OAI222D0 U379 ( .A1(n761), .A2(n633), .B1(n451), .B2(n632), .C1(n755), .C2(
        n772), .ZN(n636) );
  OAI222D0 U380 ( .A1(n482), .A2(n711), .B1(n475), .B2(n709), .C1(n731), .C2(
        n732), .ZN(n479) );
  OAI222D0 U381 ( .A1(n642), .A2(n803), .B1(n619), .B2(n612), .C1(n451), .C2(
        n725), .ZN(n617) );
  OAI221D0 U382 ( .A1(n742), .A2(n731), .B1(n437), .B2(n787), .C(n730), .ZN(
        n737) );
  ND2D1 U383 ( .A1(n451), .A2(n450), .ZN(n648) );
  ND2D1 U384 ( .A1(n436), .A2(n451), .ZN(n786) );
  NR4D0 U385 ( .A1(n513), .A2(n512), .A3(n528), .A4(n529), .ZN(n514) );
  AOI211XD0 U386 ( .A1(n860), .A2(n502), .B(n501), .C(n500), .ZN(n516) );
  ND2D1 U387 ( .A1(a[1]), .A2(n450), .ZN(n751) );
  OAI222D0 U388 ( .A1(n767), .A2(n766), .B1(n765), .B2(n764), .C1(n437), .C2(
        n763), .ZN(n792) );
  OAI222D0 U389 ( .A1(n762), .A2(n761), .B1(n760), .B2(n759), .C1(n449), .C2(
        n758), .ZN(n793) );
  NR4D0 U390 ( .A1(n636), .A2(n635), .A3(n851), .A4(n634), .ZN(n637) );
  NR3D0 U391 ( .A1(n742), .A2(n452), .A3(n619), .ZN(n651) );
  ND2D1 U392 ( .A1(n449), .A2(n450), .ZN(n764) );
  NR4D0 U393 ( .A1(n449), .A2(n836), .A3(n773), .A4(n779), .ZN(n586) );
  OAI221D0 U394 ( .A1(n624), .A2(n70), .B1(n754), .B2(n764), .C(n503), .ZN(
        n506) );
  NR2D1 U395 ( .A1(n451), .A2(n453), .ZN(n686) );
  AOI211XD0 U396 ( .A1(n806), .A2(n825), .B(n828), .C(n700), .ZN(n701) );
  NR4D0 U397 ( .A1(n436), .A2(n841), .A3(n767), .A4(n759), .ZN(n700) );
  NR3D0 U398 ( .A1(n742), .A2(n451), .A3(n70), .ZN(n540) );
  ND2D1 U399 ( .A1(n453), .A2(n454), .ZN(n707) );
  NR3D0 U400 ( .A1(n779), .A2(n454), .A3(n452), .ZN(n672) );
  AOI21D1 U401 ( .A1(n799), .A2(n652), .B(n651), .ZN(n655) );
  OAI222D0 U402 ( .A1(n756), .A2(n690), .B1(n491), .B2(n70), .C1(n436), .C2(
        n754), .ZN(n502) );
  NR2D1 U403 ( .A1(n763), .A2(n449), .ZN(n716) );
  NR3D0 U404 ( .A1(n724), .A2(n452), .A3(n841), .ZN(n662) );
  ND2D1 U405 ( .A1(n452), .A2(n803), .ZN(n594) );
  INVD1 U406 ( .I(n709), .ZN(n850) );
  ND2D1 U407 ( .A1(n452), .A2(n829), .ZN(n620) );
  ND2D1 U408 ( .A1(n438), .A2(n449), .ZN(n566) );
  INVD1 U409 ( .I(n449), .ZN(n798) );
  INVD1 U410 ( .I(n780), .ZN(n840) );
  OAI222D0 U411 ( .A1(n437), .A2(n780), .B1(n748), .B2(n761), .C1(n755), .C2(
        n751), .ZN(n495) );
  OAI222D0 U412 ( .A1(n511), .A2(n748), .B1(n821), .B2(n510), .C1(n509), .C2(
        n723), .ZN(n513) );
  INR2D1 U413 ( .A1(n765), .B1(n508), .ZN(n509) );
  NR4D0 U414 ( .A1(a[6]), .A2(n815), .A3(n731), .A4(n764), .ZN(n512) );
  INVD2 U415 ( .I(a[6]), .ZN(n836) );
  ND2D1 U416 ( .A1(n675), .A2(n860), .ZN(n778) );
  ND2D0 U417 ( .A1(n142), .A2(n834), .ZN(n650) );
  NR2D0 U418 ( .A1(n142), .A2(n800), .ZN(n624) );
  AOI222D0 U419 ( .A1(n810), .A2(n826), .B1(n824), .B2(n142), .C1(n833), .C2(
        n808), .ZN(n560) );
  INVD1 U420 ( .I(n563), .ZN(n442) );
  CKND0 U421 ( .I(n563), .ZN(n806) );
  NR3D0 U422 ( .A1(n676), .A2(n438), .A3(n817), .ZN(n653) );
  AO221D0 U423 ( .A1(n438), .A2(n835), .B1(n802), .B2(n817), .C(n705), .Z(n657) );
  AOI22D0 U424 ( .A1(n811), .A2(n859), .B1(n438), .B2(n839), .ZN(n578) );
  OAI31D0 U425 ( .A1(n438), .A2(n801), .A3(n430), .B(n861), .ZN(n498) );
  NR2D1 U426 ( .A1(n807), .A2(n438), .ZN(n482) );
  AOI32D0 U427 ( .A1(n454), .A2(n821), .A3(n438), .B1(n808), .B2(n461), .ZN(
        n462) );
  AOI32D0 U428 ( .A1(n438), .A2(n455), .A3(n835), .B1(n802), .B2(n559), .ZN(
        n561) );
  INVD1 U429 ( .I(n764), .ZN(n812) );
  OA32D0 U430 ( .A1(n829), .A2(n449), .A3(n786), .B1(n773), .B2(n444), .Z(n640) );
  INVD1 U431 ( .I(n773), .ZN(n830) );
  AOI211XD0 U432 ( .A1(n864), .A2(n811), .B(n490), .C(n668), .ZN(n517) );
  ND2D1 U433 ( .A1(n450), .A2(n742), .ZN(n740) );
  OAI222D0 U434 ( .A1(n450), .A2(n655), .B1(n654), .B2(n788), .C1(n653), .C2(
        n787), .ZN(n656) );
  ND2D1 U435 ( .A1(n450), .A2(n453), .ZN(n749) );
  ND2D1 U436 ( .A1(n450), .A2(n821), .ZN(n633) );
  ND2D1 U437 ( .A1(n452), .A2(n450), .ZN(n708) );
  OA221D1 U438 ( .A1(n761), .A2(n445), .B1(n641), .B2(n789), .C(n446), .Z(n666) );
  OA221D0 U439 ( .A1(n754), .A2(n756), .B1(n714), .B2(n789), .C(n640), .Z(n445) );
  INVD1 U440 ( .I(n641), .ZN(n857) );
  OAI22D0 U441 ( .A1(n747), .A2(n759), .B1(n611), .B2(n748), .ZN(n618) );
  NR2D1 U442 ( .A1(n455), .A2(n763), .ZN(n745) );
  OA21D0 U443 ( .A1(n689), .A2(n455), .B(n623), .Z(n627) );
  OAI22D0 U444 ( .A1(n648), .A2(n747), .B1(n748), .B2(n776), .ZN(n507) );
  OA222D0 U445 ( .A1(n751), .A2(n750), .B1(n749), .B2(n748), .C1(n753), .C2(
        n747), .Z(n762) );
  AOI22D0 U446 ( .A1(n455), .A2(n819), .B1(n815), .B2(n807), .ZN(n600) );
  OAI22D0 U447 ( .A1(n455), .A2(n725), .B1(n458), .B2(n735), .ZN(n535) );
  INVD1 U448 ( .I(n748), .ZN(n800) );
  NR3D0 U449 ( .A1(n455), .A2(n452), .A3(n690), .ZN(n603) );
  AOI21D0 U450 ( .A1(n620), .A2(n660), .B(n689), .ZN(n508) );
  OAI22D0 U451 ( .A1(n451), .A2(n620), .B1(n455), .B2(n619), .ZN(n621) );
  NR4D0 U452 ( .A1(n714), .A2(n767), .A3(n761), .A4(n829), .ZN(n739) );
  NR3D0 U453 ( .A1(n709), .A2(n829), .A3(n714), .ZN(n530) );
  OAI22D0 U454 ( .A1(n836), .A2(n714), .B1(n821), .B2(n660), .ZN(n652) );
  INVD1 U455 ( .I(n714), .ZN(n826) );
  NR4D0 U456 ( .A1(n773), .A2(n761), .A3(n669), .A4(n451), .ZN(n743) );
  OAI222D0 U457 ( .A1(n648), .A2(n727), .B1(n600), .B2(n735), .C1(n642), .C2(
        n669), .ZN(n490) );
  AOI22D0 U458 ( .A1(n827), .A2(n800), .B1(n825), .B2(n450), .ZN(n582) );
  AOI31D0 U459 ( .A1(n450), .A2(n829), .A3(n801), .B(n828), .ZN(n503) );
  AOI21D0 U460 ( .A1(n734), .A2(n674), .B(n450), .ZN(n635) );
  AOI22D0 U461 ( .A1(n838), .A2(n752), .B1(n840), .B2(n808), .ZN(n760) );
  AOI22D0 U462 ( .A1(n831), .A2(n808), .B1(n805), .B2(n833), .ZN(n459) );
  AOI22D0 U463 ( .A1(n840), .A2(n808), .B1(n811), .B2(n839), .ZN(n477) );
  NR2D1 U464 ( .A1(n800), .A2(n808), .ZN(n654) );
  AOI21D0 U465 ( .A1(n779), .A2(n749), .B(n784), .ZN(n634) );
  NR4D0 U466 ( .A1(n690), .A2(n756), .A3(n784), .A4(n821), .ZN(n661) );
endmodule


module aes_sbox_8 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n35, n64, n65, n70, n72, n73, n74, n185, n192, n205, n244, n245, n277,
         n310, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856;

  OA21D1 U35 ( .A1(n701), .A2(n700), .B(n699), .Z(n706) );
  OR3D1 U88 ( .A1(n670), .A2(n805), .A3(n447), .Z(n632) );
  OR4D1 U199 ( .A1(n656), .A2(n577), .A3(n522), .A4(n521), .Z(n524) );
  MAOI22D1 U209 ( .A1(n850), .A2(n277), .B1(n625), .B2(n771), .ZN(n515) );
  AN2XD1 U215 ( .A1(n523), .A2(n803), .Z(n522) );
  AN2XD1 U271 ( .A1(n536), .A2(n729), .Z(n469) );
  AO31D1 U286 ( .A1(n796), .A2(n852), .A3(n429), .B(n715), .Z(n462) );
  AO21D1 U297 ( .A1(n792), .A2(n828), .B(n732), .Z(n461) );
  OAI222D1 U1 ( .A1(n728), .A2(n717), .B1(n695), .B2(n443), .C1(n694), .C2(
        n771), .ZN(n696) );
  AOI211D1 U2 ( .A1(n797), .A2(n817), .B(n820), .C(n693), .ZN(n694) );
  AOI211XD1 U3 ( .A1(n852), .A2(n495), .B(n494), .C(n493), .ZN(n509) );
  INVD2 U4 ( .I(n682), .ZN(n808) );
  INVD2 U5 ( .I(n663), .ZN(n799) );
  AOI222D1 U6 ( .A1(n796), .A2(n815), .B1(n817), .B2(n798), .C1(n800), .C2(
        n441), .ZN(n597) );
  ND2D2 U7 ( .A1(n823), .A2(n841), .ZN(n728) );
  INVD2 U8 ( .I(n702), .ZN(n841) );
  CKND2D1 U9 ( .A1(n433), .A2(n841), .ZN(n598) );
  CKND2D1 U10 ( .A1(n841), .A2(n825), .ZN(n635) );
  ND4D2 U11 ( .A1(n481), .A2(n480), .A3(n482), .A4(n479), .ZN(d[7]) );
  INVD2 U12 ( .I(n439), .ZN(n807) );
  NR4D1 U13 ( .A1(n628), .A2(n627), .A3(n842), .A4(n626), .ZN(n629) );
  AOI211XD1 U14 ( .A1(n433), .A2(n589), .B(n587), .C(n588), .ZN(n590) );
  OAI32D1 U15 ( .A1(n586), .A2(n742), .A3(n683), .B1(n585), .B2(n763), .ZN(
        n587) );
  OAI22D0 U16 ( .A1(n456), .A2(n778), .B1(n745), .B2(n634), .ZN(n457) );
  INVD2 U17 ( .I(n778), .ZN(n835) );
  AOI221D2 U18 ( .A1(n840), .A2(n443), .B1(n850), .B2(n445), .C(n639), .ZN(
        n640) );
  ND2D2 U19 ( .A1(n845), .A2(n443), .ZN(n636) );
  OAI22D1 U20 ( .A1(n763), .A2(n773), .B1(n445), .B2(n762), .ZN(n764) );
  AOI221D1 U21 ( .A1(n425), .A2(n851), .B1(n803), .B2(n830), .C(n461), .ZN(
        n465) );
  AOI221D2 U22 ( .A1(n463), .A2(n801), .B1(n845), .B2(n811), .C(n462), .ZN(
        n464) );
  OAI221D1 U23 ( .A1(n748), .A2(n750), .B1(n707), .B2(n783), .C(n633), .ZN(
        n644) );
  AOI221D2 U24 ( .A1(n852), .A2(n644), .B1(n849), .B2(n796), .C(n643), .ZN(
        n661) );
  OAI22D1 U25 ( .A1(n443), .A2(n718), .B1(n447), .B2(n729), .ZN(n528) );
  INVD2 U26 ( .I(n556), .ZN(n797) );
  ND2D2 U27 ( .A1(n796), .A2(n443), .ZN(n556) );
  OAI222D1 U28 ( .A1(n743), .A2(n716), .B1(n767), .B2(n584), .C1(n748), .C2(
        n758), .ZN(n588) );
  AOI21D4 U29 ( .A1(n808), .A2(n445), .B(n797), .ZN(n585) );
  OAI221D1 U30 ( .A1(n736), .A2(n729), .B1(n702), .B2(n742), .C(n594), .ZN(
        n602) );
  AOI222D1 U31 ( .A1(n801), .A2(n823), .B1(n799), .B2(n485), .C1(n795), .C2(
        n826), .ZN(n490) );
  OAI221D2 U32 ( .A1(n559), .A2(n630), .B1(n716), .B2(n782), .C(n70), .ZN(n35)
         );
  AOI221D2 U33 ( .A1(n445), .A2(n467), .B1(n820), .B2(n829), .C(n466), .ZN(
        n481) );
  CKND1 U34 ( .I(a[1]), .ZN(n447) );
  BUFFD6 U36 ( .I(a[3]), .Z(n439) );
  INVD1 U37 ( .I(n770), .ZN(n805) );
  ND2D3 U38 ( .A1(n439), .A2(n444), .ZN(n770) );
  CKND2D2 U39 ( .A1(n442), .A2(a[6]), .ZN(n702) );
  INVD4 U40 ( .I(n440), .ZN(n813) );
  CKND2D2 U41 ( .A1(n445), .A2(n437), .ZN(n716) );
  ND2D1 U42 ( .A1(n823), .A2(n835), .ZN(n720) );
  INVD1 U43 ( .I(n436), .ZN(n722) );
  INVD1 U44 ( .I(n716), .ZN(n790) );
  ND2D1 U45 ( .A1(n440), .A2(n821), .ZN(n612) );
  NR4D0 U46 ( .A1(n740), .A2(n739), .A3(n738), .A4(n737), .ZN(n789) );
  ND4D2 U47 ( .A1(n661), .A2(n426), .A3(n660), .A4(n659), .ZN(d[2]) );
  AOI221D1 U48 ( .A1(n838), .A2(n610), .B1(n609), .B2(n443), .C(n608), .ZN(
        n623) );
  ND2D1 U49 ( .A1(n813), .A2(n821), .ZN(n767) );
  ND2D1 U50 ( .A1(n444), .A2(n807), .ZN(n682) );
  INVD3 U51 ( .I(n783), .ZN(n796) );
  ND2D1 U52 ( .A1(n821), .A2(n827), .ZN(n655) );
  ND2D1 U53 ( .A1(n807), .A2(n813), .ZN(n753) );
  INVD1 U54 ( .I(n758), .ZN(n803) );
  INVD1 U55 ( .I(n745), .ZN(n801) );
  AOI221D0 U56 ( .A1(n854), .A2(n446), .B1(n836), .B2(n716), .C(n528), .ZN(
        n531) );
  INVD1 U57 ( .I(n749), .ZN(n838) );
  AOI211D1 U58 ( .A1(n856), .A2(n802), .B(n483), .C(n432), .ZN(n510) );
  IIND4D4 U59 ( .A1(n35), .A2(n64), .B1(n623), .B2(n622), .ZN(d[3]) );
  AO221D1 U60 ( .A1(n602), .A2(n809), .B1(n835), .B2(n601), .C(n600), .Z(n64)
         );
  INVD0 U61 ( .I(n742), .ZN(n791) );
  OAI222D0 U62 ( .A1(n445), .A2(n774), .B1(n742), .B2(n755), .C1(n749), .C2(
        n745), .ZN(n488) );
  CKND2 U63 ( .I(a[1]), .ZN(n446) );
  AN3XD1 U64 ( .A1(n581), .A2(n580), .A3(n583), .Z(n65) );
  ND2D1 U65 ( .A1(n443), .A2(n446), .ZN(n742) );
  AOI22D1 U66 ( .A1(n831), .A2(n799), .B1(n802), .B2(n830), .ZN(n470) );
  ND4D2 U67 ( .A1(n510), .A2(n509), .A3(n508), .A4(n507), .ZN(d[6]) );
  ND2D4 U68 ( .A1(n445), .A2(n444), .ZN(n783) );
  OAI22D1 U69 ( .A1(n638), .A2(n736), .B1(n742), .B2(n704), .ZN(n639) );
  OAI22D1 U70 ( .A1(n744), .A2(n750), .B1(n763), .B2(n783), .ZN(n684) );
  OAI222D1 U71 ( .A1(n570), .A2(n707), .B1(n569), .B2(n741), .C1(n445), .C2(
        n568), .ZN(n571) );
  AOI21D1 U72 ( .A1(n854), .A2(n810), .B(n848), .ZN(n568) );
  AOI22D1 U73 ( .A1(n802), .A2(n851), .B1(n425), .B2(n830), .ZN(n570) );
  CKND2D1 U74 ( .A1(n438), .A2(n807), .ZN(n773) );
  ND2D2 U75 ( .A1(n441), .A2(n813), .ZN(n763) );
  AOI21D0 U76 ( .A1(n683), .A2(n763), .B(n722), .ZN(n679) );
  INVD2 U77 ( .I(n442), .ZN(n832) );
  OAI33D0 U78 ( .A1(n750), .A2(n749), .A3(n748), .B1(n771), .B2(n444), .B3(
        n747), .ZN(n751) );
  OAI222D1 U79 ( .A1(n750), .A2(n759), .B1(n687), .B2(n718), .C1(n686), .C2(
        n778), .ZN(n688) );
  CKND2D0 U80 ( .A1(n780), .A2(n556), .ZN(n557) );
  AOI221D1 U81 ( .A1(n690), .A2(n742), .B1(n445), .B2(n847), .C(n558), .ZN(
        n562) );
  CKND2D2 U82 ( .A1(n835), .A2(n822), .ZN(n718) );
  AOI21D0 U83 ( .A1(n826), .A2(n835), .B(n844), .ZN(n664) );
  OA222D1 U84 ( .A1(n663), .A2(n766), .B1(n437), .B2(n560), .C1(n748), .C2(
        n559), .Z(n435) );
  ND2D1 U85 ( .A1(n445), .A2(n443), .ZN(n736) );
  CKND0 U86 ( .I(n736), .ZN(n793) );
  CKND2D0 U87 ( .A1(n438), .A2(n736), .ZN(n734) );
  INVD2 U89 ( .I(n641), .ZN(n810) );
  ND2D2 U90 ( .A1(n442), .A2(n827), .ZN(n755) );
  AOI211XD0 U91 ( .A1(n836), .A2(n437), .B(n637), .C(n846), .ZN(n642) );
  OAI22D1 U92 ( .A1(n447), .A2(n718), .B1(n445), .B2(n635), .ZN(n637) );
  NR2XD0 U93 ( .A1(n776), .A2(n775), .ZN(n777) );
  CKND2D1 U94 ( .A1(n838), .A2(n825), .ZN(n781) );
  INVD1 U95 ( .I(n781), .ZN(n840) );
  CKND2D1 U96 ( .A1(n825), .A2(n832), .ZN(n624) );
  OAI222D1 U97 ( .A1(n722), .A2(n536), .B1(n490), .B2(n749), .C1(n489), .C2(
        n753), .ZN(n494) );
  ND2D1 U98 ( .A1(n437), .A2(n799), .ZN(n726) );
  AOI221D1 U99 ( .A1(n792), .A2(n680), .B1(n429), .B2(n799), .C(n679), .ZN(
        n681) );
  NR2D0 U100 ( .A1(n791), .A2(n799), .ZN(n649) );
  AOI22D1 U101 ( .A1(n823), .A2(n810), .B1(n799), .B2(n821), .ZN(n560) );
  OAI221D1 U102 ( .A1(n665), .A2(n675), .B1(n664), .B2(n663), .C(n839), .ZN(
        n667) );
  NR2D1 U103 ( .A1(n807), .A2(n441), .ZN(n433) );
  AOI221D2 U104 ( .A1(n437), .A2(n566), .B1(n835), .B2(n565), .C(n564), .ZN(
        n582) );
  AOI221D1 U105 ( .A1(n806), .A2(n573), .B1(n572), .B2(n816), .C(n571), .ZN(
        n581) );
  OAI221D1 U106 ( .A1(n611), .A2(n586), .B1(n439), .B2(n772), .C(n699), .ZN(
        n529) );
  AOI221D1 U107 ( .A1(n835), .A2(n653), .B1(n838), .B2(n652), .C(n651), .ZN(
        n660) );
  CKND2D1 U108 ( .A1(n442), .A2(n821), .ZN(n725) );
  AOI221D1 U109 ( .A1(n829), .A2(n818), .B1(n816), .B2(n573), .C(n844), .ZN(
        n497) );
  AOI221D1 U110 ( .A1(n793), .A2(n685), .B1(n826), .B2(n436), .C(n684), .ZN(
        n686) );
  OA222D1 U111 ( .A1(n641), .A2(n634), .B1(n592), .B2(n591), .C1(n755), .C2(
        n590), .Z(n70) );
  INVD1 U112 ( .I(n559), .ZN(n795) );
  INVD6 U113 ( .I(n446), .ZN(n445) );
  AOI221D1 U114 ( .A1(n853), .A2(n443), .B1(n845), .B2(n801), .C(n631), .ZN(
        n426) );
  OAI222D1 U115 ( .A1(n465), .A2(n747), .B1(n683), .B2(n516), .C1(n443), .C2(
        n464), .ZN(n466) );
  ND2D1 U116 ( .A1(n439), .A2(n441), .ZN(n683) );
  CKND0 U117 ( .I(n683), .ZN(n824) );
  OA221D1 U118 ( .A1(n747), .A2(n742), .B1(n683), .B2(n745), .C(n435), .Z(n561) );
  ND2D1 U119 ( .A1(n437), .A2(n446), .ZN(n741) );
  OAI222D1 U120 ( .A1(n531), .A2(n773), .B1(n722), .B2(n624), .C1(n716), .C2(
        n530), .ZN(n543) );
  AOI221D1 U121 ( .A1(n828), .A2(n790), .B1(n593), .B2(n446), .C(n732), .ZN(
        n594) );
  OA221D1 U122 ( .A1(n682), .A2(n673), .B1(n672), .B2(n783), .C(n671), .Z(n430) );
  CKND2D2 U123 ( .A1(n582), .A2(n65), .ZN(d[4]) );
  CKAN2D1 U124 ( .A1(n843), .A2(n803), .Z(n72) );
  CKAN2D1 U125 ( .A1(n690), .A2(n796), .Z(n73) );
  NR3D2 U126 ( .A1(n72), .A2(n73), .A3(n678), .ZN(n714) );
  NR2D0 U127 ( .A1(n437), .A2(n677), .ZN(n74) );
  NR2D0 U128 ( .A1(n676), .A2(n749), .ZN(n185) );
  NR2D0 U129 ( .A1(n675), .A2(n674), .ZN(n192) );
  OR3D1 U130 ( .A1(n74), .A2(n185), .A3(n192), .Z(n678) );
  CKND2D3 U131 ( .A1(n714), .A2(n424), .ZN(d[1]) );
  ND2D2 U132 ( .A1(n827), .A2(n832), .ZN(n749) );
  ND2D1 U133 ( .A1(n439), .A2(n447), .ZN(n675) );
  ND2D1 U134 ( .A1(n823), .A2(n852), .ZN(n674) );
  ND3D2 U135 ( .A1(n545), .A2(n546), .A3(n547), .ZN(d[5]) );
  NR4D1 U136 ( .A1(n543), .A2(n544), .A3(n542), .A4(n541), .ZN(n545) );
  AOI221D1 U137 ( .A1(n473), .A2(n446), .B1(n815), .B2(n472), .C(n471), .ZN(
        n480) );
  OAI222D1 U138 ( .A1(n642), .A2(n641), .B1(n758), .B2(n760), .C1(n770), .C2(
        n640), .ZN(n643) );
  OAI22D1 U139 ( .A1(n470), .A2(n707), .B1(n469), .B2(n758), .ZN(n471) );
  ND2D2 U140 ( .A1(a[6]), .A2(n821), .ZN(n771) );
  INVD6 U141 ( .I(n441), .ZN(n821) );
  OAI211D0 U142 ( .A1(n555), .A2(n716), .B(n554), .C(n553), .ZN(n565) );
  AN2D1 U143 ( .A1(n717), .A2(n716), .Z(n721) );
  CKND2D1 U144 ( .A1(n445), .A2(n434), .ZN(n486) );
  CKND2D1 U145 ( .A1(n805), .A2(n445), .ZN(n584) );
  CKND2D1 U146 ( .A1(n445), .A2(n439), .ZN(n780) );
  CKND2D1 U147 ( .A1(n445), .A2(n438), .ZN(n745) );
  BUFFD4 U148 ( .I(a[7]), .Z(n442) );
  AOI221D1 U149 ( .A1(n835), .A2(n499), .B1(n795), .B2(n512), .C(n498), .ZN(
        n508) );
  AOI22D1 U150 ( .A1(n805), .A2(n825), .B1(n808), .B2(n821), .ZN(n762) );
  ND4D2 U151 ( .A1(n427), .A2(n428), .A3(n789), .A4(n788), .ZN(d[0]) );
  NR4D1 U152 ( .A1(n785), .A2(n786), .A3(n787), .A4(n784), .ZN(n788) );
  BUFFD8 U153 ( .I(n794), .Z(n444) );
  AOI221D1 U154 ( .A1(n849), .A2(n790), .B1(n852), .B2(n689), .C(n688), .ZN(
        n713) );
  OAI221D0 U155 ( .A1(n736), .A2(n682), .B1(n744), .B2(n701), .C(n681), .ZN(
        n689) );
  AOI32D0 U156 ( .A1(n441), .A2(n443), .A3(n811), .B1(n822), .B2(n632), .ZN(
        n633) );
  CKND1 U157 ( .I(n725), .ZN(n851) );
  CKND2D1 U158 ( .A1(n438), .A2(n441), .ZN(n743) );
  CKND2D1 U159 ( .A1(n441), .A2(n434), .ZN(n774) );
  CKND2D1 U160 ( .A1(n771), .A2(n725), .ZN(n573) );
  CKND2D1 U161 ( .A1(n441), .A2(n442), .ZN(n700) );
  ND2D0 U162 ( .A1(n441), .A2(n827), .ZN(n511) );
  NR2XD0 U163 ( .A1(n813), .A2(n821), .ZN(n669) );
  ND2D0 U164 ( .A1(n441), .A2(n832), .ZN(n704) );
  OA21D0 U165 ( .A1(n682), .A2(n443), .B(n615), .Z(n619) );
  OAI222D1 U166 ( .A1(n563), .A2(n755), .B1(n682), .B2(n562), .C1(n561), .C2(
        n749), .ZN(n564) );
  OAI22D0 U167 ( .A1(n763), .A2(n682), .B1(n687), .B2(n707), .ZN(n454) );
  INVD2 U168 ( .I(n612), .ZN(n823) );
  OR2D0 U169 ( .A1(n722), .A2(n747), .Z(n205) );
  OR2D0 U170 ( .A1(n687), .A2(n683), .Z(n244) );
  OR2D0 U171 ( .A1(n753), .A2(n556), .Z(n245) );
  ND3D1 U172 ( .A1(n205), .A2(n244), .A3(n245), .ZN(n534) );
  ND2D1 U173 ( .A1(n439), .A2(n813), .ZN(n747) );
  NR2XD0 U174 ( .A1(n436), .A2(n792), .ZN(n687) );
  NR4D1 U175 ( .A1(n534), .A2(n533), .A3(n532), .A4(n595), .ZN(n535) );
  AOI221D1 U176 ( .A1(n838), .A2(n459), .B1(n458), .B2(n443), .C(n457), .ZN(
        n482) );
  OAI222D1 U177 ( .A1(n779), .A2(n778), .B1(n439), .B2(n833), .C1(n777), .C2(
        n443), .ZN(n785) );
  AOI221D1 U178 ( .A1(n425), .A2(n818), .B1(n802), .B2(n824), .C(n764), .ZN(
        n779) );
  BUFFD4 U179 ( .I(a[0]), .Z(n437) );
  CKND0 U180 ( .I(n439), .ZN(n277) );
  ND3D1 U181 ( .A1(n713), .A2(n712), .A3(n711), .ZN(n310) );
  CKND1 U182 ( .I(n310), .ZN(n424) );
  AOI221D1 U183 ( .A1(n698), .A2(n851), .B1(n810), .B2(n697), .C(n696), .ZN(
        n712) );
  AN2D2 U184 ( .A1(n447), .A2(n444), .Z(n425) );
  ND2D1 U185 ( .A1(a[6]), .A2(n832), .ZN(n778) );
  ND2D1 U186 ( .A1(n447), .A2(n444), .ZN(n750) );
  ND2D0 U187 ( .A1(n805), .A2(n847), .ZN(n567) );
  ND2D0 U188 ( .A1(n793), .A2(n852), .ZN(n516) );
  NR2D0 U189 ( .A1(n625), .A2(n716), .ZN(n698) );
  ND2D0 U190 ( .A1(n441), .A2(n807), .ZN(n766) );
  CKND2D0 U191 ( .A1(n801), .A2(n443), .ZN(n703) );
  CKND0 U192 ( .I(n782), .ZN(n856) );
  INVD1 U193 ( .I(n591), .ZN(n850) );
  INVD1 U194 ( .I(n635), .ZN(n847) );
  AOI21D1 U195 ( .A1(n814), .A2(n855), .B(n842), .ZN(n569) );
  CKND2D0 U196 ( .A1(n726), .A2(n736), .ZN(n589) );
  CKND2D0 U197 ( .A1(n722), .A2(n750), .ZN(n526) );
  NR2XD0 U198 ( .A1(n853), .A2(n512), .ZN(n513) );
  NR2XD0 U200 ( .A1(n646), .A2(n765), .ZN(n606) );
  NR2D0 U201 ( .A1(n830), .A2(n841), .ZN(n638) );
  BUFFD4 U202 ( .I(n431), .Z(n443) );
  BUFFD4 U203 ( .I(a[4]), .Z(n440) );
  BUFFD4 U204 ( .I(a[5]), .Z(n441) );
  CKND0 U205 ( .I(n584), .ZN(n806) );
  AOI22D0 U206 ( .A1(n854), .A2(n796), .B1(n811), .B2(n840), .ZN(n550) );
  ND2D0 U207 ( .A1(n809), .A2(n445), .ZN(n717) );
  NR2D0 U208 ( .A1(n801), .A2(n790), .ZN(n615) );
  NR2D0 U210 ( .A1(n810), .A2(n817), .ZN(n654) );
  NR2D0 U211 ( .A1(n798), .A2(n425), .ZN(n475) );
  ND2D0 U212 ( .A1(n816), .A2(n855), .ZN(n759) );
  CKND2D0 U213 ( .A1(n815), .A2(n838), .ZN(n668) );
  NR2D0 U214 ( .A1(n715), .A2(n850), .ZN(n723) );
  ND2D0 U216 ( .A1(n828), .A2(n818), .ZN(n536) );
  CKND0 U217 ( .I(n718), .ZN(n837) );
  OA222D0 U218 ( .A1(n723), .A2(n722), .B1(n721), .B2(n720), .C1(n719), .C2(
        n718), .Z(n427) );
  OAI33D0 U219 ( .A1(n753), .A2(n444), .A3(n725), .B1(n655), .B2(n445), .B3(
        n654), .ZN(n658) );
  NR2D0 U220 ( .A1(n749), .A2(n767), .ZN(n690) );
  OAI211D0 U221 ( .A1(n821), .A2(n753), .B(n770), .C(n748), .ZN(n680) );
  NR2D0 U222 ( .A1(n825), .A2(n805), .ZN(n517) );
  OAI31D0 U223 ( .A1(n736), .A2(n817), .A3(n749), .B(n735), .ZN(n740) );
  AOI31D0 U224 ( .A1(n841), .A2(n734), .A3(n817), .B(n733), .ZN(n735) );
  AOI211D0 U225 ( .A1(n774), .A2(n655), .B(n586), .C(n741), .ZN(n476) );
  OAI22D0 U226 ( .A1(n641), .A2(n741), .B1(n742), .B2(n770), .ZN(n500) );
  NR2D0 U227 ( .A1(n805), .A2(n798), .ZN(n449) );
  CKND2D0 U228 ( .A1(n780), .A2(n682), .ZN(n525) );
  ND2D0 U229 ( .A1(n821), .A2(n832), .ZN(n611) );
  OAI21D0 U230 ( .A1(n748), .A2(n611), .B(n634), .ZN(n512) );
  CKND0 U231 ( .I(n748), .ZN(n817) );
  AOI31D0 U232 ( .A1(n729), .A2(n728), .A3(n727), .B(n726), .ZN(n730) );
  INR2D0 U233 ( .A1(n523), .B1(n663), .ZN(n708) );
  AOI22D0 U234 ( .A1(n829), .A2(n746), .B1(n831), .B2(n799), .ZN(n754) );
  CKND2D0 U235 ( .A1(n761), .A2(n758), .ZN(n746) );
  CKND0 U236 ( .I(n707), .ZN(n818) );
  NR2D0 U237 ( .A1(n511), .A2(n663), .ZN(n572) );
  CKND2D0 U238 ( .A1(n822), .A2(n841), .ZN(n634) );
  CKND1 U239 ( .I(n433), .ZN(n744) );
  CKND2D0 U240 ( .A1(n791), .A2(n277), .ZN(n719) );
  OAI21D0 U241 ( .A1(n641), .A2(n728), .B(n782), .ZN(n473) );
  CKND2D0 U242 ( .A1(n429), .A2(n841), .ZN(n630) );
  CKND0 U243 ( .I(n700), .ZN(n855) );
  CKAN2D1 U244 ( .A1(n807), .A2(n821), .Z(n429) );
  CKND2D0 U245 ( .A1(n824), .A2(n841), .ZN(n760) );
  OAI22D0 U246 ( .A1(n741), .A2(n753), .B1(n603), .B2(n742), .ZN(n610) );
  CKND2D0 U247 ( .A1(n816), .A2(n841), .ZN(n607) );
  CKND0 U248 ( .I(n774), .ZN(n831) );
  CKND2D1 U249 ( .A1(n492), .A2(n491), .ZN(n493) );
  OAI31D0 U250 ( .A1(n425), .A2(n792), .A3(n805), .B(n853), .ZN(n491) );
  OAI31D0 U251 ( .A1(n277), .A2(n797), .A3(n803), .B(n690), .ZN(n492) );
  NR2XD0 U252 ( .A1(n836), .A2(n847), .ZN(n665) );
  CKND1 U253 ( .I(n662), .ZN(n839) );
  CKND2D0 U254 ( .A1(n444), .A2(n813), .ZN(n555) );
  AOI22D0 U255 ( .A1(n796), .A2(n829), .B1(n805), .B2(n813), .ZN(n769) );
  NR2D0 U256 ( .A1(n803), .A2(n801), .ZN(n468) );
  AOI21D0 U257 ( .A1(n816), .A2(n851), .B(n692), .ZN(n504) );
  OAI33D0 U258 ( .A1(n641), .A2(n442), .A3(n767), .B1(n700), .B2(n444), .B3(
        n748), .ZN(n537) );
  OAI21D0 U259 ( .A1(n655), .A2(n747), .B(n727), .ZN(n539) );
  NR2D0 U260 ( .A1(n797), .A2(n800), .ZN(n576) );
  CKND2D0 U261 ( .A1(n716), .A2(n277), .ZN(n575) );
  CKND2D0 U262 ( .A1(n436), .A2(n825), .ZN(n645) );
  CKND2D0 U263 ( .A1(n810), .A2(n813), .ZN(n604) );
  AOI21D0 U264 ( .A1(n850), .A2(n811), .B(n692), .ZN(n695) );
  NR2XD0 U265 ( .A1(n854), .A2(n840), .ZN(n460) );
  CKND2D0 U266 ( .A1(n683), .A2(n747), .ZN(n685) );
  OAI31D0 U267 ( .A1(n702), .A2(n441), .A3(n445), .B(n636), .ZN(n558) );
  AOI21D0 U268 ( .A1(n849), .A2(n445), .B(n690), .ZN(n691) );
  ND4D0 U269 ( .A1(n792), .A2(n829), .A3(n440), .A4(n442), .ZN(n724) );
  AOI32D0 U270 ( .A1(n442), .A2(n813), .A3(n425), .B1(n799), .B2(n450), .ZN(
        n451) );
  NR2D0 U272 ( .A1(n850), .A2(n690), .ZN(n452) );
  OAI22D0 U273 ( .A1(n442), .A2(n655), .B1(n748), .B2(n725), .ZN(n450) );
  OAI22D0 U274 ( .A1(n783), .A2(n782), .B1(n781), .B2(n780), .ZN(n784) );
  OAI32D0 U275 ( .A1(n766), .A2(n475), .A3(n702), .B1(n474), .B2(n736), .ZN(
        n478) );
  AOI31D0 U276 ( .A1(n440), .A2(n827), .A3(n805), .B(n692), .ZN(n474) );
  AOI33D0 U277 ( .A1(n613), .A2(n827), .A3(n796), .B1(n847), .B2(n277), .B3(
        n793), .ZN(n614) );
  OAI31D0 U278 ( .A1(n745), .A2(n774), .A3(n747), .B(n614), .ZN(n621) );
  AOI21D0 U279 ( .A1(n682), .A2(n586), .B(n741), .ZN(n453) );
  OAI22D0 U280 ( .A1(n827), .A2(n707), .B1(n813), .B2(n655), .ZN(n647) );
  OAI22D0 U281 ( .A1(n447), .A2(n630), .B1(n629), .B2(n741), .ZN(n631) );
  AOI22D0 U282 ( .A1(n443), .A2(n811), .B1(n277), .B2(n798), .ZN(n592) );
  NR2D0 U283 ( .A1(n443), .A2(n757), .ZN(n739) );
  AOI32D0 U284 ( .A1(n425), .A2(n443), .A3(n826), .B1(n793), .B2(n552), .ZN(
        n554) );
  CKND2D0 U285 ( .A1(n748), .A2(n743), .ZN(n552) );
  AOI32D0 U287 ( .A1(n440), .A2(n832), .A3(n809), .B1(n810), .B2(n549), .ZN(
        n551) );
  OAI21D0 U288 ( .A1(n706), .A2(n736), .B(n705), .ZN(n710) );
  OAI211D0 U289 ( .A1(n441), .A2(n780), .B(n625), .C(n747), .ZN(n538) );
  CKND2D1 U290 ( .A1(n597), .A2(n596), .ZN(n601) );
  AOI21D0 U291 ( .A1(n800), .A2(n838), .B(n572), .ZN(n514) );
  AOI21D0 U292 ( .A1(n840), .A2(n810), .B(n751), .ZN(n752) );
  CKND2D0 U293 ( .A1(n823), .A2(n446), .ZN(n673) );
  NR2D0 U294 ( .A1(n440), .A2(n827), .ZN(n463) );
  ND2D1 U295 ( .A1(n443), .A2(n444), .ZN(n761) );
  BUFFD4 U296 ( .I(a[2]), .Z(n438) );
  INVD1 U298 ( .I(a[0]), .ZN(n431) );
  INVD1 U299 ( .I(n674), .ZN(n854) );
  INVD1 U300 ( .I(n599), .ZN(n820) );
  INVD1 U301 ( .I(n567), .ZN(n848) );
  INVD1 U302 ( .I(n767), .ZN(n822) );
  ND2D1 U303 ( .A1(n429), .A2(n838), .ZN(n727) );
  INVD1 U304 ( .I(n634), .ZN(n849) );
  ND2D1 U305 ( .A1(n855), .A2(n818), .ZN(n782) );
  INVD1 U306 ( .I(n728), .ZN(n845) );
  INVD1 U307 ( .I(n630), .ZN(n843) );
  ND2D1 U308 ( .A1(n790), .A2(n819), .ZN(n599) );
  INVD1 U309 ( .I(n720), .ZN(n836) );
  AO221D0 U310 ( .A1(n425), .A2(n826), .B1(n793), .B2(n809), .C(n698), .Z(n652) );
  INVD1 U311 ( .I(n598), .ZN(n844) );
  ND2D1 U312 ( .A1(n814), .A2(n829), .ZN(n699) );
  INVD1 U313 ( .I(n555), .ZN(n814) );
  INVD1 U314 ( .I(n607), .ZN(n842) );
  OAI222D0 U315 ( .A1(n781), .A2(n584), .B1(n773), .B2(n636), .C1(n497), .C2(
        n761), .ZN(n498) );
  OAI221D0 U316 ( .A1(n616), .A2(n763), .B1(n748), .B2(n758), .C(n496), .ZN(
        n499) );
  OAI222D0 U317 ( .A1(n725), .A2(n599), .B1(n722), .B2(n760), .C1(n615), .C2(
        n598), .ZN(n600) );
  AOI211D1 U318 ( .A1(n834), .A2(n802), .B(n488), .C(n487), .ZN(n489) );
  INVD1 U319 ( .I(n611), .ZN(n834) );
  OAI221D0 U320 ( .A1(n449), .A2(n612), .B1(n773), .B2(n716), .C(n448), .ZN(
        n459) );
  NR4D0 U321 ( .A1(n506), .A2(n505), .A3(n521), .A4(n522), .ZN(n507) );
  AOI221D0 U322 ( .A1(n732), .A2(n809), .B1(n808), .B2(n731), .C(n730), .ZN(
        n428) );
  AOI211D1 U323 ( .A1(n855), .A2(n520), .B(n519), .C(n518), .ZN(n547) );
  INR4D0 U324 ( .A1(n757), .B1(n524), .B2(n738), .B3(n708), .ZN(n546) );
  NR4D0 U325 ( .A1(n579), .A2(n578), .A3(n577), .A4(n737), .ZN(n580) );
  AOI221D0 U326 ( .A1(n805), .A2(n837), .B1(n845), .B2(n811), .C(n548), .ZN(
        n583) );
  INVD1 U327 ( .I(n655), .ZN(n829) );
  INVD1 U328 ( .I(n747), .ZN(n816) );
  OAI221D0 U329 ( .A1(n445), .A2(n668), .B1(n719), .B2(n674), .C(n527), .ZN(
        n544) );
  NR3D0 U330 ( .A1(n821), .A2(n445), .A3(n722), .ZN(n532) );
  INVD1 U331 ( .I(n763), .ZN(n825) );
  AOI221D0 U332 ( .A1(n797), .A2(n826), .B1(n822), .B2(n557), .C(n698), .ZN(
        n563) );
  NR4D0 U333 ( .A1(n710), .A2(n733), .A3(n709), .A4(n708), .ZN(n711) );
  INVD1 U334 ( .I(n780), .ZN(n811) );
  NR3D0 U335 ( .A1(n716), .A2(n813), .A3(n727), .ZN(n577) );
  INVD1 U336 ( .I(n726), .ZN(n800) );
  INVD1 U337 ( .I(n741), .ZN(n792) );
  INVD1 U338 ( .I(n766), .ZN(n826) );
  INVD1 U339 ( .I(n773), .ZN(n809) );
  INVD1 U340 ( .I(n703), .ZN(n802) );
  NR3D0 U341 ( .A1(n511), .A2(n748), .A3(n783), .ZN(n477) );
  NR2D1 U342 ( .A1(n624), .A2(n741), .ZN(n765) );
  INVD1 U343 ( .I(n761), .ZN(n798) );
  NR2D1 U344 ( .A1(n700), .A2(n742), .ZN(n732) );
  NR2D1 U345 ( .A1(n704), .A2(n707), .ZN(n715) );
  INVD1 U346 ( .I(n755), .ZN(n852) );
  INVD1 U347 ( .I(n701), .ZN(n819) );
  INVD1 U348 ( .I(n511), .ZN(n828) );
  NR4D0 U349 ( .A1(n455), .A2(n454), .A3(n532), .A4(n453), .ZN(n456) );
  AOI221D0 U350 ( .A1(n799), .A2(n539), .B1(n838), .B2(n538), .C(n537), .ZN(
        n540) );
  OAI222D0 U351 ( .A1(n750), .A2(n607), .B1(n606), .B2(n444), .C1(n605), .C2(
        n674), .ZN(n608) );
  ND2D1 U352 ( .A1(n437), .A2(n438), .ZN(n758) );
  OAI222D0 U353 ( .A1(n442), .A2(n769), .B1(n768), .B2(n767), .C1(n778), .C2(
        n766), .ZN(n776) );
  INVD1 U354 ( .I(n765), .ZN(n833) );
  AOI221D0 U355 ( .A1(n816), .A2(n852), .B1(n805), .B2(n825), .C(n529), .ZN(
        n530) );
  AOI221D0 U356 ( .A1(n790), .A2(n808), .B1(n795), .B2(n433), .C(n595), .ZN(
        n596) );
  INVD1 U357 ( .I(n636), .ZN(n846) );
  OA221D0 U358 ( .A1(n744), .A2(n736), .B1(n753), .B2(n663), .C(n430), .Z(n676) );
  INR4D0 U359 ( .A1(n668), .B1(n667), .B2(n666), .B3(n848), .ZN(n677) );
  OAI221D0 U360 ( .A1(n460), .A2(n773), .B1(n718), .B2(n770), .C(n567), .ZN(
        n467) );
  OAI222D0 U361 ( .A1(n504), .A2(n742), .B1(n813), .B2(n503), .C1(n502), .C2(
        n716), .ZN(n506) );
  ND2D1 U362 ( .A1(n442), .A2(n500), .ZN(n503) );
  INR2D1 U363 ( .A1(n759), .B1(n501), .ZN(n502) );
  ND2D1 U364 ( .A1(n440), .A2(n439), .ZN(n748) );
  OAI222D0 U365 ( .A1(n758), .A2(n766), .B1(n780), .B2(n645), .C1(n747), .C2(
        n703), .ZN(n653) );
  OAI222D0 U366 ( .A1(n750), .A2(n683), .B1(n484), .B2(n763), .C1(n445), .C2(
        n748), .ZN(n495) );
  OAI222D0 U367 ( .A1(n756), .A2(n755), .B1(n754), .B2(n753), .C1(n437), .C2(
        n752), .ZN(n787) );
  OAI222D0 U368 ( .A1(n761), .A2(n760), .B1(n759), .B2(n758), .C1(n445), .C2(
        n757), .ZN(n786) );
  NR3D0 U369 ( .A1(n736), .A2(n440), .A3(n611), .ZN(n646) );
  NR4D0 U370 ( .A1(n658), .A2(n657), .A3(n656), .A4(n739), .ZN(n659) );
  NR3D0 U371 ( .A1(n773), .A2(n442), .A3(n440), .ZN(n666) );
  ND2D1 U372 ( .A1(n439), .A2(n438), .ZN(n641) );
  NR4D0 U373 ( .A1(n445), .A2(n832), .A3(n761), .A4(n753), .ZN(n693) );
  OAI221D0 U374 ( .A1(n736), .A2(n725), .B1(n445), .B2(n781), .C(n724), .ZN(
        n731) );
  NR2D1 U375 ( .A1(n621), .A2(n620), .ZN(n622) );
  INVD1 U376 ( .I(n771), .ZN(n830) );
  NR3D0 U377 ( .A1(n443), .A2(n440), .A3(n683), .ZN(n595) );
  OAI222D0 U378 ( .A1(n804), .A2(n630), .B1(n556), .B2(n536), .C1(n535), .C2(
        n778), .ZN(n542) );
  INVD1 U379 ( .I(n734), .ZN(n804) );
  ND2D1 U380 ( .A1(n440), .A2(n807), .ZN(n707) );
  AOI21D1 U381 ( .A1(n790), .A2(n647), .B(n646), .ZN(n650) );
  OAI222D0 U382 ( .A1(n515), .A2(n741), .B1(n514), .B2(n748), .C1(n513), .C2(
        n761), .ZN(n519) );
  NR3D0 U383 ( .A1(n717), .A2(n440), .A3(n832), .ZN(n657) );
  ND2D1 U384 ( .A1(n440), .A2(n444), .ZN(n586) );
  ND2D1 U385 ( .A1(n438), .A2(n447), .ZN(n663) );
  OAI221D0 U386 ( .A1(n452), .A2(n641), .B1(n770), .B2(n729), .C(n451), .ZN(
        n458) );
  INVD1 U387 ( .I(n438), .ZN(n794) );
  OAI31D1 U388 ( .A1(n670), .A2(n436), .A3(n812), .B(n669), .ZN(n671) );
  OAI222D0 U389 ( .A1(n619), .A2(n772), .B1(n618), .B2(n720), .C1(n617), .C2(
        n753), .ZN(n620) );
  OA22D0 U390 ( .A1(n774), .A2(n741), .B1(n725), .B2(n616), .Z(n617) );
  OAI221D0 U391 ( .A1(n443), .A2(n729), .B1(n702), .B2(n716), .C(n691), .ZN(
        n697) );
  OAI222D0 U392 ( .A1(n576), .A2(n772), .B1(n781), .B2(n575), .C1(n574), .C2(
        n774), .ZN(n579) );
  OAI222D0 U393 ( .A1(n774), .A2(n783), .B1(n773), .B2(n772), .C1(n771), .C2(
        n770), .ZN(n775) );
  ND2D1 U394 ( .A1(n425), .A2(n437), .ZN(n559) );
  INR2D1 U395 ( .A1(a[0]), .B1(n438), .ZN(n436) );
  INVD2 U396 ( .I(a[6]), .ZN(n827) );
  INVD1 U397 ( .I(n753), .ZN(n815) );
  OAI32D1 U398 ( .A1(n559), .A2(n755), .A3(n744), .B1(n517), .B2(n516), .ZN(
        n518) );
  INVD1 U399 ( .I(n772), .ZN(n853) );
  NR4D0 U400 ( .A1(n707), .A2(n761), .A3(n755), .A4(n821), .ZN(n733) );
  OAI22D0 U401 ( .A1(n753), .A2(n750), .B1(n654), .B2(n736), .ZN(n520) );
  CKND2D0 U402 ( .A1(n669), .A2(n841), .ZN(n591) );
  ND2D1 U403 ( .A1(n669), .A2(n852), .ZN(n772) );
  NR2D0 U404 ( .A1(n635), .A2(n719), .ZN(n738) );
  OAI222D0 U405 ( .A1(n641), .A2(n720), .B1(n592), .B2(n729), .C1(n635), .C2(
        n663), .ZN(n483) );
  OAI22D0 U406 ( .A1(n720), .A2(n750), .B1(n444), .B2(n727), .ZN(n432) );
  OAI22D1 U407 ( .A1(n720), .A2(n750), .B1(n444), .B2(n727), .ZN(n662) );
  INVD0 U408 ( .I(n827), .ZN(n434) );
  NR2D0 U409 ( .A1(n436), .A2(n791), .ZN(n616) );
  ND3D0 U410 ( .A1(n810), .A2(n669), .A3(n838), .ZN(n757) );
  CKND2D1 U411 ( .A1(n835), .A2(n669), .ZN(n729) );
  INVD1 U412 ( .I(n675), .ZN(n812) );
  OAI211D1 U413 ( .A1(n700), .A2(n675), .B(n551), .C(n550), .ZN(n566) );
  OAI222D0 U414 ( .A1(n722), .A2(n598), .B1(n729), .B2(n675), .C1(n635), .C2(
        n758), .ZN(n548) );
  NR2XD0 U415 ( .A1(n803), .A2(n439), .ZN(n618) );
  OAI222D0 U416 ( .A1(n635), .A2(n444), .B1(n611), .B2(n604), .C1(n439), .C2(
        n718), .ZN(n609) );
  OAI222D0 U417 ( .A1(n755), .A2(n625), .B1(n439), .B2(n624), .C1(n749), .C2(
        n766), .ZN(n628) );
  NR2XD0 U418 ( .A1(n728), .A2(n439), .ZN(n692) );
  AOI211XD0 U419 ( .A1(n812), .A2(n437), .B(n810), .C(n803), .ZN(n605) );
  NR4D0 U420 ( .A1(n437), .A2(n827), .A3(n767), .A4(n773), .ZN(n578) );
  OAI222D0 U421 ( .A1(n703), .A2(n729), .B1(n437), .B2(n540), .C1(n783), .C2(
        n772), .ZN(n541) );
  AN4D0 U422 ( .A1(n669), .A2(n811), .A3(n437), .A4(n838), .Z(n521) );
  OAI21D0 U423 ( .A1(n437), .A2(n683), .B(n747), .ZN(n485) );
  AOI22D0 U424 ( .A1(n801), .A2(n437), .B1(n445), .B2(n810), .ZN(n484) );
  NR2D0 U425 ( .A1(n757), .A2(n437), .ZN(n709) );
  OAI33D0 U426 ( .A1(n655), .A2(n437), .A3(n444), .B1(n486), .B2(n725), .B3(
        n758), .ZN(n487) );
  NR2XD0 U427 ( .A1(n826), .A2(n433), .ZN(n672) );
  NR3D0 U428 ( .A1(n670), .A2(n425), .A3(n809), .ZN(n648) );
  NR4D0 U429 ( .A1(n683), .A2(n750), .A3(n778), .A4(n813), .ZN(n656) );
  AOI21D0 U430 ( .A1(n773), .A2(n743), .B(n778), .ZN(n626) );
  OAI222D0 U431 ( .A1(n438), .A2(n650), .B1(n649), .B2(n782), .C1(n648), .C2(
        n781), .ZN(n651) );
  ND2D1 U432 ( .A1(n438), .A2(n813), .ZN(n625) );
  ND2D1 U433 ( .A1(n440), .A2(n438), .ZN(n701) );
  OA222D0 U434 ( .A1(n745), .A2(n744), .B1(n743), .B2(n742), .C1(n747), .C2(
        n741), .Z(n756) );
  AOI22D0 U435 ( .A1(n433), .A2(n799), .B1(n796), .B2(n824), .ZN(n448) );
  AOI222D0 U436 ( .A1(n801), .A2(n818), .B1(n816), .B2(n436), .C1(n824), .C2(
        n799), .ZN(n553) );
  NR4D0 U437 ( .A1(n478), .A2(n477), .A3(n709), .A4(n476), .ZN(n479) );
  NR4D0 U438 ( .A1(n767), .A2(n755), .A3(n663), .A4(n439), .ZN(n737) );
  NR3D0 U439 ( .A1(n736), .A2(n439), .A3(n763), .ZN(n533) );
  AOI21D0 U440 ( .A1(n439), .A2(n852), .B(n812), .ZN(n768) );
  NR2D1 U441 ( .A1(n443), .A2(n439), .ZN(n670) );
  AOI31D0 U442 ( .A1(n438), .A2(n821), .A3(n792), .B(n820), .ZN(n496) );
  AOI22D0 U443 ( .A1(n819), .A2(n791), .B1(n817), .B2(n438), .ZN(n574) );
  AOI21D0 U444 ( .A1(n728), .A2(n668), .B(n438), .ZN(n627) );
  OAI222D0 U445 ( .A1(n475), .A2(n704), .B1(n468), .B2(n702), .C1(n725), .C2(
        n726), .ZN(n472) );
  OAI222D0 U446 ( .A1(n744), .A2(n556), .B1(n641), .B2(n716), .C1(n745), .C2(
        n683), .ZN(n455) );
  NR2D1 U447 ( .A1(n819), .A2(n823), .ZN(n603) );
  OAI22D0 U448 ( .A1(n439), .A2(n612), .B1(n443), .B2(n611), .ZN(n613) );
  AOI21D0 U449 ( .A1(n612), .A2(n655), .B(n682), .ZN(n501) );
  OAI21D1 U450 ( .A1(n749), .A2(n612), .B(n718), .ZN(n593) );
  AOI22D0 U451 ( .A1(n845), .A2(n526), .B1(n690), .B2(n525), .ZN(n527) );
  NR4D0 U452 ( .A1(n434), .A2(n277), .A3(n725), .A4(n758), .ZN(n505) );
  OA33D0 U453 ( .A1(n704), .A2(n748), .A3(n741), .B1(n703), .B2(n702), .B3(
        n766), .Z(n705) );
  NR3D0 U454 ( .A1(n702), .A2(n821), .A3(n707), .ZN(n523) );
  OAI22D0 U455 ( .A1(n434), .A2(n440), .B1(n441), .B2(n755), .ZN(n549) );
endmodule


module aes_sbox_7 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n62, n64, n65, n70, n81, n175, n176, n192, n277, n404, n405, n408,
         n409, n410, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857;

  AN2XD1 U28 ( .A1(n716), .A2(n715), .Z(n720) );
  OA21D1 U35 ( .A1(n700), .A2(n699), .B(n698), .Z(n705) );
  OR4D1 U199 ( .A1(n655), .A2(n574), .A3(n518), .A4(n517), .Z(n520) );
  AN2XD1 U215 ( .A1(n519), .A2(n803), .Z(n518) );
  OAI22D1 U1 ( .A1(n762), .A2(n772), .B1(n446), .B2(n761), .ZN(n763) );
  CKND2D1 U2 ( .A1(n445), .A2(n795), .ZN(n760) );
  ND3D2 U3 ( .A1(n427), .A2(n428), .A3(n429), .ZN(n678) );
  ND2D0 U4 ( .A1(n440), .A2(n443), .ZN(n742) );
  CKND2D1 U5 ( .A1(n821), .A2(n833), .ZN(n608) );
  CKND2D1 U6 ( .A1(n443), .A2(a[6]), .ZN(n773) );
  NR2XD0 U7 ( .A1(n813), .A2(n821), .ZN(n669) );
  CKND2D1 U8 ( .A1(a[6]), .A2(n821), .ZN(n770) );
  ND2D0 U9 ( .A1(n443), .A2(n444), .ZN(n699) );
  CKND2D1 U10 ( .A1(n821), .A2(n828), .ZN(n654) );
  OAI222D1 U11 ( .A1(n804), .A2(n629), .B1(n552), .B2(n532), .C1(n531), .C2(
        n777), .ZN(n538) );
  OAI22D1 U12 ( .A1(n448), .A2(n629), .B1(n628), .B2(n740), .ZN(n630) );
  INVD2 U13 ( .I(n777), .ZN(n836) );
  ND2D1 U14 ( .A1(n669), .A2(n853), .ZN(n771) );
  AOI221D1 U15 ( .A1(n855), .A2(n447), .B1(n837), .B2(n715), .C(n524), .ZN(
        n527) );
  CKND2D2 U16 ( .A1(n446), .A2(n445), .ZN(n735) );
  AOI221D2 U17 ( .A1(n794), .A2(n686), .B1(n827), .B2(n438), .C(n685), .ZN(
        n687) );
  OAI22D2 U18 ( .A1(n743), .A2(n424), .B1(n762), .B2(n426), .ZN(n685) );
  ND2D1 U19 ( .A1(a[6]), .A2(n833), .ZN(n777) );
  INVD2 U20 ( .I(n444), .ZN(n833) );
  NR4D1 U21 ( .A1(n627), .A2(n626), .A3(n843), .A4(n625), .ZN(n628) );
  OAI222D1 U22 ( .A1(n663), .A2(n765), .B1(n439), .B2(n556), .C1(n747), .C2(
        n555), .ZN(n557) );
  AOI221D1 U23 ( .A1(n439), .A2(n563), .B1(n836), .B2(n562), .C(n561), .ZN(
        n579) );
  OAI222D1 U24 ( .A1(n755), .A2(n754), .B1(n753), .B2(n752), .C1(n439), .C2(
        n751), .ZN(n785) );
  AOI21D0 U25 ( .A1(n841), .A2(n810), .B(n750), .ZN(n751) );
  OAI222D1 U26 ( .A1(n440), .A2(n649), .B1(n648), .B2(n781), .C1(n647), .C2(
        n780), .ZN(n650) );
  ND2D0 U27 ( .A1(n443), .A2(n807), .ZN(n765) );
  INVD4 U29 ( .I(n441), .ZN(n807) );
  BUFFD2 U30 ( .I(n621), .Z(n65) );
  CKND2 U31 ( .I(n662), .ZN(n840) );
  OAI22D2 U32 ( .A1(n719), .A2(n424), .B1(n795), .B2(n726), .ZN(n662) );
  ND2D0 U33 ( .A1(n448), .A2(n795), .ZN(n749) );
  ND2D1 U34 ( .A1(n795), .A2(n807), .ZN(n683) );
  INVD2 U36 ( .I(n409), .ZN(n410) );
  INVD1 U37 ( .I(a[6]), .ZN(n828) );
  INVD4 U38 ( .I(n443), .ZN(n821) );
  CKBD4 U39 ( .I(a[7]), .Z(n444) );
  INVD1 U40 ( .I(n754), .ZN(n853) );
  CKND2D1 U41 ( .A1(n807), .A2(n813), .ZN(n752) );
  ND2D2 U42 ( .A1(n444), .A2(n828), .ZN(n754) );
  CKND2D1 U43 ( .A1(n813), .A2(n821), .ZN(n766) );
  INVD2 U44 ( .I(n663), .ZN(n799) );
  OA221D0 U45 ( .A1(n749), .A2(n724), .B1(n757), .B2(n770), .C(n70), .Z(n463)
         );
  CKBD4 U46 ( .I(a[2]), .Z(n440) );
  INVD1 U47 ( .I(n654), .ZN(n830) );
  INVD1 U48 ( .I(n746), .ZN(n816) );
  OA221D1 U49 ( .A1(n555), .A2(n629), .B1(n715), .B2(n781), .C(n404), .Z(n622)
         );
  ND4D2 U50 ( .A1(n713), .A2(n711), .A3(n712), .A4(n710), .ZN(d[1]) );
  NR3D0 U51 ( .A1(n405), .A2(n408), .A3(n642), .ZN(n660) );
  OAI222D0 U52 ( .A1(n444), .A2(n768), .B1(n767), .B2(n766), .C1(n777), .C2(
        n765), .ZN(n775) );
  OAI31D1 U53 ( .A1(n438), .A2(n670), .A3(n812), .B(n669), .ZN(n671) );
  AOI21D1 U54 ( .A1(n808), .A2(n446), .B(n797), .ZN(n582) );
  ND2D1 U55 ( .A1(n823), .A2(n435), .ZN(n595) );
  INVD1 U56 ( .I(n743), .ZN(n823) );
  NR4D0 U57 ( .A1(n783), .A2(n784), .A3(n785), .A4(n782), .ZN(n786) );
  NR2D1 U58 ( .A1(n645), .A2(n764), .ZN(n603) );
  AN2XD1 U59 ( .A1(n853), .A2(n643), .Z(n405) );
  AOI221D0 U60 ( .A1(n836), .A2(n652), .B1(n839), .B2(n651), .C(n650), .ZN(
        n659) );
  AOI221D0 U61 ( .A1(n434), .A2(n827), .B1(n822), .B2(n553), .C(n697), .ZN(
        n560) );
  INVD1 U62 ( .I(n727), .ZN(n846) );
  INVD1 U63 ( .I(n752), .ZN(n815) );
  NR4D0 U64 ( .A1(n456), .A2(n455), .A3(n528), .A4(n454), .ZN(n457) );
  OA222D1 U65 ( .A1(n463), .A2(n746), .B1(n684), .B2(n512), .C1(n462), .C2(
        n445), .Z(n277) );
  AOI211D1 U66 ( .A1(n853), .A2(n491), .B(n490), .C(n489), .ZN(n505) );
  OAI222D1 U67 ( .A1(n721), .A2(n532), .B1(n486), .B2(n748), .C1(n485), .C2(
        n752), .ZN(n490) );
  ND2D2 U68 ( .A1(n446), .A2(n439), .ZN(n715) );
  CKND2D1 U69 ( .A1(n446), .A2(n440), .ZN(n744) );
  INVD4 U70 ( .I(n447), .ZN(n446) );
  INVD3 U71 ( .I(a[1]), .ZN(n447) );
  INVD1 U72 ( .I(n749), .ZN(n425) );
  AN2XD1 U73 ( .A1(n446), .A2(n795), .Z(n62) );
  ND2D2 U74 ( .A1(n444), .A2(a[6]), .ZN(n701) );
  ND2D2 U75 ( .A1(n62), .A2(n445), .ZN(n552) );
  AN3XD1 U76 ( .A1(n659), .A2(n661), .A3(n658), .Z(n64) );
  INVD2 U77 ( .I(n440), .ZN(n795) );
  AOI31D1 U78 ( .A1(n62), .A2(n853), .A3(n680), .B(n714), .ZN(n433) );
  CKND2D1 U79 ( .A1(n441), .A2(n443), .ZN(n684) );
  ND2D1 U80 ( .A1(n441), .A2(n813), .ZN(n746) );
  NR2D0 U81 ( .A1(n441), .A2(n443), .ZN(n680) );
  ND2D1 U82 ( .A1(n441), .A2(n795), .ZN(n769) );
  CKND2D0 U83 ( .A1(n779), .A2(n552), .ZN(n553) );
  ND4D2 U84 ( .A1(n579), .A2(n580), .A3(n578), .A4(n577), .ZN(d[4]) );
  AOI221D2 U85 ( .A1(n806), .A2(n570), .B1(n569), .B2(n816), .C(n568), .ZN(
        n578) );
  INVD2 U86 ( .I(n762), .ZN(n826) );
  ND2D1 U87 ( .A1(n824), .A2(n836), .ZN(n719) );
  IND4D1 U88 ( .A1(n789), .B1(n788), .B2(n787), .B3(n786), .ZN(d[0]) );
  OAI222D1 U89 ( .A1(n527), .A2(n772), .B1(n721), .B2(n623), .C1(n526), .C2(
        n715), .ZN(n539) );
  AOI21D1 U90 ( .A1(n793), .A2(n829), .B(n731), .ZN(n70) );
  AOI221D1 U91 ( .A1(n816), .A2(n853), .B1(n805), .B2(n826), .C(n525), .ZN(
        n526) );
  OAI222D2 U92 ( .A1(n567), .A2(n410), .B1(n566), .B2(n740), .C1(n446), .C2(
        n565), .ZN(n568) );
  CKND2D1 U93 ( .A1(n441), .A2(n821), .ZN(n743) );
  NR2D1 U94 ( .A1(n438), .A2(n793), .ZN(n688) );
  AOI221D1 U95 ( .A1(n839), .A2(n460), .B1(n459), .B2(n445), .C(n458), .ZN(
        n478) );
  CKND2D1 U96 ( .A1(n446), .A2(n441), .ZN(n779) );
  INVD2 U97 ( .I(n425), .ZN(n424) );
  AOI211XD0 U98 ( .A1(n835), .A2(n802), .B(n484), .C(n483), .ZN(n485) );
  AOI32D0 U99 ( .A1(n443), .A2(n445), .A3(n811), .B1(n822), .B2(n631), .ZN(
        n632) );
  INVD2 U100 ( .I(n757), .ZN(n803) );
  OAI22D0 U101 ( .A1(n457), .A2(n777), .B1(n744), .B2(n633), .ZN(n458) );
  ND4D2 U102 ( .A1(n478), .A2(n477), .A3(n476), .A4(n475), .ZN(d[7]) );
  OA221D1 U103 ( .A1(n743), .A2(n735), .B1(n752), .B2(n663), .C(n81), .Z(n676)
         );
  OA221D1 U104 ( .A1(n683), .A2(n673), .B1(n672), .B2(n426), .C(n671), .Z(n81)
         );
  OA221D1 U105 ( .A1(n633), .A2(n715), .B1(n754), .B2(n175), .C(n176), .Z(n712) );
  OA221D0 U106 ( .A1(n735), .A2(n683), .B1(n743), .B2(n700), .C(n682), .Z(n175) );
  OA222D1 U107 ( .A1(n424), .A2(n758), .B1(n688), .B2(n717), .C1(n777), .C2(
        n687), .Z(n176) );
  OA21D0 U108 ( .A1(n683), .A2(n445), .B(n612), .Z(n616) );
  INVD2 U109 ( .I(n609), .ZN(n824) );
  ND2D2 U110 ( .A1(n442), .A2(n821), .ZN(n609) );
  OA221D1 U111 ( .A1(n432), .A2(n744), .B1(n727), .B2(n779), .C(n433), .Z(n462) );
  OAI21D0 U112 ( .A1(n748), .A2(n609), .B(n717), .ZN(n590) );
  CKND2D1 U113 ( .A1(n444), .A2(n821), .ZN(n724) );
  OA221D1 U114 ( .A1(n447), .A2(n192), .B1(n596), .B2(n654), .C(n277), .Z(n477) );
  OA221D0 U115 ( .A1(n461), .A2(n772), .B1(n717), .B2(n769), .C(n564), .Z(n192) );
  OA222D1 U116 ( .A1(n640), .A2(n633), .B1(n589), .B2(n588), .C1(n587), .C2(
        n754), .Z(n404) );
  ND4D4 U117 ( .A1(n622), .A2(n65), .A3(n620), .A4(n619), .ZN(d[3]) );
  OAI222D1 U118 ( .A1(n780), .A2(n581), .B1(n772), .B2(n635), .C1(n493), .C2(
        n760), .ZN(n494) );
  AOI221D1 U119 ( .A1(n830), .A2(n818), .B1(n816), .B2(n570), .C(n845), .ZN(
        n493) );
  OR2XD1 U120 ( .A1(n676), .A2(n748), .Z(n428) );
  ND2D1 U121 ( .A1(n440), .A2(n807), .ZN(n772) );
  OAI222D1 U122 ( .A1(n641), .A2(n640), .B1(n757), .B2(n759), .C1(n639), .C2(
        n769), .ZN(n642) );
  CKND2D1 U123 ( .A1(n770), .A2(n724), .ZN(n570) );
  CKND0 U124 ( .I(n724), .ZN(n852) );
  AOI222D1 U125 ( .A1(n801), .A2(n824), .B1(n799), .B2(n481), .C1(n796), .C2(
        n827), .ZN(n486) );
  ND2D2 U126 ( .A1(n846), .A2(n445), .ZN(n635) );
  AOI211XD1 U127 ( .A1(n823), .A2(n586), .B(n584), .C(n585), .ZN(n587) );
  OAI222D1 U128 ( .A1(n754), .A2(n624), .B1(n441), .B2(n623), .C1(n748), .C2(
        n765), .ZN(n627) );
  ND2D0 U129 ( .A1(n826), .A2(n833), .ZN(n623) );
  AOI221D4 U130 ( .A1(n839), .A2(n607), .B1(n606), .B2(n445), .C(n605), .ZN(
        n620) );
  ND3D2 U131 ( .A1(n543), .A2(n542), .A3(n541), .ZN(d[5]) );
  AOI221D1 U132 ( .A1(n469), .A2(n447), .B1(n815), .B2(n468), .C(n467), .ZN(
        n476) );
  ND2D0 U133 ( .A1(n446), .A2(n795), .ZN(n426) );
  AOI221D1 U134 ( .A1(n793), .A2(n681), .B1(n680), .B2(n799), .C(n679), .ZN(
        n682) );
  AOI211XD1 U135 ( .A1(n434), .A2(n817), .B(n692), .C(n820), .ZN(n693) );
  OAI222D1 U136 ( .A1(n560), .A2(n754), .B1(n683), .B2(n559), .C1(n558), .C2(
        n748), .ZN(n561) );
  NR4D1 U137 ( .A1(n539), .A2(n540), .A3(n538), .A4(n537), .ZN(n541) );
  INVD6 U138 ( .I(n442), .ZN(n813) );
  OAI221D1 U139 ( .A1(n735), .A2(n728), .B1(n701), .B2(n741), .C(n591), .ZN(
        n599) );
  AOI221D1 U140 ( .A1(n697), .A2(n852), .B1(n810), .B2(n696), .C(n695), .ZN(
        n711) );
  CKND2D2 U141 ( .A1(n441), .A2(n440), .ZN(n640) );
  ND4D2 U142 ( .A1(n504), .A2(n505), .A3(n506), .A4(n503), .ZN(d[6]) );
  AOI211XD0 U143 ( .A1(n857), .A2(n802), .B(n479), .C(n662), .ZN(n506) );
  OAI222D0 U144 ( .A1(n727), .A2(n716), .B1(n694), .B2(n445), .C1(n693), .C2(
        n770), .ZN(n695) );
  ND2D0 U145 ( .A1(n824), .A2(n447), .ZN(n673) );
  AOI22D1 U146 ( .A1(n824), .A2(n810), .B1(n799), .B2(n821), .ZN(n556) );
  ND2D2 U147 ( .A1(n824), .A2(n842), .ZN(n727) );
  OAI222D1 U148 ( .A1(n778), .A2(n777), .B1(n441), .B2(n834), .C1(n776), .C2(
        n445), .ZN(n783) );
  ND2D1 U149 ( .A1(n836), .A2(n669), .ZN(n728) );
  CKND1 U150 ( .I(n715), .ZN(n791) );
  OA222D0 U151 ( .A1(n744), .A2(n743), .B1(n742), .B2(n741), .C1(n746), .C2(
        n740), .Z(n755) );
  AOI221D1 U152 ( .A1(n854), .A2(n445), .B1(n846), .B2(n801), .C(n630), .ZN(
        n661) );
  NR3D1 U153 ( .A1(n430), .A2(n431), .A3(n678), .ZN(n713) );
  ND2D2 U154 ( .A1(n828), .A2(n833), .ZN(n748) );
  ND2D1 U155 ( .A1(n801), .A2(n445), .ZN(n702) );
  INVD2 U156 ( .I(n744), .ZN(n801) );
  AOI31D0 U157 ( .A1(n440), .A2(n821), .A3(n793), .B(n820), .ZN(n492) );
  CKND2D1 U158 ( .A1(n442), .A2(n440), .ZN(n700) );
  CKND2D2 U159 ( .A1(n440), .A2(n448), .ZN(n663) );
  CKND2D1 U160 ( .A1(n439), .A2(n440), .ZN(n757) );
  CKND2D1 U161 ( .A1(n444), .A2(n496), .ZN(n499) );
  OAI31D0 U162 ( .A1(n701), .A2(n443), .A3(n446), .B(n635), .ZN(n554) );
  CKND1 U163 ( .I(n701), .ZN(n435) );
  INR2XD0 U164 ( .A1(n519), .B1(n663), .ZN(n707) );
  NR2XD0 U165 ( .A1(n507), .A2(n663), .ZN(n569) );
  NR2D0 U166 ( .A1(n792), .A2(n799), .ZN(n648) );
  OAI221D1 U167 ( .A1(n665), .A2(n675), .B1(n664), .B2(n663), .C(n840), .ZN(
        n667) );
  CKND2D1 U168 ( .A1(n439), .A2(n799), .ZN(n725) );
  INVD2 U169 ( .I(n769), .ZN(n805) );
  ND2D1 U170 ( .A1(n442), .A2(n807), .ZN(n706) );
  CKAN2D1 U171 ( .A1(n850), .A2(n62), .Z(n408) );
  CKND2D2 U172 ( .A1(n660), .A2(n64), .ZN(d[2]) );
  AOI221D1 U173 ( .A1(n425), .A2(n818), .B1(n802), .B2(n825), .C(n763), .ZN(
        n778) );
  AOI221D1 U174 ( .A1(n599), .A2(n809), .B1(n836), .B2(n598), .C(n597), .ZN(
        n621) );
  OAI222D1 U175 ( .A1(n742), .A2(n715), .B1(n766), .B2(n581), .C1(n747), .C2(
        n757), .ZN(n585) );
  OAI33D0 U176 ( .A1(n752), .A2(n795), .A3(n724), .B1(n654), .B2(n446), .B3(
        n653), .ZN(n657) );
  INVD1 U177 ( .I(n706), .ZN(n409) );
  AOI221D1 U178 ( .A1(n689), .A2(n741), .B1(n446), .B2(n848), .C(n554), .ZN(
        n559) );
  ND2D2 U179 ( .A1(n439), .A2(n447), .ZN(n740) );
  ND2D2 U180 ( .A1(n445), .A2(n447), .ZN(n741) );
  AOI221D1 U181 ( .A1(n829), .A2(n791), .B1(n590), .B2(n447), .C(n731), .ZN(
        n591) );
  BUFFD8 U182 ( .I(n790), .Z(n445) );
  INVD1 U183 ( .I(n735), .ZN(n794) );
  BUFFD6 U184 ( .I(a[0]), .Z(n439) );
  OAI22D0 U185 ( .A1(n741), .A2(n703), .B1(n637), .B2(n735), .ZN(n638) );
  AOI22D0 U186 ( .A1(n832), .A2(n799), .B1(n802), .B2(n831), .ZN(n466) );
  BUFFD4 U187 ( .I(a[3]), .Z(n441) );
  ND2D1 U188 ( .A1(n836), .A2(n822), .ZN(n717) );
  AOI22D0 U189 ( .A1(n802), .A2(n852), .B1(n425), .B2(n831), .ZN(n567) );
  CKND1 U190 ( .I(n438), .ZN(n721) );
  ND2D1 U191 ( .A1(n816), .A2(n435), .ZN(n604) );
  ND2D0 U192 ( .A1(n443), .A2(n833), .ZN(n703) );
  ND2D0 U193 ( .A1(n824), .A2(n853), .ZN(n674) );
  NR2D0 U194 ( .A1(n831), .A2(n435), .ZN(n637) );
  NR2D0 U195 ( .A1(n748), .A2(n766), .ZN(n689) );
  OR2D0 U196 ( .A1(n439), .A2(n677), .Z(n427) );
  OR2D0 U197 ( .A1(n675), .A2(n674), .Z(n429) );
  CKAN2D1 U198 ( .A1(n844), .A2(n803), .Z(n430) );
  CKAN2D1 U200 ( .A1(n689), .A2(n62), .Z(n431) );
  OAI33D0 U201 ( .A1(n424), .A2(n748), .A3(n747), .B1(n770), .B2(n795), .B3(
        n746), .ZN(n750) );
  OAI22D0 U202 ( .A1(n752), .A2(n424), .B1(n653), .B2(n735), .ZN(n516) );
  CKND2D0 U203 ( .A1(n856), .A2(n818), .ZN(n781) );
  ND2D0 U204 ( .A1(n805), .A2(n848), .ZN(n564) );
  NR2D0 U205 ( .A1(n810), .A2(n817), .ZN(n653) );
  AOI21D1 U206 ( .A1(n814), .A2(n856), .B(n843), .ZN(n566) );
  NR2XD0 U207 ( .A1(n827), .A2(n823), .ZN(n672) );
  CKND2D0 U208 ( .A1(n747), .A2(n742), .ZN(n548) );
  CKND0 U209 ( .I(n747), .ZN(n817) );
  CKAN2D1 U210 ( .A1(n532), .A2(n728), .Z(n465) );
  OAI32D1 U211 ( .A1(n583), .A2(n741), .A3(n684), .B1(n582), .B2(n762), .ZN(
        n584) );
  CKND0 U212 ( .I(n555), .ZN(n796) );
  ND2D0 U213 ( .A1(n443), .A2(n828), .ZN(n507) );
  BUFFD4 U214 ( .I(a[4]), .Z(n442) );
  NR2D0 U216 ( .A1(n798), .A2(n425), .ZN(n471) );
  CKND0 U217 ( .I(n581), .ZN(n806) );
  ND3D0 U218 ( .A1(n810), .A2(n669), .A3(n839), .ZN(n756) );
  ND2D0 U219 ( .A1(n839), .A2(n826), .ZN(n780) );
  AOI22D0 U220 ( .A1(n855), .A2(n62), .B1(n811), .B2(n841), .ZN(n546) );
  ND2D0 U221 ( .A1(n809), .A2(n446), .ZN(n716) );
  NR2D0 U222 ( .A1(n634), .A2(n718), .ZN(n737) );
  NR2D0 U223 ( .A1(n801), .A2(n791), .ZN(n612) );
  ND2D0 U224 ( .A1(n816), .A2(n856), .ZN(n758) );
  CKND2D0 U225 ( .A1(n815), .A2(n839), .ZN(n668) );
  CKND2D0 U226 ( .A1(n829), .A2(n818), .ZN(n532) );
  ND2D0 U227 ( .A1(n794), .A2(n853), .ZN(n512) );
  NR2D0 U228 ( .A1(n851), .A2(n689), .ZN(n453) );
  NR2D0 U229 ( .A1(n714), .A2(n851), .ZN(n722) );
  CKND2D0 U230 ( .A1(n725), .A2(n735), .ZN(n586) );
  CKND2D0 U231 ( .A1(n438), .A2(n826), .ZN(n644) );
  OAI22D0 U232 ( .A1(n445), .A2(n717), .B1(n448), .B2(n728), .ZN(n524) );
  AOI22D0 U233 ( .A1(n846), .A2(n522), .B1(n689), .B2(n521), .ZN(n523) );
  CKND2D0 U234 ( .A1(n721), .A2(n424), .ZN(n522) );
  CKND2D0 U235 ( .A1(n779), .A2(n683), .ZN(n521) );
  NR2D0 U236 ( .A1(n855), .A2(n841), .ZN(n461) );
  CKND2D1 U237 ( .A1(n488), .A2(n487), .ZN(n489) );
  AOI21D0 U238 ( .A1(n683), .A2(n583), .B(n740), .ZN(n454) );
  OAI31D0 U239 ( .A1(n735), .A2(n817), .A3(n748), .B(n734), .ZN(n739) );
  AOI31D0 U240 ( .A1(n435), .A2(n733), .A3(n817), .B(n732), .ZN(n734) );
  AOI22D0 U241 ( .A1(n445), .A2(n811), .B1(n807), .B2(n798), .ZN(n589) );
  AOI21D0 U242 ( .A1(n684), .A2(n762), .B(n721), .ZN(n679) );
  OAI21D0 U243 ( .A1(n747), .A2(n608), .B(n633), .ZN(n508) );
  OAI22D0 U244 ( .A1(n740), .A2(n752), .B1(n600), .B2(n741), .ZN(n607) );
  NR2D0 U245 ( .A1(n819), .A2(n824), .ZN(n600) );
  NR2D0 U246 ( .A1(n445), .A2(n756), .ZN(n738) );
  AOI22D0 U247 ( .A1(n830), .A2(n745), .B1(n832), .B2(n799), .ZN(n753) );
  CKND2D0 U248 ( .A1(n760), .A2(n757), .ZN(n745) );
  ND2D0 U249 ( .A1(n795), .A2(n813), .ZN(n551) );
  CKND2D0 U250 ( .A1(n792), .A2(n807), .ZN(n718) );
  CKND0 U251 ( .I(n699), .ZN(n856) );
  NR2D0 U252 ( .A1(n438), .A2(n792), .ZN(n613) );
  CKND2D0 U253 ( .A1(n825), .A2(n435), .ZN(n759) );
  NR2D0 U254 ( .A1(n803), .A2(n801), .ZN(n464) );
  AOI21D0 U255 ( .A1(n800), .A2(n839), .B(n569), .ZN(n510) );
  MAOI22D0 U256 ( .A1(n851), .A2(n807), .B1(n624), .B2(n770), .ZN(n511) );
  AOI21D0 U257 ( .A1(n441), .A2(n853), .B(n812), .ZN(n767) );
  NR2D0 U258 ( .A1(n803), .A2(n441), .ZN(n615) );
  CKND2D0 U259 ( .A1(n684), .A2(n746), .ZN(n686) );
  CKND0 U260 ( .I(n764), .ZN(n834) );
  NR2XD0 U261 ( .A1(n775), .A2(n774), .ZN(n776) );
  AOI21D0 U262 ( .A1(n816), .A2(n852), .B(n691), .ZN(n500) );
  OAI33D0 U263 ( .A1(n640), .A2(n444), .A3(n766), .B1(n699), .B2(n795), .B3(
        n747), .ZN(n533) );
  AOI22D0 U264 ( .A1(n819), .A2(n792), .B1(n817), .B2(n440), .ZN(n571) );
  CKND2D0 U265 ( .A1(n715), .A2(n807), .ZN(n572) );
  CKND0 U266 ( .I(n733), .ZN(n804) );
  CKND2D0 U267 ( .A1(n810), .A2(n813), .ZN(n601) );
  AOI21D0 U268 ( .A1(n850), .A2(n446), .B(n689), .ZN(n690) );
  ND4D0 U269 ( .A1(n793), .A2(n830), .A3(n442), .A4(n444), .ZN(n723) );
  OAI211D0 U270 ( .A1(n699), .A2(n675), .B(n547), .C(n546), .ZN(n563) );
  OAI22D0 U271 ( .A1(n426), .A2(n781), .B1(n780), .B2(n779), .ZN(n782) );
  OAI32D0 U272 ( .A1(n765), .A2(n471), .A3(n701), .B1(n470), .B2(n735), .ZN(
        n474) );
  OAI31D0 U273 ( .A1(n744), .A2(n773), .A3(n746), .B(n611), .ZN(n618) );
  AOI33D0 U274 ( .A1(n610), .A2(n828), .A3(n62), .B1(n848), .B2(n807), .B3(
        n794), .ZN(n611) );
  OAI22D0 U275 ( .A1(n441), .A2(n609), .B1(n445), .B2(n608), .ZN(n610) );
  CKND0 U276 ( .I(n608), .ZN(n835) );
  AOI21D0 U277 ( .A1(n851), .A2(n811), .B(n691), .ZN(n694) );
  AOI32D0 U278 ( .A1(n444), .A2(n813), .A3(n425), .B1(n799), .B2(n451), .ZN(
        n452) );
  CKND2D0 U279 ( .A1(n442), .A2(n795), .ZN(n583) );
  CKND2D0 U280 ( .A1(n440), .A2(n813), .ZN(n624) );
  CKND2D0 U281 ( .A1(n440), .A2(n735), .ZN(n733) );
  CKND2D1 U282 ( .A1(n594), .A2(n593), .ZN(n598) );
  OAI21D0 U283 ( .A1(n705), .A2(n735), .B(n704), .ZN(n709) );
  OA33D0 U284 ( .A1(n703), .A2(n747), .A3(n740), .B1(n702), .B2(n701), .B3(
        n765), .Z(n704) );
  OAI22D0 U285 ( .A1(n448), .A2(n717), .B1(n446), .B2(n634), .ZN(n636) );
  CKND0 U286 ( .I(n635), .ZN(n847) );
  AOI32D0 U287 ( .A1(n442), .A2(n833), .A3(n809), .B1(n810), .B2(n545), .ZN(
        n547) );
  ND2D0 U288 ( .A1(n446), .A2(a[6]), .ZN(n482) );
  BUFFD4 U289 ( .I(a[5]), .Z(n443) );
  INVD1 U290 ( .I(n674), .ZN(n855) );
  INVD1 U291 ( .I(n780), .ZN(n841) );
  INVD1 U292 ( .I(n771), .ZN(n854) );
  INVD1 U293 ( .I(n781), .ZN(n857) );
  INVD1 U294 ( .I(n564), .ZN(n849) );
  INVD1 U295 ( .I(n596), .ZN(n820) );
  INVD1 U296 ( .I(n702), .ZN(n802) );
  INVD1 U297 ( .I(n719), .ZN(n837) );
  INVD1 U298 ( .I(n633), .ZN(n850) );
  ND2D1 U299 ( .A1(n805), .A2(n446), .ZN(n581) );
  INVD1 U300 ( .I(n629), .ZN(n844) );
  INVD1 U301 ( .I(n588), .ZN(n851) );
  INVD1 U302 ( .I(n683), .ZN(n808) );
  INVD1 U303 ( .I(n634), .ZN(n848) );
  INVD1 U304 ( .I(n760), .ZN(n798) );
  ND2D1 U305 ( .A1(n791), .A2(n819), .ZN(n596) );
  INVD1 U306 ( .I(n766), .ZN(n822) );
  ND2D1 U307 ( .A1(n814), .A2(n830), .ZN(n698) );
  INVD1 U308 ( .I(n552), .ZN(n797) );
  INVD1 U309 ( .I(n604), .ZN(n843) );
  INVD1 U310 ( .I(n717), .ZN(n838) );
  INVD1 U311 ( .I(n551), .ZN(n814) );
  INVD1 U312 ( .I(n595), .ZN(n845) );
  OAI222D0 U313 ( .A1(n721), .A2(n746), .B1(n688), .B2(n684), .C1(n752), .C2(
        n552), .ZN(n530) );
  AOI222D0 U314 ( .A1(n801), .A2(n818), .B1(n816), .B2(n438), .C1(n825), .C2(
        n799), .ZN(n549) );
  NR4D0 U315 ( .A1(n474), .A2(n473), .A3(n708), .A4(n472), .ZN(n475) );
  OAI222D0 U316 ( .A1(n757), .A2(n765), .B1(n779), .B2(n644), .C1(n746), .C2(
        n702), .ZN(n652) );
  OAI222D0 U317 ( .A1(n724), .A2(n596), .B1(n721), .B2(n759), .C1(n612), .C2(
        n595), .ZN(n597) );
  OAI222D0 U318 ( .A1(n721), .A2(n595), .B1(n728), .B2(n675), .C1(n634), .C2(
        n757), .ZN(n544) );
  OAI222D0 U319 ( .A1(n722), .A2(n721), .B1(n720), .B2(n719), .C1(n718), .C2(
        n717), .ZN(n789) );
  NR4D0 U320 ( .A1(n739), .A2(n738), .A3(n737), .A4(n736), .ZN(n787) );
  AOI221D0 U321 ( .A1(n731), .A2(n809), .B1(n808), .B2(n730), .C(n729), .ZN(
        n788) );
  NR4D0 U322 ( .A1(n657), .A2(n656), .A3(n655), .A4(n738), .ZN(n658) );
  AOI221D0 U323 ( .A1(n805), .A2(n838), .B1(n846), .B2(n811), .C(n544), .ZN(
        n580) );
  NR4D0 U324 ( .A1(n576), .A2(n575), .A3(n574), .A4(n736), .ZN(n577) );
  NR2D1 U325 ( .A1(n618), .A2(n617), .ZN(n619) );
  OAI221D0 U326 ( .A1(n446), .A2(n668), .B1(n718), .B2(n674), .C(n523), .ZN(
        n540) );
  NR4D0 U327 ( .A1(n709), .A2(n732), .A3(n708), .A4(n707), .ZN(n710) );
  OAI222D0 U328 ( .A1(n424), .A2(n684), .B1(n480), .B2(n762), .C1(n446), .C2(
        n747), .ZN(n491) );
  AOI211D1 U329 ( .A1(n856), .A2(n516), .B(n515), .C(n514), .ZN(n543) );
  INR4D0 U330 ( .A1(n756), .B1(n520), .B2(n737), .B3(n707), .ZN(n542) );
  AOI221D0 U331 ( .A1(n841), .A2(n445), .B1(n851), .B2(n446), .C(n638), .ZN(
        n639) );
  NR3D0 U332 ( .A1(n715), .A2(n813), .A3(n726), .ZN(n574) );
  NR2D1 U333 ( .A1(n624), .A2(n715), .ZN(n697) );
  ND2D1 U334 ( .A1(n680), .A2(n839), .ZN(n726) );
  ND2D1 U335 ( .A1(n435), .A2(n826), .ZN(n634) );
  INVD1 U336 ( .I(n772), .ZN(n809) );
  NR2D1 U337 ( .A1(n699), .A2(n741), .ZN(n731) );
  NR3D0 U338 ( .A1(n507), .A2(n747), .A3(n426), .ZN(n473) );
  INVD1 U339 ( .I(n740), .ZN(n793) );
  NR2D1 U340 ( .A1(n623), .A2(n740), .ZN(n764) );
  NR2D1 U341 ( .A1(n703), .A2(n410), .ZN(n714) );
  AOI21D1 U342 ( .A1(n855), .A2(n810), .B(n849), .ZN(n565) );
  INVD1 U343 ( .I(n675), .ZN(n812) );
  INVD1 U344 ( .I(n725), .ZN(n800) );
  INVD1 U345 ( .I(n765), .ZN(n827) );
  INVD1 U346 ( .I(n700), .ZN(n819) );
  INVD1 U347 ( .I(n507), .ZN(n829) );
  INVD1 U348 ( .I(n748), .ZN(n839) );
  OAI222D0 U349 ( .A1(n640), .A2(n719), .B1(n589), .B2(n728), .C1(n634), .C2(
        n663), .ZN(n479) );
  INVD1 U350 ( .I(n640), .ZN(n810) );
  INR2D1 U351 ( .A1(n439), .B1(n440), .ZN(n438) );
  AOI221D0 U352 ( .A1(n799), .A2(n535), .B1(n839), .B2(n534), .C(n533), .ZN(
        n536) );
  NR4D0 U353 ( .A1(n446), .A2(n833), .A3(n760), .A4(n752), .ZN(n692) );
  OAI222D0 U354 ( .A1(n424), .A2(n604), .B1(n603), .B2(n795), .C1(n602), .C2(
        n674), .ZN(n605) );
  OAI222D0 U355 ( .A1(n634), .A2(n795), .B1(n608), .B2(n601), .C1(n441), .C2(
        n717), .ZN(n606) );
  OAI221D0 U356 ( .A1(n747), .A2(n424), .B1(n410), .B2(n426), .C(n632), .ZN(
        n643) );
  OAI222D0 U357 ( .A1(n471), .A2(n703), .B1(n464), .B2(n701), .C1(n724), .C2(
        n725), .ZN(n468) );
  OAI222D0 U358 ( .A1(n773), .A2(n426), .B1(n772), .B2(n771), .C1(n770), .C2(
        n769), .ZN(n774) );
  NR4D0 U359 ( .A1(n502), .A2(n501), .A3(n517), .A4(n518), .ZN(n503) );
  OAI222D0 U360 ( .A1(n616), .A2(n771), .B1(n615), .B2(n719), .C1(n614), .C2(
        n752), .ZN(n617) );
  OA22D0 U361 ( .A1(n773), .A2(n740), .B1(n724), .B2(n613), .Z(n614) );
  INR4D0 U362 ( .A1(n668), .B1(n667), .B2(n666), .B3(n849), .ZN(n677) );
  OAI211D1 U363 ( .A1(n551), .A2(n715), .B(n550), .C(n549), .ZN(n562) );
  OAI221D0 U364 ( .A1(n445), .A2(n728), .B1(n701), .B2(n715), .C(n690), .ZN(
        n696) );
  OAI221D0 U365 ( .A1(n735), .A2(n724), .B1(n446), .B2(n780), .C(n723), .ZN(
        n730) );
  NR3D0 U366 ( .A1(n735), .A2(n442), .A3(n608), .ZN(n645) );
  OAI222D0 U367 ( .A1(n760), .A2(n759), .B1(n758), .B2(n757), .C1(n446), .C2(
        n756), .ZN(n784) );
  OAI221D0 U368 ( .A1(n608), .A2(n583), .B1(n441), .B2(n771), .C(n698), .ZN(
        n525) );
  NR3D0 U369 ( .A1(n772), .A2(n444), .A3(n442), .ZN(n666) );
  OAI222D0 U370 ( .A1(n573), .A2(n771), .B1(n780), .B2(n572), .C1(n571), .C2(
        n773), .ZN(n576) );
  NR3D0 U371 ( .A1(n445), .A2(n442), .A3(n684), .ZN(n592) );
  ND2D1 U372 ( .A1(n441), .A2(n448), .ZN(n675) );
  NR3D0 U373 ( .A1(n436), .A2(n437), .A3(n557), .ZN(n558) );
  NR2XD0 U374 ( .A1(n837), .A2(n848), .ZN(n665) );
  AOI21D1 U375 ( .A1(n791), .A2(n646), .B(n645), .ZN(n649) );
  NR3D0 U376 ( .A1(n716), .A2(n442), .A3(n833), .ZN(n656) );
  ND2D1 U377 ( .A1(n443), .A2(n813), .ZN(n762) );
  INVD1 U378 ( .I(n770), .ZN(n831) );
  ND2D1 U379 ( .A1(n442), .A2(n441), .ZN(n747) );
  INVD1 U380 ( .I(n773), .ZN(n832) );
  INVD1 U381 ( .I(n439), .ZN(n790) );
  AOI222D0 U382 ( .A1(n62), .A2(n815), .B1(n817), .B2(n798), .C1(n800), .C2(
        n443), .ZN(n594) );
  AOI221D0 U383 ( .A1(n791), .A2(n808), .B1(n796), .B2(n823), .C(n592), .ZN(
        n593) );
  OAI222D0 U384 ( .A1(n500), .A2(n741), .B1(n813), .B2(n499), .C1(n498), .C2(
        n715), .ZN(n502) );
  INR2D1 U385 ( .A1(n758), .B1(n497), .ZN(n498) );
  OAI222D0 U386 ( .A1(n511), .A2(n740), .B1(n510), .B2(n747), .C1(n509), .C2(
        n760), .ZN(n515) );
  NR2D1 U387 ( .A1(n854), .A2(n508), .ZN(n509) );
  INVD1 U388 ( .I(n701), .ZN(n842) );
  NR2D1 U389 ( .A1(n445), .A2(n441), .ZN(n670) );
  OAI221D0 U390 ( .A1(n453), .A2(n640), .B1(n769), .B2(n728), .C(n452), .ZN(
        n459) );
  OAI221D0 U391 ( .A1(n450), .A2(n609), .B1(n772), .B2(n715), .C(n449), .ZN(
        n460) );
  NR4D0 U392 ( .A1(n530), .A2(n529), .A3(n528), .A4(n592), .ZN(n531) );
  NR3D0 U393 ( .A1(n735), .A2(n441), .A3(n762), .ZN(n529) );
  INVD1 U394 ( .I(a[1]), .ZN(n448) );
  OAI221D0 U395 ( .A1(n613), .A2(n762), .B1(n747), .B2(n757), .C(n492), .ZN(
        n495) );
  ND2D1 U396 ( .A1(n680), .A2(n435), .ZN(n629) );
  ND2D1 U397 ( .A1(n822), .A2(n435), .ZN(n633) );
  OR2D1 U398 ( .A1(n442), .A2(n828), .Z(n432) );
  INVD1 U399 ( .I(n779), .ZN(n811) );
  OAI32D0 U400 ( .A1(n555), .A2(n754), .A3(n743), .B1(n513), .B2(n512), .ZN(
        n514) );
  OAI222D0 U401 ( .A1(n446), .A2(n773), .B1(n741), .B2(n754), .C1(n748), .C2(
        n744), .ZN(n484) );
  OAI33D0 U402 ( .A1(n654), .A2(n439), .A3(n795), .B1(n482), .B2(n724), .B3(
        n757), .ZN(n483) );
  AOI211XD0 U403 ( .A1(n837), .A2(n439), .B(n636), .C(n847), .ZN(n641) );
  AOI211XD0 U404 ( .A1(n812), .A2(n439), .B(n810), .C(n803), .ZN(n602) );
  AN4D0 U405 ( .A1(n669), .A2(n811), .A3(n439), .A4(n839), .Z(n517) );
  OAI21D0 U406 ( .A1(n439), .A2(n684), .B(n746), .ZN(n481) );
  AOI22D0 U407 ( .A1(n801), .A2(n439), .B1(n446), .B2(n810), .ZN(n480) );
  NR2XD0 U408 ( .A1(n756), .A2(n439), .ZN(n708) );
  NR4D0 U409 ( .A1(n439), .A2(n828), .A3(n766), .A4(n772), .ZN(n575) );
  OAI222D0 U410 ( .A1(n702), .A2(n728), .B1(n439), .B2(n536), .C1(n426), .C2(
        n771), .ZN(n537) );
  INVD1 U411 ( .I(n552), .ZN(n434) );
  OAI211D0 U412 ( .A1(n443), .A2(n779), .B(n624), .C(n746), .ZN(n534) );
  ND2D1 U413 ( .A1(n425), .A2(n439), .ZN(n555) );
  OR3D0 U414 ( .A1(n670), .A2(n805), .A3(n448), .Z(n631) );
  AO221D0 U415 ( .A1(n425), .A2(n827), .B1(n794), .B2(n809), .C(n697), .Z(n651) );
  AOI32D0 U416 ( .A1(n425), .A2(n445), .A3(n827), .B1(n794), .B2(n548), .ZN(
        n550) );
  AOI211D1 U417 ( .A1(n773), .A2(n654), .B(n583), .C(n740), .ZN(n472) );
  AOI21D0 U418 ( .A1(n609), .A2(n654), .B(n683), .ZN(n497) );
  OAI21D0 U419 ( .A1(n654), .A2(n746), .B(n726), .ZN(n535) );
  OAI22D0 U420 ( .A1(n444), .A2(n654), .B1(n747), .B2(n724), .ZN(n451) );
  IAO21D1 U421 ( .A1(n765), .A2(n777), .B(n845), .ZN(n664) );
  AOI31D0 U422 ( .A1(n728), .A2(n727), .A3(n726), .B(n725), .ZN(n729) );
  AOI21D0 U423 ( .A1(n727), .A2(n668), .B(n440), .ZN(n626) );
  NR2D0 U424 ( .A1(n727), .A2(n441), .ZN(n691) );
  OAI21D0 U425 ( .A1(n640), .A2(n727), .B(n781), .ZN(n469) );
  OAI222D0 U426 ( .A1(n743), .A2(n552), .B1(n640), .B2(n715), .C1(n744), .C2(
        n684), .ZN(n456) );
  CKND2D1 U427 ( .A1(n669), .A2(n435), .ZN(n588) );
  AN2XD1 U428 ( .A1(n816), .A2(n792), .Z(n436) );
  AN2XD1 U429 ( .A1(n825), .A2(n801), .Z(n437) );
  CKND0 U430 ( .I(n741), .ZN(n792) );
  INVD1 U431 ( .I(n684), .ZN(n825) );
  OAI22D0 U432 ( .A1(n466), .A2(n410), .B1(n465), .B2(n757), .ZN(n467) );
  OAI22D0 U433 ( .A1(n828), .A2(n410), .B1(n813), .B2(n654), .ZN(n646) );
  INVD1 U434 ( .I(n410), .ZN(n818) );
  OAI22D0 U435 ( .A1(n762), .A2(n683), .B1(n688), .B2(n410), .ZN(n455) );
  NR3D0 U436 ( .A1(n670), .A2(n425), .A3(n809), .ZN(n647) );
  NR2D1 U437 ( .A1(n826), .A2(n805), .ZN(n513) );
  OAI31D0 U438 ( .A1(n425), .A2(n793), .A3(n805), .B(n854), .ZN(n487) );
  AOI31D0 U439 ( .A1(n442), .A2(n828), .A3(n805), .B(n691), .ZN(n470) );
  OAI22D0 U440 ( .A1(n640), .A2(n740), .B1(n741), .B2(n769), .ZN(n496) );
  NR2D1 U441 ( .A1(n805), .A2(n798), .ZN(n450) );
  AOI22D0 U442 ( .A1(n62), .A2(n830), .B1(n805), .B2(n813), .ZN(n768) );
  NR2D1 U443 ( .A1(n434), .A2(n800), .ZN(n573) );
  OAI31D0 U444 ( .A1(n807), .A2(n434), .A3(n803), .B(n689), .ZN(n488) );
  NR4D0 U445 ( .A1(a[6]), .A2(n807), .A3(n724), .A4(n757), .ZN(n501) );
  NR4D0 U446 ( .A1(n766), .A2(n754), .A3(n663), .A4(n441), .ZN(n736) );
  OAI22D0 U447 ( .A1(a[6]), .A2(n442), .B1(n443), .B2(n754), .ZN(n545) );
  NR3D0 U448 ( .A1(n701), .A2(n821), .A3(n410), .ZN(n519) );
  NR4D0 U449 ( .A1(n410), .A2(n760), .A3(n754), .A4(n821), .ZN(n732) );
  OAI211D0 U450 ( .A1(n821), .A2(n752), .B(n769), .C(n747), .ZN(n681) );
  AOI22D0 U451 ( .A1(n823), .A2(n799), .B1(n62), .B2(n825), .ZN(n449) );
  NR3D0 U452 ( .A1(n821), .A2(n446), .A3(n721), .ZN(n528) );
  AOI22D1 U453 ( .A1(n805), .A2(n826), .B1(n808), .B2(n821), .ZN(n761) );
  AOI221D1 U454 ( .A1(n836), .A2(n495), .B1(n796), .B2(n508), .C(n494), .ZN(
        n504) );
  NR4D0 U455 ( .A1(n684), .A2(n424), .A3(n777), .A4(n813), .ZN(n655) );
  AOI21D0 U456 ( .A1(n772), .A2(n742), .B(n777), .ZN(n625) );
endmodule


module aes_sbox_6 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n4, n5, n6, n8, n10, n11, n12, n16, n17, n18, n19, n21, n22,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n40, n41, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53, n55, n56,
         n57, n59, n60, n61, n64, n65, n66, n68, n71, n72, n82, n83, n84, n86,
         n90, n91, n92, n93, n94, n97, n98, n101, n103, n104, n105, n106, n109,
         n111, n114, n115, n116, n119, n120, n122, n123, n135, n136, n137,
         n139, n142, n144, n157, n161, n162, n164, n172, n174, n181, n182,
         n190, n197, n202, n203, n204, n212, n226, n231, n232, n233, n253,
         n254, n257, n258, n269, n270, n278, n286, n297, n312, n315, n323,
         n335, n348, n349, n350, n359, n360, net7259, net7257, net7255,
         net7573, net7579, net7581, net7583, net7585, net7587, net7589,
         net8759, net8948, net9018, net11484, net12162, net12727, net12782,
         n373, n271, n13, n42, n63, n67, n69, n70, n117, n148, n304, n305,
         n306, n389, n390, n398, n399, n400, n404, n405, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716;

  AN2XD1 U28 ( .A1(n662), .A2(net12727), .Z(n665) );
  OA21D1 U35 ( .A1(n650), .A2(n164), .B(n649), .Z(n653) );
  OR3D1 U88 ( .A1(n623), .A2(n53), .A3(net8759), .Z(n593) );
  OR4D1 U199 ( .A1(n612), .A2(n544), .A3(n349), .A4(n350), .Z(n498) );
  AO21D1 U297 ( .A1(n68), .A2(n29), .B(n671), .Z(n475) );
  AN2XD1 U215 ( .A1(n348), .A2(n55), .Z(n349) );
  OAI222D1 U1 ( .A1(n538), .A2(n157), .B1(n537), .B2(n123), .C1(net7255), .C2(
        n536), .ZN(n539) );
  OAI32D2 U2 ( .A1(n552), .A2(n122), .A3(n181), .B1(n551), .B2(n101), .ZN(n553) );
  NR4D1 U3 ( .A1(n589), .A2(n588), .A3(n712), .A4(n587), .ZN(n590) );
  OAI221D1 U4 ( .A1(n675), .A2(n135), .B1(n162), .B2(n122), .C(n560), .ZN(n565) );
  INVD2 U5 ( .I(n63), .ZN(n5) );
  AOI221D2 U6 ( .A1(n117), .A2(n304), .B1(n33), .B2(n57), .C(n531), .ZN(n532)
         );
  NR4D1 U7 ( .A1(n469), .A2(n468), .A3(n506), .A4(n467), .ZN(n470) );
  AOI22D1 U8 ( .A1(n53), .A2(n32), .B1(n50), .B2(n37), .ZN(n687) );
  AOI221D1 U9 ( .A1(n64), .A2(n40), .B1(n56), .B2(n33), .C(n688), .ZN(n695) );
  OAI22D0 U10 ( .A1(n101), .A2(n91), .B1(net7255), .B2(n687), .ZN(n688) );
  IAO22D0 U11 ( .B1(n715), .B2(n51), .A1(n586), .A2(n93), .ZN(n492) );
  ND2D1 U12 ( .A1(a[6]), .A2(n37), .ZN(n93) );
  CKND2D1 U13 ( .A1(n53), .A2(net7255), .ZN(n286) );
  INVD1 U14 ( .I(n114), .ZN(n64) );
  ND4D3 U15 ( .A1(n550), .A2(n549), .A3(n548), .A4(n547), .ZN(d[4]) );
  AOI221XD4 U16 ( .A1(net8948), .A2(n713), .B1(n71), .B2(n1), .C(n558), .ZN(
        n584) );
  OAI222D2 U17 ( .A1(n226), .A2(n233), .B1(n278), .B2(n557), .C1(n63), .C2(
        n556), .ZN(n558) );
  INVD3 U18 ( .I(n162), .ZN(n16) );
  NR2XD1 U19 ( .A1(n27), .A2(n16), .ZN(n596) );
  ND2D2 U20 ( .A1(n16), .A2(n32), .ZN(n232) );
  NR2D0 U21 ( .A1(n136), .A2(net7585), .ZN(n172) );
  OAI222D1 U22 ( .A1(n680), .A2(net12727), .B1(n97), .B2(n286), .C1(n116), 
        .C2(n106), .ZN(n554) );
  OA221D4 U23 ( .A1(n72), .A2(n305), .B1(n86), .B2(n306), .C(n389), .Z(n549)
         );
  OAI221D1 U24 ( .A1(n116), .A2(n148), .B1(n157), .B2(n696), .C(n594), .ZN(
        n601) );
  ND2D2 U25 ( .A1(n12), .A2(n72), .ZN(n231) );
  INVD1 U26 ( .I(n109), .ZN(n42) );
  CKND4 U27 ( .I(n42), .ZN(n63) );
  ND2D0 U29 ( .A1(net7579), .A2(n30), .ZN(n109) );
  AOI221D2 U30 ( .A1(n52), .A2(n297), .B1(n540), .B2(n117), .C(n539), .ZN(n548) );
  INVD2 U31 ( .I(n257), .ZN(n34) );
  ND2D2 U32 ( .A1(net7585), .A2(net7587), .ZN(n226) );
  INVD2 U33 ( .I(net7259), .ZN(net7255) );
  INVD6 U34 ( .I(net7583), .ZN(n45) );
  BUFFD6 U36 ( .I(a[3]), .Z(net7585) );
  ND2D1 U37 ( .A1(net7589), .A2(net7259), .ZN(n123) );
  INVD2 U38 ( .I(n70), .ZN(net12727) );
  ND2D1 U39 ( .A1(net7587), .A2(net7259), .ZN(n203) );
  INVD3 U40 ( .I(net7579), .ZN(n25) );
  BUFFD6 U41 ( .I(a[4]), .Z(net7583) );
  ND2D2 U42 ( .A1(net7583), .A2(n37), .ZN(n257) );
  AOI221D0 U43 ( .A1(n716), .A2(net7259), .B1(n21), .B2(net12727), .C(n502), 
        .ZN(n505) );
  INVD4 U44 ( .I(net7585), .ZN(n51) );
  AOI221D1 U45 ( .A1(n648), .A2(n6), .B1(n48), .B2(n647), .C(n646), .ZN(n658)
         );
  AOI221D0 U46 ( .A1(n53), .A2(n711), .B1(n12), .B2(n47), .C(n323), .ZN(n550)
         );
  INVD1 U47 ( .I(n120), .ZN(n35) );
  AOI211D1 U48 ( .A1(n21), .A2(net12162), .B(n595), .C(n11), .ZN(n599) );
  ND2D2 U49 ( .A1(net7257), .A2(net7573), .ZN(n696) );
  ND2D1 U50 ( .A1(net7585), .A2(n37), .ZN(n120) );
  ND2D1 U51 ( .A1(net7581), .A2(n45), .ZN(n101) );
  ND2D1 U52 ( .A1(net7585), .A2(net7581), .ZN(n181) );
  ND2D1 U53 ( .A1(net7585), .A2(net7573), .ZN(n94) );
  INVD1 U54 ( .I(n203), .ZN(n59) );
  INVD2 U55 ( .I(n696), .ZN(n705) );
  ND2D1 U56 ( .A1(net7581), .A2(n25), .ZN(n651) );
  ND2D2 U57 ( .A1(n34), .A2(n16), .ZN(n136) );
  OA22D0 U58 ( .A1(n90), .A2(n123), .B1(n139), .B2(n253), .Z(n576) );
  NR2D1 U59 ( .A1(n164), .A2(n122), .ZN(n671) );
  NR2D2 U60 ( .A1(n114), .A2(n72), .ZN(net8948) );
  INVD1 U61 ( .I(n86), .ZN(n22) );
  ND3D1 U62 ( .A1(n454), .A2(n455), .A3(n456), .ZN(n516) );
  OAI222D0 U63 ( .A1(n543), .A2(n92), .B1(n83), .B2(n542), .C1(n541), .C2(n90), 
        .ZN(n546) );
  INVD2 U64 ( .I(n94), .ZN(n53) );
  IIND4D4 U65 ( .A1(n67), .A2(n69), .B1(n489), .B2(n488), .ZN(d[7]) );
  AO221D1 U66 ( .A1(n19), .A2(n473), .B1(n472), .B2(n72), .C(n471), .Z(n67) );
  OAI221D1 U67 ( .A1(net7259), .A2(n449), .B1(n270), .B2(n212), .C(n450), .ZN(
        n69) );
  OAI222D1 U68 ( .A1(n226), .A2(n144), .B1(n278), .B2(n135), .C1(n232), .C2(
        net9018), .ZN(n448) );
  CKND3 U69 ( .I(a[1]), .ZN(net7259) );
  CKND2D2 U70 ( .A1(n72), .A2(net7259), .ZN(n122) );
  AN2D1 U71 ( .A1(net7585), .A2(n45), .Z(n117) );
  INVD1 U72 ( .I(n675), .ZN(n461) );
  ND2D1 U73 ( .A1(net7255), .A2(n72), .ZN(n675) );
  OA221D0 U74 ( .A1(n390), .A2(a[1]), .B1(n111), .B2(n398), .C(n399), .Z(n489)
         );
  AN2XD1 U75 ( .A1(net7257), .A2(net7589), .Z(n70) );
  INVD3 U76 ( .I(net7589), .ZN(n72) );
  INVD1 U77 ( .I(n111), .ZN(n43) );
  ND2D1 U78 ( .A1(n51), .A2(n45), .ZN(n111) );
  AOI31D1 U79 ( .A1(net11484), .A2(n37), .A3(n68), .B(n38), .ZN(n435) );
  OAI221D0 U80 ( .A1(n253), .A2(n101), .B1(n116), .B2(n106), .C(n435), .ZN(
        n434) );
  ND4D2 U81 ( .A1(n618), .A2(n617), .A3(n616), .A4(n615), .ZN(d[2]) );
  CKND2D1 U82 ( .A1(net7583), .A2(net7573), .ZN(n552) );
  CKND2D1 U83 ( .A1(n72), .A2(net7573), .ZN(n103) );
  AOI221D1 U84 ( .A1(n59), .A2(n512), .B1(n19), .B2(n511), .C(n510), .ZN(n513)
         );
  OAI222D0 U85 ( .A1(n161), .A2(n135), .B1(net12162), .B2(n513), .C1(n696), 
        .C2(n92), .ZN(n514) );
  AOI221D1 U86 ( .A1(n64), .A2(n6), .B1(n55), .B2(n27), .C(n475), .ZN(n479) );
  ND2D3 U87 ( .A1(net7259), .A2(net7573), .ZN(n114) );
  OAI221D1 U89 ( .A1(n258), .A2(n552), .B1(net7585), .B2(n92), .C(n649), .ZN(
        n503) );
  ND4D2 U90 ( .A1(n660), .A2(n658), .A3(n659), .A4(n657), .ZN(d[1]) );
  AOI221D2 U91 ( .A1(n477), .A2(n57), .B1(n12), .B2(n47), .C(n476), .ZN(n478)
         );
  AOI221D1 U92 ( .A1(n22), .A2(n610), .B1(n19), .B2(n609), .C(n608), .ZN(n616)
         );
  OAI222D0 U93 ( .A1(net11484), .A2(n607), .B1(n606), .B2(n82), .C1(n605), 
        .C2(n83), .ZN(n608) );
  INVD2 U94 ( .I(n136), .ZN(n12) );
  OAI221D1 U95 ( .A1(n619), .A2(n190), .B1(n202), .B2(net9018), .C(n18), .ZN(
        n621) );
  OA222D1 U96 ( .A1(n479), .A2(net12782), .B1(n181), .B2(n493), .C1(n72), .C2(
        n478), .Z(n450) );
  CKND2D0 U97 ( .A1(net7589), .A2(n59), .ZN(n668) );
  NR2D0 U98 ( .A1(n304), .A2(n59), .ZN(n606) );
  INVD1 U99 ( .I(n64), .ZN(n148) );
  AOI221D1 U100 ( .A1(n29), .A2(n71), .B1(n559), .B2(net7259), .C(n671), .ZN(
        n560) );
  AOI221D1 U101 ( .A1(n49), .A2(n565), .B1(n22), .B2(n564), .C(n269), .ZN(n583) );
  AOI221D1 U102 ( .A1(n68), .A2(n634), .B1(n633), .B2(n59), .C(n632), .ZN(n635) );
  OAI22D0 U103 ( .A1(n144), .A2(n114), .B1(net7573), .B2(n137), .ZN(n204) );
  ND4D2 U104 ( .A1(n584), .A2(n583), .A3(n582), .A4(n581), .ZN(d[3]) );
  OR2XD1 U105 ( .A1(n533), .A2(n182), .Z(n452) );
  AOI221D1 U106 ( .A1(n61), .A2(n31), .B1(n36), .B2(n528), .C(n648), .ZN(n534)
         );
  OAI222D2 U107 ( .A1(net9018), .A2(n98), .B1(net7589), .B2(n530), .C1(n116), 
        .C2(n312), .ZN(n531) );
  CKND2D1 U108 ( .A1(net7579), .A2(n37), .ZN(n139) );
  OAI222D1 U109 ( .A1(n142), .A2(n335), .B1(n441), .B2(n115), .C1(n442), .C2(
        n111), .ZN(n437) );
  AOI211D1 U110 ( .A1(n404), .A2(n56), .B(n443), .C(n444), .ZN(n442) );
  AOI221D1 U111 ( .A1(n461), .A2(n637), .B1(n31), .B2(n65), .C(n636), .ZN(n638) );
  OAI222D1 U112 ( .A1(n136), .A2(n662), .B1(n645), .B2(n72), .C1(n644), .C2(
        n93), .ZN(n646) );
  CKND0 U113 ( .I(n122), .ZN(n304) );
  OAI222D0 U114 ( .A1(net7255), .A2(n90), .B1(n122), .B2(n63), .C1(n115), .C2(
        n119), .ZN(n443) );
  AOI22D2 U115 ( .A1(n34), .A2(n48), .B1(n59), .B2(n37), .ZN(n530) );
  ND3D2 U116 ( .A1(n520), .A2(n519), .A3(n518), .ZN(d[5]) );
  OR2XD1 U117 ( .A1(n532), .A2(n115), .Z(n453) );
  ND2D2 U118 ( .A1(net7257), .A2(net7587), .ZN(n119) );
  CKND2 U119 ( .I(net8948), .ZN(n312) );
  AOI222D1 U120 ( .A1(n57), .A2(n34), .B1(n59), .B2(n446), .C1(net8948), .C2(
        n31), .ZN(n441) );
  AO31D1 U121 ( .A1(n705), .A2(n5), .A3(n633), .B(n661), .Z(n476) );
  CKND2D2 U122 ( .A1(a[6]), .A2(n25), .ZN(n86) );
  CKND2D0 U123 ( .A1(n37), .A2(n25), .ZN(n258) );
  ND2D4 U124 ( .A1(n30), .A2(n25), .ZN(n115) );
  ND2D1 U125 ( .A1(n22), .A2(n197), .ZN(n135) );
  NR2D1 U126 ( .A1(n45), .A2(n37), .ZN(n197) );
  ND2D1 U127 ( .A1(n19), .A2(n32), .ZN(n83) );
  AOI221D1 U128 ( .A1(n19), .A2(n573), .B1(n572), .B2(n72), .C(n571), .ZN(n582) );
  NR3D1 U129 ( .A1(n631), .A2(n458), .A3(n457), .ZN(n660) );
  CKND2D1 U130 ( .A1(n93), .A2(n139), .ZN(n297) );
  CKND0 U131 ( .I(n139), .ZN(n6) );
  OAI222D0 U132 ( .A1(n83), .A2(n286), .B1(n91), .B2(n231), .C1(n400), .C2(
        n103), .ZN(n373) );
  AOI221D1 U133 ( .A1(n28), .A2(n40), .B1(n117), .B2(n297), .C(n13), .ZN(n400)
         );
  OAI222D1 U134 ( .A1(n685), .A2(n63), .B1(n684), .B2(n111), .C1(net12162), 
        .C2(n683), .ZN(n700) );
  CKND2D1 U135 ( .A1(n45), .A2(n37), .ZN(n97) );
  OA211D0 U136 ( .A1(n164), .A2(n190), .B(n523), .C(n522), .Z(n305) );
  OA211D0 U137 ( .A1(n527), .A2(net12727), .B(n526), .C(n525), .Z(n306) );
  AN3XD1 U138 ( .A1(n451), .A2(n452), .A3(n453), .Z(n389) );
  AOI211XD0 U139 ( .A1(n61), .A2(n41), .B(n38), .C(n643), .ZN(n644) );
  INVD1 U140 ( .I(n212), .ZN(n28) );
  ND2D1 U141 ( .A1(n37), .A2(n30), .ZN(n212) );
  OAI21D0 U142 ( .A1(n212), .A2(net12782), .B(n137), .ZN(n512) );
  AOI221D1 U143 ( .A1(n117), .A2(n5), .B1(n53), .B2(n32), .C(n503), .ZN(n504)
         );
  OAI22D1 U144 ( .A1(net8759), .A2(n591), .B1(n590), .B2(n123), .ZN(n592) );
  OA21D0 U145 ( .A1(n226), .A2(n136), .B(n82), .Z(n390) );
  OA222D0 U146 ( .A1(n484), .A2(n651), .B1(n480), .B2(n162), .C1(n139), .C2(
        n668), .Z(n398) );
  OA22D0 U147 ( .A1(n482), .A2(n157), .B1(n481), .B2(n106), .Z(n399) );
  AN2D1 U148 ( .A1(n335), .A2(n135), .Z(n481) );
  OAI22D1 U149 ( .A1(n72), .A2(n663), .B1(net8759), .B2(n135), .ZN(n502) );
  OAI22D0 U150 ( .A1(n111), .A2(n148), .B1(n611), .B2(n675), .ZN(n497) );
  AOI221D1 U151 ( .A1(n4), .A2(n72), .B1(n12), .B2(n57), .C(n592), .ZN(n618)
         );
  CKND1 U152 ( .I(n72), .ZN(net12162) );
  AN4D1 U153 ( .A1(n197), .A2(n47), .A3(net12162), .A4(n19), .Z(n350) );
  NR2D0 U154 ( .A1(n686), .A2(net12162), .ZN(n655) );
  OA222D0 U155 ( .A1(n119), .A2(n120), .B1(n680), .B2(n122), .C1(net12782), 
        .C2(n123), .Z(n685) );
  INVD8 U156 ( .I(net7581), .ZN(n37) );
  CKND0 U157 ( .I(n157), .ZN(n40) );
  INVD1 U158 ( .I(n271), .ZN(n13) );
  ND2D1 U159 ( .A1(n35), .A2(n16), .ZN(n271) );
  AOI21D1 U160 ( .A1(n31), .A2(n22), .B(n13), .ZN(n202) );
  OAI222D0 U161 ( .A1(n139), .A2(n270), .B1(n142), .B2(n104), .C1(n254), .C2(
        n271), .ZN(n269) );
  OAI222D0 U162 ( .A1(n142), .A2(n271), .B1(n135), .B2(n190), .C1(n232), .C2(
        n106), .ZN(n323) );
  ND4D2 U163 ( .A1(n405), .A2(n424), .A3(n425), .A4(n426), .ZN(d[6]) );
  AOI211D0 U164 ( .A1(n1), .A2(n56), .B(n448), .C(n204), .ZN(n405) );
  CKND0 U165 ( .I(n82), .ZN(n1) );
  INVD1 U166 ( .I(n161), .ZN(n56) );
  OR2XD1 U167 ( .A1(n257), .A2(n86), .Z(n144) );
  AOI22D1 U168 ( .A1(n72), .A2(n47), .B1(n51), .B2(n60), .ZN(n278) );
  BUFFD1 U169 ( .I(n203), .Z(net9018) );
  AOI211XD0 U170 ( .A1(n5), .A2(n436), .B(n437), .C(n438), .ZN(n424) );
  OAI222D0 U171 ( .A1(n148), .A2(n181), .B1(n447), .B2(n101), .C1(net7255), 
        .C2(n116), .ZN(n436) );
  AOI22D0 U172 ( .A1(n57), .A2(net12162), .B1(net7255), .B2(n48), .ZN(n447) );
  INVD1 U173 ( .I(n119), .ZN(n57) );
  INVD2 U174 ( .I(n226), .ZN(n48) );
  ND2D1 U175 ( .A1(net7583), .A2(net7585), .ZN(n116) );
  ND2D3 U176 ( .A1(net7589), .A2(net7573), .ZN(n142) );
  ND2D0 U177 ( .A1(n29), .A2(n40), .ZN(n335) );
  OAI21D0 U178 ( .A1(net12162), .A2(n181), .B(net12782), .ZN(n446) );
  INVD1 U179 ( .I(n98), .ZN(n31) );
  CKND0 U180 ( .I(n258), .ZN(n404) );
  ND2D0 U181 ( .A1(net7581), .A2(a[6]), .ZN(n90) );
  OAI33D0 U182 ( .A1(n212), .A2(net12162), .A3(net7573), .B1(n445), .B2(n139), 
        .B3(n106), .ZN(n444) );
  BUFFD8 U183 ( .I(n66), .Z(net7573) );
  CKND2D0 U184 ( .A1(net7255), .A2(a[6]), .ZN(n445) );
  ND2D1 U185 ( .A1(net7589), .A2(net7587), .ZN(n106) );
  ND2D1 U186 ( .A1(n439), .A2(n440), .ZN(n438) );
  OAI31D0 U187 ( .A1(n51), .A2(n61), .A3(n55), .B(n174), .ZN(n439) );
  INVD1 U188 ( .I(n315), .ZN(n61) );
  INVD1 U189 ( .I(n106), .ZN(n55) );
  NR2D0 U190 ( .A1(n115), .A2(n97), .ZN(n174) );
  OAI31D0 U191 ( .A1(n64), .A2(n68), .A3(n53), .B(n4), .ZN(n440) );
  INVD1 U192 ( .I(n123), .ZN(n68) );
  CKND0 U193 ( .I(n92), .ZN(n4) );
  AOI221D1 U194 ( .A1(n22), .A2(n434), .B1(net8948), .B2(n359), .C(n373), .ZN(
        n425) );
  NR2D1 U195 ( .A1(n65), .A2(n304), .ZN(n253) );
  CKND0 U196 ( .I(net7573), .ZN(net11484) );
  INVD1 U197 ( .I(n270), .ZN(n38) );
  OAI21D0 U198 ( .A1(n116), .A2(n258), .B(n233), .ZN(n359) );
  ND2D1 U200 ( .A1(net7587), .A2(n51), .ZN(n91) );
  NR4D0 U201 ( .A1(n427), .A2(n428), .A3(n350), .A4(n349), .ZN(n426) );
  OAI222D0 U202 ( .A1(n429), .A2(n122), .B1(n45), .B2(n430), .C1(n431), .C2(
        net12727), .ZN(n427) );
  AOI21D0 U203 ( .A1(n117), .A2(n6), .B(n172), .ZN(n429) );
  ND2D1 U204 ( .A1(net7579), .A2(n433), .ZN(n430) );
  BUFFD4 U205 ( .I(a[7]), .Z(net7579) );
  OAI22D0 U206 ( .A1(n226), .A2(n123), .B1(n122), .B2(n94), .ZN(n433) );
  INR2D1 U207 ( .A1(n105), .B1(n432), .ZN(n431) );
  ND2D0 U208 ( .A1(n117), .A2(n2), .ZN(n105) );
  AOI21D0 U209 ( .A1(n257), .A2(n212), .B(n182), .ZN(n432) );
  ND2D2 U210 ( .A1(net7573), .A2(n51), .ZN(n182) );
  NR4D0 U211 ( .A1(a[6]), .A2(n51), .A3(n139), .A4(n106), .ZN(n428) );
  CKND2D0 U212 ( .A1(net7255), .A2(net7585), .ZN(n84) );
  OAI222D1 U213 ( .A1(n599), .A2(n226), .B1(n106), .B2(n104), .C1(n94), .C2(
        n598), .ZN(n600) );
  OAI222D1 U214 ( .A1(n707), .A2(n591), .B1(n315), .B2(n335), .C1(n509), .C2(
        n86), .ZN(n515) );
  OA221D0 U216 ( .A1(n474), .A2(n91), .B1(n663), .B2(n94), .C(n535), .Z(n449)
         );
  BUFFD16 U217 ( .I(a[5]), .Z(net7581) );
  AOI221D1 U218 ( .A1(n8), .A2(n71), .B1(n5), .B2(n641), .C(n640), .ZN(n659)
         );
  IND4D2 U219 ( .A1(n704), .B1(n703), .B2(n702), .B3(n701), .ZN(d[0]) );
  NR4D1 U220 ( .A1(n698), .A2(n699), .A3(n700), .A4(n697), .ZN(n701) );
  OAI222D1 U221 ( .A1(n695), .A2(n86), .B1(net7585), .B2(n710), .C1(n694), 
        .C2(n72), .ZN(n698) );
  INVD3 U222 ( .I(a[6]), .ZN(n30) );
  ND2D2 U223 ( .A1(net7579), .A2(a[6]), .ZN(n162) );
  AOI211XD1 U224 ( .A1(n35), .A2(n555), .B(n553), .C(n554), .ZN(n556) );
  OR2D0 U225 ( .A1(n534), .A2(n63), .Z(n451) );
  OR2D0 U226 ( .A1(n505), .A2(n91), .Z(n454) );
  OR2D0 U227 ( .A1(n142), .A2(n585), .Z(n455) );
  OR2D0 U228 ( .A1(n504), .A2(net12727), .Z(n456) );
  CKND2D0 U229 ( .A1(n32), .A2(n25), .ZN(n585) );
  NR4D1 U230 ( .A1(n517), .A2(n516), .A3(n515), .A4(n514), .ZN(n518) );
  AOI221D1 U231 ( .A1(n5), .A2(n601), .B1(n8), .B2(n705), .C(n600), .ZN(n617)
         );
  AOI221D1 U232 ( .A1(n174), .A2(n122), .B1(net7255), .B2(n10), .C(n529), .ZN(
        n533) );
  AOI221D1 U233 ( .A1(n17), .A2(n72), .B1(n715), .B2(net7255), .C(n597), .ZN(
        n598) );
  CKND2 U234 ( .I(n117), .ZN(net12782) );
  INVD2 U235 ( .I(n182), .ZN(n50) );
  IAO21D2 U236 ( .A1(n182), .A2(net8759), .B(n61), .ZN(n551) );
  OAI211D0 U237 ( .A1(net7581), .A2(n84), .B(n586), .C(net12782), .ZN(n511) );
  OAI31D0 U238 ( .A1(n162), .A2(net7581), .A3(net7255), .B(n231), .ZN(n529) );
  CKND2D0 U239 ( .A1(net7587), .A2(net7581), .ZN(n680) );
  ND2D0 U240 ( .A1(net7581), .A2(n30), .ZN(n360) );
  ND2D0 U241 ( .A1(net7581), .A2(net7579), .ZN(n164) );
  NR2D0 U242 ( .A1(net7585), .A2(net7581), .ZN(n633) );
  CKAN2D1 U243 ( .A1(n713), .A2(n55), .Z(n457) );
  CKAN2D1 U244 ( .A1(n174), .A2(n705), .Z(n458) );
  CKAN2D1 U245 ( .A1(n35), .A2(n461), .Z(n459) );
  CKAN2D1 U246 ( .A1(n43), .A2(n59), .Z(n460) );
  NR3D0 U247 ( .A1(n459), .A2(n460), .A3(n627), .ZN(n629) );
  OAI22D1 U248 ( .A1(n122), .A2(n651), .B1(n596), .B2(n675), .ZN(n597) );
  ND2D0 U249 ( .A1(net7585), .A2(net7259), .ZN(n190) );
  BUFFD4 U250 ( .I(a[0]), .Z(net7589) );
  NR2D0 U251 ( .A1(n57), .A2(n71), .ZN(n254) );
  CKND2D0 U252 ( .A1(n668), .A2(n675), .ZN(n555) );
  AOI21D1 U253 ( .A1(n716), .A2(n48), .B(n714), .ZN(n536) );
  ND2D0 U254 ( .A1(n34), .A2(net7259), .ZN(n626) );
  OAI31D1 U255 ( .A1(n623), .A2(n46), .A3(n65), .B(n197), .ZN(n624) );
  NR2D1 U256 ( .A1(n651), .A2(n157), .ZN(n661) );
  INVD1 U257 ( .I(n181), .ZN(n33) );
  NR2XD0 U258 ( .A1(n4), .A2(n359), .ZN(n490) );
  ND2D0 U259 ( .A1(net7581), .A2(n51), .ZN(n98) );
  CKND2D0 U260 ( .A1(n181), .A2(net12782), .ZN(n637) );
  BUFFD4 U261 ( .I(a[2]), .Z(net7587) );
  NR2D0 U262 ( .A1(n60), .A2(n64), .ZN(n484) );
  CKND0 U263 ( .I(n286), .ZN(n52) );
  ND3D0 U264 ( .A1(n48), .A2(n197), .A3(n19), .ZN(n686) );
  AOI22D0 U265 ( .A1(n716), .A2(n705), .B1(n47), .B2(n17), .ZN(n522) );
  ND2D0 U266 ( .A1(n49), .A2(net7255), .ZN(n662) );
  ND2D0 U267 ( .A1(n34), .A2(n5), .ZN(n628) );
  ND2D0 U268 ( .A1(n53), .A2(n10), .ZN(n535) );
  CKND2D0 U269 ( .A1(n43), .A2(n19), .ZN(n622) );
  ND2D0 U270 ( .A1(n461), .A2(n5), .ZN(n493) );
  NR2D0 U271 ( .A1(n661), .A2(n715), .ZN(n666) );
  CKND0 U272 ( .I(n663), .ZN(n711) );
  NR2D0 U273 ( .A1(n716), .A2(n17), .ZN(n474) );
  AOI21D0 U274 ( .A1(n708), .A2(n2), .B(n712), .ZN(n537) );
  AOI22D0 U275 ( .A1(n56), .A2(n6), .B1(n64), .B2(n27), .ZN(n538) );
  OAI33D0 U276 ( .A1(n111), .A2(net7573), .A3(n139), .B1(n212), .B2(net7255), 
        .B3(n611), .ZN(n614) );
  CKND2D0 U277 ( .A1(n84), .A2(n315), .ZN(n528) );
  NR2XD0 U278 ( .A1(n21), .A2(n10), .ZN(n619) );
  CKND1 U279 ( .I(n204), .ZN(n18) );
  CKND2D0 U280 ( .A1(n84), .A2(n182), .ZN(n499) );
  CKND2D0 U281 ( .A1(n142), .A2(n148), .ZN(n500) );
  OAI32D0 U282 ( .A1(n312), .A2(n63), .A3(n120), .B1(n494), .B2(n493), .ZN(
        n495) );
  CKND2D0 U283 ( .A1(n103), .A2(n106), .ZN(n681) );
  OAI31D0 U284 ( .A1(n675), .A2(n41), .A3(n115), .B(n674), .ZN(n679) );
  AOI31D0 U285 ( .A1(n16), .A2(n673), .A3(n41), .B(n672), .ZN(n674) );
  NR2D0 U286 ( .A1(n53), .A2(n60), .ZN(n463) );
  AOI32D0 U287 ( .A1(n64), .A2(n72), .A3(n31), .B1(n461), .B2(n524), .ZN(n526)
         );
  CKND2D0 U288 ( .A1(n116), .A2(n680), .ZN(n524) );
  CKND0 U289 ( .I(n116), .ZN(n41) );
  OAI22D0 U290 ( .A1(n123), .A2(n111), .B1(n566), .B2(n122), .ZN(n573) );
  NR2D0 U291 ( .A1(n709), .A2(n34), .ZN(n566) );
  OAI22D0 U292 ( .A1(n101), .A2(n182), .B1(n639), .B2(n157), .ZN(n468) );
  NR2D0 U293 ( .A1(n585), .A2(n123), .ZN(n689) );
  CKND2D0 U294 ( .A1(n36), .A2(n16), .ZN(n233) );
  CKND2D0 U295 ( .A1(net7573), .A2(n45), .ZN(n527) );
  CKND2D0 U296 ( .A1(n197), .A2(n16), .ZN(n557) );
  CKND2D0 U298 ( .A1(n304), .A2(n51), .ZN(n664) );
  CKND0 U299 ( .I(n164), .ZN(n2) );
  CKND2D0 U300 ( .A1(n633), .A2(n16), .ZN(n591) );
  CKND2D0 U301 ( .A1(n33), .A2(n16), .ZN(n104) );
  CKND0 U302 ( .I(net7255), .ZN(net8759) );
  CKND2D0 U303 ( .A1(n117), .A2(n16), .ZN(n570) );
  AOI21D0 U304 ( .A1(n706), .A2(n19), .B(n540), .ZN(n491) );
  NR2D0 U305 ( .A1(n55), .A2(net7585), .ZN(n577) );
  OAI22D0 U306 ( .A1(n120), .A2(n114), .B1(n101), .B2(n696), .ZN(n636) );
  AOI32D0 U307 ( .A1(net7581), .A2(n72), .A3(n47), .B1(n36), .B2(n593), .ZN(
        n594) );
  CKND0 U308 ( .I(n689), .ZN(n710) );
  NR2D0 U309 ( .A1(n55), .A2(n57), .ZN(n480) );
  CKND0 U310 ( .I(n673), .ZN(n707) );
  AOI31D0 U311 ( .A1(net7583), .A2(n30), .A3(n53), .B(n172), .ZN(n483) );
  CKND2D0 U312 ( .A1(n48), .A2(n45), .ZN(n567) );
  AOI211D0 U313 ( .A1(n46), .A2(net7589), .B(n48), .C(n55), .ZN(n568) );
  AOI21D0 U314 ( .A1(n17), .A2(n48), .B(n682), .ZN(n683) );
  OAI33D0 U315 ( .A1(n114), .A2(n115), .A3(n116), .B1(n93), .B2(net7573), .B3(
        net12782), .ZN(n682) );
  OAI33D0 U316 ( .A1(n226), .A2(net7579), .A3(n97), .B1(n164), .B2(net7573), 
        .B3(n116), .ZN(n510) );
  AOI21D0 U317 ( .A1(n8), .A2(net7255), .B(n174), .ZN(n642) );
  ND4D0 U318 ( .A1(n68), .A2(n28), .A3(net7583), .A4(net7579), .ZN(n667) );
  OAI21D0 U319 ( .A1(n115), .A2(n257), .B(n663), .ZN(n559) );
  OAI22D0 U320 ( .A1(net7579), .A2(n212), .B1(n116), .B2(n139), .ZN(n464) );
  NR2D0 U321 ( .A1(n715), .A2(n174), .ZN(n466) );
  AOI21D0 U322 ( .A1(n91), .A2(n680), .B(n86), .ZN(n587) );
  OAI22D0 U323 ( .A1(n696), .A2(n82), .B1(n83), .B2(n84), .ZN(n697) );
  OAI22D0 U324 ( .A1(n470), .A2(n86), .B1(n119), .B2(n233), .ZN(n471) );
  AOI21D0 U325 ( .A1(n182), .A2(n552), .B(n123), .ZN(n467) );
  AOI33D0 U326 ( .A1(n574), .A2(n30), .A3(n705), .B1(n10), .B2(n51), .B3(n461), 
        .ZN(n575) );
  OAI31D0 U327 ( .A1(n119), .A2(n90), .A3(net12782), .B(n575), .ZN(n580) );
  AOI211D0 U328 ( .A1(n90), .A2(n212), .B(n552), .C(n123), .ZN(n485) );
  OAI22D0 U329 ( .A1(n30), .A2(n157), .B1(n45), .B2(n212), .ZN(n604) );
  AOI21D0 U330 ( .A1(n715), .A2(n47), .B(n172), .ZN(n645) );
  CKND2D0 U331 ( .A1(net7587), .A2(n45), .ZN(n586) );
  OAI21D0 U332 ( .A1(n653), .A2(n675), .B(n652), .ZN(n656) );
  AOI21D0 U333 ( .A1(net7585), .A2(n5), .B(n46), .ZN(n690) );
  CKND2D0 U334 ( .A1(net11484), .A2(n675), .ZN(n673) );
  CKND2D0 U335 ( .A1(net12727), .A2(n51), .ZN(n542) );
  AOI22D0 U336 ( .A1(n709), .A2(n304), .B1(n41), .B2(net11484), .ZN(n541) );
  NR2D0 U337 ( .A1(n61), .A2(n706), .ZN(n543) );
  CKND2D1 U338 ( .A1(n563), .A2(n562), .ZN(n564) );
  CKND0 U339 ( .I(n231), .ZN(n11) );
  AOI32D0 U340 ( .A1(net7583), .A2(n25), .A3(n49), .B1(n48), .B2(n521), .ZN(
        n523) );
  OAI22D0 U341 ( .A1(a[6]), .A2(net7583), .B1(net7581), .B2(n63), .ZN(n521) );
  INVD1 U342 ( .I(n628), .ZN(n716) );
  INVD1 U343 ( .I(n83), .ZN(n17) );
  INVD1 U344 ( .I(n535), .ZN(n714) );
  ND2D1 U345 ( .A1(n197), .A2(n5), .ZN(n92) );
  INVD1 U346 ( .I(n103), .ZN(n60) );
  INVD1 U347 ( .I(n97), .ZN(n36) );
  INVD1 U348 ( .I(n233), .ZN(n8) );
  AO221D0 U349 ( .A1(n64), .A2(n31), .B1(n461), .B2(n49), .C(n648), .Z(n609)
         );
  NR2D1 U350 ( .A1(n48), .A2(n41), .ZN(n611) );
  INVD1 U351 ( .I(n232), .ZN(n10) );
  ND2D1 U352 ( .A1(n2), .A2(n40), .ZN(n82) );
  INVD1 U353 ( .I(n557), .ZN(n715) );
  INVD1 U354 ( .I(n591), .ZN(n713) );
  ND2D1 U355 ( .A1(n71), .A2(n709), .ZN(n270) );
  ND2D1 U356 ( .A1(n708), .A2(n28), .ZN(n649) );
  INVD1 U357 ( .I(n527), .ZN(n708) );
  INVD1 U358 ( .I(n570), .ZN(n712) );
  OAI222D0 U359 ( .A1(n142), .A2(net12782), .B1(n639), .B2(n181), .C1(n111), 
        .C2(n315), .ZN(n508) );
  NR4D0 U360 ( .A1(n157), .A2(n103), .A3(n63), .A4(n37), .ZN(n672) );
  OAI221D0 U361 ( .A1(n675), .A2(n182), .B1(n120), .B2(n650), .C(n635), .ZN(
        n641) );
  OAI222D0 U362 ( .A1(n666), .A2(n142), .B1(n665), .B2(n144), .C1(n664), .C2(
        n663), .ZN(n704) );
  AOI221D0 U363 ( .A1(n671), .A2(n49), .B1(n50), .B2(n670), .C(n669), .ZN(n703) );
  NR4D0 U364 ( .A1(n679), .A2(n678), .A3(n677), .A4(n676), .ZN(n702) );
  NR2D1 U365 ( .A1(n586), .A2(net12727), .ZN(n648) );
  NR4D0 U366 ( .A1(n546), .A2(n545), .A3(n544), .A4(n676), .ZN(n547) );
  INVD1 U367 ( .I(net12727), .ZN(n71) );
  NR4D0 U368 ( .A1(n614), .A2(n613), .A3(n612), .A4(n678), .ZN(n615) );
  NR2D1 U369 ( .A1(n580), .A2(n579), .ZN(n581) );
  OAI221D0 U370 ( .A1(n182), .A2(n626), .B1(n625), .B2(n696), .C(n624), .ZN(
        n627) );
  OAI221D0 U371 ( .A1(net7255), .A2(n622), .B1(n664), .B2(n628), .C(n501), 
        .ZN(n517) );
  NR4D0 U372 ( .A1(n656), .A2(n672), .A3(n655), .A4(n654), .ZN(n657) );
  OAI221D0 U373 ( .A1(n463), .A2(n257), .B1(n91), .B2(net12727), .C(n462), 
        .ZN(n473) );
  ND2D1 U374 ( .A1(n22), .A2(n36), .ZN(n663) );
  INR4D0 U375 ( .A1(n686), .B1(n498), .B2(n677), .B3(n654), .ZN(n519) );
  AOI211D1 U376 ( .A1(n2), .A2(n497), .B(n496), .C(n495), .ZN(n520) );
  INVD1 U377 ( .I(n91), .ZN(n49) );
  INVD1 U378 ( .I(n84), .ZN(n47) );
  NR3D0 U379 ( .A1(net12727), .A2(n45), .A3(n137), .ZN(n544) );
  INVD1 U380 ( .I(n101), .ZN(n32) );
  INVD1 U381 ( .I(n668), .ZN(n706) );
  ND2D1 U382 ( .A1(n633), .A2(n19), .ZN(n137) );
  NR3D0 U383 ( .A1(n360), .A2(n116), .A3(n696), .ZN(n486) );
  INVD1 U384 ( .I(n190), .ZN(n46) );
  INVD1 U385 ( .I(n144), .ZN(n21) );
  INVD1 U386 ( .I(n360), .ZN(n29) );
  ND2D1 U387 ( .A1(n705), .A2(n72), .ZN(n315) );
  INVD1 U388 ( .I(n142), .ZN(n65) );
  INVD1 U389 ( .I(n650), .ZN(n709) );
  INVD1 U390 ( .I(n115), .ZN(n19) );
  INVD1 U391 ( .I(net7259), .ZN(net7257) );
  NR4D0 U392 ( .A1(net7257), .A2(n25), .A3(n103), .A4(n111), .ZN(n643) );
  OAI222D0 U393 ( .A1(n148), .A2(n105), .B1(n639), .B2(n663), .C1(n638), .C2(
        n86), .ZN(n640) );
  AOI21D1 U394 ( .A1(n71), .A2(n604), .B(n603), .ZN(n607) );
  OAI222D0 U395 ( .A1(n492), .A2(n123), .B1(n491), .B2(n116), .C1(n490), .C2(
        n103), .ZN(n496) );
  OAI222D0 U396 ( .A1(net7579), .A2(n691), .B1(n690), .B2(n97), .C1(n86), .C2(
        n98), .ZN(n693) );
  OAI222D0 U397 ( .A1(n578), .A2(n92), .B1(n577), .B2(n144), .C1(n576), .C2(
        n111), .ZN(n579) );
  OAI222D0 U398 ( .A1(net12162), .A2(n630), .B1(n629), .B2(n115), .C1(n190), 
        .C2(n628), .ZN(n631) );
  INR4D0 U399 ( .A1(n622), .B1(n621), .B2(n620), .B3(n714), .ZN(n630) );
  NR4D0 U400 ( .A1(n508), .A2(n507), .A3(n506), .A4(n561), .ZN(n509) );
  NR3D0 U401 ( .A1(n675), .A2(net7585), .A3(n101), .ZN(n507) );
  OAI222D0 U402 ( .A1(n63), .A2(n586), .B1(net7585), .B2(n585), .C1(n115), 
        .C2(n98), .ZN(n589) );
  OAI222D0 U403 ( .A1(n148), .A2(n570), .B1(n569), .B2(net7573), .C1(n568), 
        .C2(n628), .ZN(n571) );
  NR2XD0 U404 ( .A1(n603), .A2(n689), .ZN(n569) );
  OAI221D0 U405 ( .A1(n675), .A2(n139), .B1(net7257), .B2(n83), .C(n667), .ZN(
        n670) );
  NR4D0 U406 ( .A1(n181), .A2(n114), .A3(n86), .A4(n45), .ZN(n612) );
  NR2D1 U407 ( .A1(net7583), .A2(n30), .ZN(n477) );
  OAI222D0 U408 ( .A1(n103), .A2(n104), .B1(n105), .B2(n106), .C1(net7255), 
        .C2(n686), .ZN(n699) );
  OAI222D0 U409 ( .A1(n120), .A2(n315), .B1(n226), .B2(net12727), .C1(n119), 
        .C2(n181), .ZN(n469) );
  NR3D0 U410 ( .A1(n675), .A2(net7583), .A3(n258), .ZN(n603) );
  NR4D0 U411 ( .A1(net12162), .A2(n30), .A3(n97), .A4(n91), .ZN(n545) );
  NR3D0 U412 ( .A1(n91), .A2(net7579), .A3(net7583), .ZN(n620) );
  ND2D1 U413 ( .A1(net7583), .A2(n51), .ZN(n157) );
  NR3D0 U414 ( .A1(n162), .A2(n37), .A3(n157), .ZN(n348) );
  AOI222D0 U415 ( .A1(n705), .A2(n43), .B1(n41), .B2(n60), .C1(n706), .C2(
        net7581), .ZN(n563) );
  NR3D0 U416 ( .A1(n662), .A2(net7583), .A3(n25), .ZN(n613) );
  OAI221D0 U417 ( .A1(n72), .A2(n135), .B1(n162), .B2(net12727), .C(n642), 
        .ZN(n647) );
  ND2D1 U418 ( .A1(net7583), .A2(net7587), .ZN(n650) );
  INVD1 U419 ( .I(net7587), .ZN(n66) );
  INVD1 U420 ( .I(n93), .ZN(n27) );
  INVD1 U421 ( .I(n90), .ZN(n26) );
  OAI222D0 U422 ( .A1(n232), .A2(net7573), .B1(n258), .B2(n567), .C1(net7585), 
        .C2(n663), .ZN(n572) );
  OAI211D0 U423 ( .A1(n37), .A2(n111), .B(n94), .C(n116), .ZN(n634) );
  OAI222D0 U424 ( .A1(n90), .A2(n696), .B1(n91), .B2(n92), .C1(n93), .C2(n94), 
        .ZN(n692) );
  OAI221D0 U425 ( .A1(n466), .A2(n226), .B1(n94), .B2(n135), .C(n465), .ZN(
        n472) );
  AOI32D0 U426 ( .A1(net7579), .A2(n45), .A3(n64), .B1(n59), .B2(n464), .ZN(
        n465) );
  AOI221D0 U427 ( .A1(n71), .A2(n50), .B1(net8948), .B2(n35), .C(n561), .ZN(
        n562) );
  NR2D1 U428 ( .A1(n693), .A2(n692), .ZN(n694) );
  AOI22D1 U429 ( .A1(n705), .A2(n28), .B1(n53), .B2(n45), .ZN(n691) );
  AN2D1 U430 ( .A1(net7589), .A2(n51), .Z(n623) );
  NR4D0 U431 ( .A1(n97), .A2(n63), .A3(net9018), .A4(net7585), .ZN(n676) );
  INR2D1 U432 ( .A1(n348), .B1(net9018), .ZN(n654) );
  NR2D1 U433 ( .A1(n360), .A2(net9018), .ZN(n540) );
  NR4D0 U434 ( .A1(n487), .A2(n486), .A3(n655), .A4(n485), .ZN(n488) );
  CKND2D1 U435 ( .A1(n57), .A2(n72), .ZN(n161) );
  NR3D0 U436 ( .A1(n72), .A2(net7583), .A3(n181), .ZN(n561) );
  OAI22D0 U437 ( .A1(net7585), .A2(n257), .B1(n72), .B2(n258), .ZN(n574) );
  OA21D0 U438 ( .A1(n182), .A2(n72), .B(n254), .Z(n578) );
  NR2D0 U439 ( .A1(n72), .A2(n686), .ZN(n678) );
  NR2D1 U440 ( .A1(n32), .A2(n53), .ZN(n494) );
  NR2D1 U441 ( .A1(n232), .A2(n664), .ZN(n677) );
  ND2D1 U442 ( .A1(n65), .A2(n32), .ZN(n602) );
  OAI22D1 U443 ( .A1(net8759), .A2(n663), .B1(net7255), .B2(n232), .ZN(n595)
         );
  NR3D0 U444 ( .A1(n623), .A2(n64), .A3(n49), .ZN(n605) );
  OAI32D0 U445 ( .A1(n98), .A2(n484), .A3(n162), .B1(n483), .B2(n675), .ZN(
        n487) );
  OA33D0 U446 ( .A1(n651), .A2(n116), .A3(n123), .B1(n161), .B2(n162), .B3(n98), .Z(n652) );
  OAI222D0 U447 ( .A1(n106), .A2(n98), .B1(n84), .B2(n602), .C1(net12782), 
        .C2(n161), .ZN(n610) );
  AOI22D0 U448 ( .A1(n28), .A2(n681), .B1(n26), .B2(n59), .ZN(n684) );
  AOI22D0 U449 ( .A1(n35), .A2(n59), .B1(n705), .B2(n33), .ZN(n462) );
  AOI22D0 U450 ( .A1(n26), .A2(n59), .B1(n56), .B2(n27), .ZN(n482) );
  AOI222D0 U451 ( .A1(n57), .A2(n40), .B1(n117), .B2(n65), .C1(n33), .C2(n59), 
        .ZN(n525) );
  NR3D0 U452 ( .A1(n37), .A2(net7257), .A3(n142), .ZN(n506) );
  AOI21D0 U453 ( .A1(n181), .A2(n101), .B(n142), .ZN(n632) );
  NR2D1 U454 ( .A1(n65), .A2(n68), .ZN(n639) );
  NR2XD0 U455 ( .A1(n31), .A2(n35), .ZN(n625) );
  AOI31D0 U456 ( .A1(n135), .A2(n136), .A3(n137), .B(n668), .ZN(n669) );
  AOI22D0 U457 ( .A1(n12), .A2(n500), .B1(n174), .B2(n499), .ZN(n501) );
  AOI21D0 U458 ( .A1(n136), .A2(n622), .B(net11484), .ZN(n588) );
endmodule


module aes_sbox_5 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n65, n70, n114, n304, n305, n306, n310, n313, n404, n405, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864;

  AN2XD1 U28 ( .A1(n721), .A2(n720), .Z(n725) );
  OA21D1 U35 ( .A1(n705), .A2(n704), .B(n703), .Z(n710) );
  OR3D1 U88 ( .A1(n430), .A2(n812), .A3(n451), .Z(n633) );
  OA21D1 U101 ( .A1(n686), .A2(n795), .B(n614), .Z(n618) );
  OR4D1 U199 ( .A1(n657), .A2(n575), .A3(n524), .A4(n523), .Z(n526) );
  MAOI22D1 U209 ( .A1(n858), .A2(n814), .B1(n626), .B2(n774), .ZN(n517) );
  AN2XD1 U215 ( .A1(n525), .A2(n810), .Z(n524) );
  AO21D1 U297 ( .A1(n798), .A2(n836), .B(n736), .Z(n465) );
  OAI222D2 U1 ( .A1(n432), .A2(n635), .B1(n590), .B2(n589), .C1(n758), .C2(
        n588), .ZN(n591) );
  OAI222D1 U2 ( .A1(n477), .A2(n708), .B1(n470), .B2(n706), .C1(n729), .C2(
        n730), .ZN(n474) );
  ND4D2 U3 ( .A1(n662), .A2(n663), .A3(n661), .A4(n660), .ZN(d[2]) );
  ND3D2 U4 ( .A1(n549), .A2(n548), .A3(n547), .ZN(d[5]) );
  OAI22D1 U5 ( .A1(n451), .A2(n631), .B1(n630), .B2(n745), .ZN(n632) );
  CKND2D1 U6 ( .A1(n812), .A2(n449), .ZN(n582) );
  AOI211XD1 U7 ( .A1(n440), .A2(n587), .B(n585), .C(n586), .ZN(n588) );
  AOI221D2 U8 ( .A1(n851), .A2(n810), .B1(n694), .B2(n803), .C(n681), .ZN(n718) );
  INVD3 U9 ( .I(n451), .ZN(n450) );
  AOI31D1 U10 ( .A1(n443), .A2(n828), .A3(n798), .B(n827), .ZN(n498) );
  OAI222D1 U11 ( .A1(n784), .A2(n582), .B1(n776), .B2(n637), .C1(n499), .C2(
        n764), .ZN(n500) );
  NR4D0 U12 ( .A1(n536), .A2(n535), .A3(n534), .A4(n594), .ZN(n537) );
  AOI221D2 U13 ( .A1(n860), .A2(n645), .B1(n857), .B2(n803), .C(n644), .ZN(
        n662) );
  AOI222D1 U14 ( .A1(n803), .A2(n822), .B1(n824), .B2(n805), .C1(n807), .C2(
        n446), .ZN(n596) );
  OAI221D1 U15 ( .A1(n752), .A2(n426), .B1(n711), .B2(n786), .C(n634), .ZN(
        n645) );
  AOI221D1 U16 ( .A1(n836), .A2(n796), .B1(n592), .B2(n451), .C(n736), .ZN(
        n593) );
  INVD1 U17 ( .I(n746), .ZN(n65) );
  CKND2 U18 ( .I(n65), .ZN(n70) );
  CKND1 U19 ( .I(n65), .ZN(n114) );
  ND2D0 U20 ( .A1(n449), .A2(n444), .ZN(n783) );
  BUFFD4 U21 ( .I(a[2]), .Z(n443) );
  CKND2D1 U22 ( .A1(a[0]), .A2(n443), .ZN(n761) );
  INVD1 U23 ( .I(n758), .ZN(n860) );
  OR2D0 U24 ( .A1(a[0]), .A2(n443), .Z(n764) );
  AN2XD1 U25 ( .A1(n853), .A2(n818), .Z(n405) );
  ND2D1 U26 ( .A1(a[6]), .A2(n828), .ZN(n774) );
  ND2D1 U27 ( .A1(n444), .A2(n820), .ZN(n751) );
  ND2D1 U29 ( .A1(n450), .A2(a[0]), .ZN(n720) );
  CKND2D1 U30 ( .A1(n447), .A2(n828), .ZN(n729) );
  CKND2D1 U31 ( .A1(n795), .A2(n451), .ZN(n746) );
  NR2D1 U32 ( .A1(n704), .A2(n70), .ZN(n736) );
  ND2D1 U33 ( .A1(n443), .A2(n451), .ZN(n665) );
  INVD1 U34 ( .I(n611), .ZN(n831) );
  INVD3 U36 ( .I(n443), .ZN(n800) );
  ND2D1 U37 ( .A1(n444), .A2(n828), .ZN(n748) );
  AOI221D0 U38 ( .A1(n837), .A2(n825), .B1(n823), .B2(n571), .C(n852), .ZN(
        n499) );
  CKBD4 U39 ( .I(a[7]), .Z(n447) );
  ND2D1 U40 ( .A1(n444), .A2(n800), .ZN(n773) );
  ND2D1 U41 ( .A1(n683), .A2(n846), .ZN(n731) );
  AOI221D0 U42 ( .A1(n804), .A2(n834), .B1(n829), .B2(n559), .C(n702), .ZN(
        n564) );
  ND2D2 U43 ( .A1(n800), .A2(n814), .ZN(n686) );
  ND2D1 U44 ( .A1(n450), .A2(n443), .ZN(n749) );
  ND2D1 U45 ( .A1(n445), .A2(n444), .ZN(n752) );
  ND2D2 U46 ( .A1(n447), .A2(n835), .ZN(n758) );
  AOI221D0 U47 ( .A1(n796), .A2(n815), .B1(n802), .B2(n440), .C(n594), .ZN(
        n595) );
  ND2D2 U48 ( .A1(n447), .A2(a[6]), .ZN(n706) );
  INVD1 U49 ( .I(n776), .ZN(n816) );
  ND2D1 U50 ( .A1(n843), .A2(n829), .ZN(n722) );
  INVD1 U51 ( .I(n781), .ZN(n843) );
  OAI222D0 U52 ( .A1(n811), .A2(n631), .B1(n558), .B2(n538), .C1(n537), .C2(
        n781), .ZN(n544) );
  AOI221D1 U53 ( .A1(n801), .A2(n859), .B1(n810), .B2(n838), .C(n465), .ZN(
        n469) );
  ND2D1 U54 ( .A1(n828), .A2(n835), .ZN(n656) );
  INVD1 U55 ( .I(n753), .ZN(n846) );
  AOI21D1 U56 ( .A1(n862), .A2(n817), .B(n856), .ZN(n566) );
  INVD1 U57 ( .I(n773), .ZN(n812) );
  ND4D3 U58 ( .A1(n580), .A2(n581), .A3(n579), .A4(n578), .ZN(d[4]) );
  NR2D1 U59 ( .A1(n834), .A2(n830), .ZN(n674) );
  AOI21D4 U60 ( .A1(n815), .A2(n449), .B(n804), .ZN(n583) );
  AOI222D1 U61 ( .A1(n808), .A2(n825), .B1(n823), .B2(n442), .C1(n832), .C2(
        n806), .ZN(n555) );
  INVD0 U62 ( .I(n687), .ZN(n832) );
  AOI211XD0 U63 ( .A1(n863), .A2(n522), .B(n521), .C(n520), .ZN(n549) );
  OAI32D2 U64 ( .A1(n584), .A2(n114), .A3(n687), .B1(n583), .B2(n766), .ZN(
        n585) );
  ND2D1 U65 ( .A1(n803), .A2(n795), .ZN(n558) );
  INVD1 U66 ( .I(n678), .ZN(n819) );
  INVD1 U67 ( .I(n726), .ZN(n442) );
  INVD4 U68 ( .I(a[0]), .ZN(n795) );
  AN2XD1 U69 ( .A1(n451), .A2(n800), .Z(n304) );
  AN3XD1 U70 ( .A1(n623), .A2(n622), .A3(n621), .Z(n305) );
  AOI221D2 U71 ( .A1(n813), .A2(n571), .B1(n570), .B2(n823), .C(n569), .ZN(
        n579) );
  ND2D1 U72 ( .A1(a[0]), .A2(n800), .ZN(n726) );
  CKND2D1 U73 ( .A1(n443), .A2(n814), .ZN(n776) );
  BUFFD6 U74 ( .I(a[3]), .Z(n444) );
  CKND2D1 U75 ( .A1(n446), .A2(n814), .ZN(n769) );
  OAI22D1 U76 ( .A1(n795), .A2(n722), .B1(n451), .B2(n733), .ZN(n530) );
  OAI221D1 U77 ( .A1(n740), .A2(n733), .B1(n706), .B2(n114), .C(n593), .ZN(
        n601) );
  ND2D1 U78 ( .A1(n444), .A2(n443), .ZN(n642) );
  ND2D1 U79 ( .A1(n445), .A2(n828), .ZN(n611) );
  INVD6 U80 ( .I(n446), .ZN(n828) );
  ND2D2 U81 ( .A1(n801), .A2(a[0]), .ZN(n560) );
  INVD4 U82 ( .I(n424), .ZN(n801) );
  AOI21D0 U83 ( .A1(n834), .A2(n843), .B(n852), .ZN(n666) );
  CKND2D1 U84 ( .A1(n814), .A2(n820), .ZN(n756) );
  INVD2 U85 ( .I(a[6]), .ZN(n835) );
  AOI221D1 U86 ( .A1(n846), .A2(n463), .B1(n462), .B2(n795), .C(n461), .ZN(
        n484) );
  ND2D1 U87 ( .A1(n444), .A2(n451), .ZN(n678) );
  OAI22D1 U89 ( .A1(n114), .A2(n708), .B1(n639), .B2(n740), .ZN(n640) );
  INR4D1 U90 ( .A1(n670), .B1(n856), .B2(n668), .B3(n669), .ZN(n680) );
  OA22D1 U91 ( .A1(n665), .A2(n446), .B1(n611), .B2(n642), .Z(n561) );
  INVD4 U92 ( .I(n444), .ZN(n814) );
  AO31D1 U93 ( .A1(n803), .A2(n860), .A3(n683), .B(n719), .Z(n466) );
  INVD0 U94 ( .I(n560), .ZN(n802) );
  OAI222D1 U95 ( .A1(n782), .A2(n781), .B1(n444), .B2(n841), .C1(n780), .C2(
        n795), .ZN(n788) );
  OAI22D0 U96 ( .A1(n472), .A2(n711), .B1(n471), .B2(n761), .ZN(n473) );
  OAI222D1 U97 ( .A1(n568), .A2(n711), .B1(n567), .B2(n745), .C1(n449), .C2(
        n566), .ZN(n569) );
  NR3D1 U98 ( .A1(n404), .A2(n405), .A3(n466), .ZN(n468) );
  ND2D0 U99 ( .A1(n443), .A2(n446), .ZN(n747) );
  CKND2D1 U100 ( .A1(n445), .A2(n443), .ZN(n705) );
  INVD1 U102 ( .I(n304), .ZN(n425) );
  CKND2D0 U103 ( .A1(n443), .A2(n820), .ZN(n626) );
  CKND2D1 U104 ( .A1(n446), .A2(n835), .ZN(n513) );
  AOI221D1 U105 ( .A1(n799), .A2(n689), .B1(n834), .B2(n441), .C(n688), .ZN(
        n690) );
  AOI211XD0 U106 ( .A1(n844), .A2(a[0]), .B(n638), .C(n854), .ZN(n643) );
  OAI31D2 U107 ( .A1(n672), .A2(n442), .A3(n819), .B(n671), .ZN(n673) );
  OA221D1 U108 ( .A1(n795), .A2(n306), .B1(n781), .B2(n310), .C(n313), .Z(n580) );
  OA211D0 U109 ( .A1(n704), .A2(n678), .B(n553), .C(n552), .Z(n306) );
  OA211D0 U110 ( .A1(n557), .A2(n720), .B(n556), .C(n555), .Z(n310) );
  OA222D1 U111 ( .A1(n564), .A2(n758), .B1(n563), .B2(n686), .C1(n562), .C2(
        n753), .Z(n313) );
  CKND2D2 U112 ( .A1(a[6]), .A2(n840), .ZN(n781) );
  ND2D1 U113 ( .A1(a[0]), .A2(n451), .ZN(n745) );
  INVD2 U114 ( .I(n745), .ZN(n798) );
  ND2D1 U115 ( .A1(n445), .A2(n814), .ZN(n711) );
  INVD1 U116 ( .I(n711), .ZN(n825) );
  OAI222D1 U117 ( .A1(n533), .A2(n776), .B1(n437), .B2(n625), .C1(n532), .C2(
        n720), .ZN(n545) );
  CKND2 U118 ( .I(n304), .ZN(n424) );
  OAI222D1 U119 ( .A1(n732), .A2(n721), .B1(n699), .B2(n795), .C1(n698), .C2(
        n774), .ZN(n700) );
  NR2XD0 U120 ( .A1(n808), .A2(n796), .ZN(n614) );
  CKND2D2 U121 ( .A1(n449), .A2(n795), .ZN(n740) );
  ND2D2 U122 ( .A1(n853), .A2(n795), .ZN(n637) );
  AOI22D1 U123 ( .A1(n795), .A2(n818), .B1(n814), .B2(n805), .ZN(n590) );
  AOI221D1 U124 ( .A1(n848), .A2(n795), .B1(n858), .B2(n449), .C(n640), .ZN(
        n641) );
  NR4D1 U125 ( .A1(n544), .A2(n545), .A3(n546), .A4(n543), .ZN(n547) );
  AOI211XD1 U126 ( .A1(n804), .A2(n824), .B(n827), .C(n697), .ZN(n698) );
  AOI221D1 U127 ( .A1(n861), .A2(n795), .B1(n853), .B2(n808), .C(n632), .ZN(
        n663) );
  AOI221D2 U128 ( .A1(n802), .A2(n851), .B1(n796), .B2(n864), .C(n591), .ZN(
        n624) );
  INVD0 U129 ( .I(n752), .ZN(n824) );
  AOI221D1 U130 ( .A1(n798), .A2(n684), .B1(n683), .B2(n806), .C(n682), .ZN(
        n685) );
  OAI221D1 U131 ( .A1(n686), .A2(n675), .B1(n674), .B2(n786), .C(n673), .ZN(
        n676) );
  OAI221D1 U132 ( .A1(n667), .A2(n678), .B1(n666), .B2(n431), .C(n847), .ZN(
        n669) );
  ND2D0 U133 ( .A1(a[0]), .A2(n806), .ZN(n730) );
  AOI211XD0 U134 ( .A1(n819), .A2(a[0]), .B(n817), .C(n810), .ZN(n604) );
  NR2XD1 U135 ( .A1(n442), .A2(n798), .ZN(n691) );
  OA222D1 U136 ( .A1(n469), .A2(n751), .B1(n687), .B2(n518), .C1(n468), .C2(
        n795), .Z(n436) );
  CKND2D1 U137 ( .A1(n444), .A2(n446), .ZN(n687) );
  CKND0 U138 ( .I(n114), .ZN(n797) );
  AOI221D1 U139 ( .A1(n846), .A2(n609), .B1(n608), .B2(n795), .C(n607), .ZN(
        n622) );
  INVD1 U140 ( .I(n751), .ZN(n823) );
  OA221D1 U141 ( .A1(n751), .A2(n438), .B1(n687), .B2(n749), .C(n439), .Z(n562) );
  AOI222D1 U142 ( .A1(n808), .A2(n831), .B1(n806), .B2(n487), .C1(n802), .C2(
        n834), .ZN(n492) );
  INVD2 U143 ( .I(n786), .ZN(n803) );
  ND2D2 U144 ( .A1(n450), .A2(n800), .ZN(n786) );
  AOI221D1 U145 ( .A1(n843), .A2(n501), .B1(n802), .B2(n514), .C(n500), .ZN(
        n510) );
  AOI221D1 U146 ( .A1(n816), .A2(n601), .B1(n843), .B2(n600), .C(n599), .ZN(
        n623) );
  OAI222D1 U147 ( .A1(n643), .A2(n432), .B1(n761), .B2(n763), .C1(n641), .C2(
        n773), .ZN(n644) );
  ND2D2 U148 ( .A1(n831), .A2(n849), .ZN(n732) );
  INVD4 U149 ( .I(n706), .ZN(n849) );
  OAI33D0 U150 ( .A1(n425), .A2(n753), .A3(n752), .B1(n774), .B2(n448), .B3(
        n751), .ZN(n754) );
  OAI21D0 U151 ( .A1(n656), .A2(n751), .B(n731), .ZN(n541) );
  NR2XD0 U152 ( .A1(n795), .A2(n444), .ZN(n430) );
  NR2D0 U153 ( .A1(n444), .A2(n446), .ZN(n683) );
  NR2XD0 U154 ( .A1(n795), .A2(n444), .ZN(n672) );
  INVD6 U155 ( .I(n447), .ZN(n840) );
  OAI21D0 U156 ( .A1(n753), .A2(n434), .B(n722), .ZN(n592) );
  OAI222D1 U157 ( .A1(a[0]), .A2(n680), .B1(n753), .B2(n679), .C1(n678), .C2(
        n677), .ZN(n681) );
  AOI221D1 U158 ( .A1(n823), .A2(n860), .B1(n812), .B2(n833), .C(n531), .ZN(
        n532) );
  INVD4 U159 ( .I(n445), .ZN(n820) );
  CKND2D2 U160 ( .A1(n446), .A2(n820), .ZN(n766) );
  ND2D3 U161 ( .A1(n835), .A2(n840), .ZN(n753) );
  ND2D1 U162 ( .A1(n846), .A2(n833), .ZN(n784) );
  ND2D1 U163 ( .A1(n822), .A2(n846), .ZN(n670) );
  CKND3 U164 ( .I(a[1]), .ZN(n451) );
  INVD4 U165 ( .I(n451), .ZN(n449) );
  AOI32D0 U166 ( .A1(n446), .A2(n795), .A3(n818), .B1(n829), .B2(n633), .ZN(
        n634) );
  CKND1 U167 ( .I(n729), .ZN(n859) );
  CKND2D1 U168 ( .A1(n446), .A2(n447), .ZN(n704) );
  ND2D0 U169 ( .A1(n446), .A2(a[6]), .ZN(n777) );
  AN2D1 U170 ( .A1(n445), .A2(n446), .Z(n671) );
  CKAN2D1 U171 ( .A1(n467), .A2(n808), .Z(n404) );
  ND4D2 U172 ( .A1(n718), .A2(n717), .A3(n716), .A4(n715), .ZN(d[1]) );
  AOI221D1 U173 ( .A1(n857), .A2(n796), .B1(n860), .B2(n693), .C(n692), .ZN(
        n717) );
  AOI221D1 U174 ( .A1(n801), .A2(n825), .B1(n809), .B2(n832), .C(n767), .ZN(
        n782) );
  AOI221D1 U175 ( .A1(n702), .A2(n859), .B1(n817), .B2(n701), .C(n700), .ZN(
        n716) );
  ND4D2 U176 ( .A1(n484), .A2(n483), .A3(n482), .A4(n481), .ZN(d[7]) );
  CKND0 U177 ( .I(n304), .ZN(n426) );
  NR4D1 U178 ( .A1(n788), .A2(n789), .A3(n790), .A4(n787), .ZN(n791) );
  CKND2D0 U179 ( .A1(n831), .A2(n451), .ZN(n675) );
  OAI22D0 U180 ( .A1(n766), .A2(n776), .B1(n449), .B2(n765), .ZN(n767) );
  AOI22D0 U181 ( .A1(n812), .A2(n833), .B1(n815), .B2(n828), .ZN(n765) );
  CKND2D0 U182 ( .A1(n799), .A2(n860), .ZN(n518) );
  AOI221D1 U183 ( .A1(n440), .A2(n799), .B1(n822), .B2(n806), .C(n676), .ZN(
        n679) );
  ND2D0 U184 ( .A1(n831), .A2(n860), .ZN(n677) );
  CKND2D0 U185 ( .A1(n836), .A2(n825), .ZN(n538) );
  ND2D0 U186 ( .A1(n812), .A2(n855), .ZN(n565) );
  NR2XD0 U187 ( .A1(n838), .A2(n849), .ZN(n639) );
  INVD0 U188 ( .I(n642), .ZN(n817) );
  CKND2D1 U189 ( .A1(n494), .A2(n493), .ZN(n495) );
  AOI21D0 U190 ( .A1(n858), .A2(n818), .B(n696), .ZN(n699) );
  OAI22D0 U191 ( .A1(n447), .A2(n656), .B1(n752), .B2(n729), .ZN(n454) );
  OA31D0 U192 ( .A1(n706), .A2(n446), .A3(n449), .B(n637), .Z(n429) );
  ND2D0 U193 ( .A1(n449), .A2(a[6]), .ZN(n488) );
  NR2D0 U194 ( .A1(n817), .A2(n824), .ZN(n655) );
  CKND0 U195 ( .I(n610), .ZN(n842) );
  AOI21D1 U196 ( .A1(n821), .A2(n863), .B(n850), .ZN(n567) );
  INVD1 U197 ( .I(n761), .ZN(n810) );
  ND2D1 U198 ( .A1(n820), .A2(n828), .ZN(n770) );
  CKND2D0 U200 ( .A1(n829), .A2(n849), .ZN(n635) );
  CKND2D0 U201 ( .A1(n730), .A2(n740), .ZN(n587) );
  NR2D0 U202 ( .A1(n625), .A2(n745), .ZN(n768) );
  CKND0 U203 ( .I(n764), .ZN(n805) );
  NR2XD0 U204 ( .A1(n861), .A2(n514), .ZN(n515) );
  BUFFD6 U205 ( .I(a[5]), .Z(n446) );
  BUFFD6 U206 ( .I(a[4]), .Z(n445) );
  NR2D0 U207 ( .A1(n795), .A2(n760), .ZN(n743) );
  AOI22D0 U208 ( .A1(n862), .A2(n803), .B1(n818), .B2(n848), .ZN(n552) );
  CKND2D0 U210 ( .A1(n863), .A2(n825), .ZN(n785) );
  CKND2D0 U211 ( .A1(n816), .A2(n449), .ZN(n721) );
  NR2D0 U212 ( .A1(n636), .A2(n723), .ZN(n742) );
  NR2D0 U213 ( .A1(n805), .A2(n801), .ZN(n477) );
  ND2D0 U214 ( .A1(n823), .A2(n863), .ZN(n762) );
  OAI21D0 U216 ( .A1(n432), .A2(n732), .B(n785), .ZN(n475) );
  CKND0 U217 ( .I(n775), .ZN(n861) );
  CKND0 U218 ( .I(n724), .ZN(n844) );
  NR2D0 U219 ( .A1(n719), .A2(n858), .ZN(n727) );
  CKND2D0 U220 ( .A1(n441), .A2(n833), .ZN(n646) );
  NR2D0 U221 ( .A1(n833), .A2(n812), .ZN(n519) );
  OAI33D0 U222 ( .A1(n756), .A2(n448), .A3(n729), .B1(n656), .B2(n449), .B3(
        n655), .ZN(n659) );
  NR2XD0 U223 ( .A1(n844), .A2(n855), .ZN(n667) );
  CKND1 U224 ( .I(n664), .ZN(n847) );
  CKND2D0 U225 ( .A1(n783), .A2(n686), .ZN(n527) );
  OAI22D0 U226 ( .A1(n432), .A2(n745), .B1(n114), .B2(n773), .ZN(n502) );
  OAI31D0 U227 ( .A1(n740), .A2(n824), .A3(n753), .B(n739), .ZN(n744) );
  AOI31D0 U228 ( .A1(n849), .A2(n738), .A3(n824), .B(n737), .ZN(n739) );
  NR2D0 U229 ( .A1(n812), .A2(n805), .ZN(n453) );
  OAI21D0 U230 ( .A1(n752), .A2(n610), .B(n635), .ZN(n514) );
  CKND2D0 U231 ( .A1(n828), .A2(n840), .ZN(n610) );
  AOI32D0 U232 ( .A1(n801), .A2(n795), .A3(n834), .B1(n799), .B2(n554), .ZN(
        n556) );
  CKND2D0 U233 ( .A1(n752), .A2(n747), .ZN(n554) );
  OAI22D0 U234 ( .A1(n745), .A2(n756), .B1(n602), .B2(n114), .ZN(n609) );
  NR2D0 U235 ( .A1(n826), .A2(n831), .ZN(n602) );
  OAI211D0 U236 ( .A1(n828), .A2(n756), .B(n773), .C(n752), .ZN(n684) );
  CKAN2D1 U237 ( .A1(n538), .A2(n733), .Z(n471) );
  AOI21D0 U238 ( .A1(n434), .A2(n656), .B(n686), .ZN(n503) );
  CKND2D0 U239 ( .A1(n764), .A2(n761), .ZN(n750) );
  AOI31D0 U240 ( .A1(n733), .A2(n732), .A3(n731), .B(n730), .ZN(n734) );
  NR2D0 U241 ( .A1(n513), .A2(n431), .ZN(n570) );
  INR2D0 U242 ( .A1(n525), .B1(n431), .ZN(n712) );
  CKND2D0 U243 ( .A1(n683), .A2(n849), .ZN(n631) );
  CKND2D0 U244 ( .A1(n797), .A2(n814), .ZN(n723) );
  AOI22D0 U245 ( .A1(n809), .A2(n859), .B1(n801), .B2(n838), .ZN(n568) );
  CKND0 U246 ( .I(n704), .ZN(n863) );
  CKND2D0 U247 ( .A1(n832), .A2(n849), .ZN(n763) );
  CKND2D0 U248 ( .A1(n823), .A2(n849), .ZN(n606) );
  OAI31D0 U249 ( .A1(n814), .A2(n804), .A3(n810), .B(n694), .ZN(n494) );
  OAI31D0 U250 ( .A1(n801), .A2(n798), .A3(n812), .B(n861), .ZN(n493) );
  NR2D0 U251 ( .A1(n862), .A2(n848), .ZN(n464) );
  OA221D0 U252 ( .A1(n451), .A2(n435), .B1(n598), .B2(n656), .C(n436), .Z(n483) );
  AOI21D0 U253 ( .A1(n796), .A2(n648), .B(n647), .ZN(n651) );
  NR2D0 U254 ( .A1(n810), .A2(n444), .ZN(n617) );
  AOI22D0 U255 ( .A1(n808), .A2(a[0]), .B1(n449), .B2(n817), .ZN(n486) );
  AOI21D0 U256 ( .A1(n823), .A2(n859), .B(n696), .ZN(n506) );
  CKND2D0 U257 ( .A1(n720), .A2(n814), .ZN(n573) );
  NR2D0 U258 ( .A1(n804), .A2(n807), .ZN(n574) );
  AOI22D0 U259 ( .A1(n826), .A2(n797), .B1(n824), .B2(n443), .ZN(n572) );
  CKND0 U260 ( .I(n738), .ZN(n811) );
  AOI211XD0 U261 ( .A1(n842), .A2(n809), .B(n490), .C(n489), .ZN(n491) );
  OAI21D0 U262 ( .A1(a[0]), .A2(n687), .B(n751), .ZN(n487) );
  AOI22D0 U263 ( .A1(n803), .A2(n837), .B1(n812), .B2(n820), .ZN(n772) );
  AOI211D0 U264 ( .A1(n864), .A2(n809), .B(n485), .C(n664), .ZN(n512) );
  CKND2D0 U265 ( .A1(n817), .A2(n820), .ZN(n603) );
  NR2XD0 U266 ( .A1(n647), .A2(n768), .ZN(n605) );
  CKND2D0 U267 ( .A1(n687), .A2(n751), .ZN(n689) );
  ND4D0 U268 ( .A1(n798), .A2(n837), .A3(n445), .A4(n447), .ZN(n728) );
  OAI22D0 U269 ( .A1(n786), .A2(n785), .B1(n784), .B2(n783), .ZN(n787) );
  OAI32D0 U270 ( .A1(n433), .A2(n477), .A3(n706), .B1(n476), .B2(n740), .ZN(
        n480) );
  AOI31D0 U271 ( .A1(n445), .A2(n835), .A3(n812), .B(n696), .ZN(n476) );
  AOI21D0 U272 ( .A1(n776), .A2(n747), .B(n781), .ZN(n627) );
  AOI21D0 U273 ( .A1(n732), .A2(n670), .B(n443), .ZN(n628) );
  NR2D0 U274 ( .A1(n858), .A2(n694), .ZN(n456) );
  OAI31D0 U275 ( .A1(n749), .A2(n777), .A3(n751), .B(n613), .ZN(n620) );
  AOI33D0 U276 ( .A1(n612), .A2(n835), .A3(n803), .B1(n855), .B2(n814), .B3(
        n799), .ZN(n613) );
  OAI22D0 U277 ( .A1(n444), .A2(n434), .B1(n795), .B2(n610), .ZN(n612) );
  AOI211D0 U278 ( .A1(n777), .A2(n656), .B(n584), .C(n745), .ZN(n478) );
  OAI22D0 U279 ( .A1(n451), .A2(n722), .B1(n449), .B2(n636), .ZN(n638) );
  NR2D0 U280 ( .A1(n732), .A2(n444), .ZN(n696) );
  OAI22D0 U281 ( .A1(n460), .A2(n781), .B1(n749), .B2(n635), .ZN(n461) );
  OAI22D0 U282 ( .A1(n766), .A2(n686), .B1(n691), .B2(n711), .ZN(n458) );
  AOI21D0 U283 ( .A1(n686), .A2(n584), .B(n745), .ZN(n457) );
  NR2D0 U284 ( .A1(n760), .A2(a[0]), .ZN(n713) );
  CKND2D0 U285 ( .A1(n443), .A2(n740), .ZN(n738) );
  OAI21D0 U286 ( .A1(n710), .A2(n740), .B(n709), .ZN(n714) );
  CKND2D0 U287 ( .A1(n446), .A2(n840), .ZN(n708) );
  CKND2D1 U288 ( .A1(n596), .A2(n595), .ZN(n600) );
  AOI21D0 U289 ( .A1(n848), .A2(n817), .B(n754), .ZN(n755) );
  CKND2D1 U290 ( .A1(n774), .A2(n729), .ZN(n571) );
  CKND1 U291 ( .I(n797), .ZN(n438) );
  NR2D0 U292 ( .A1(n810), .A2(n808), .ZN(n470) );
  AOI21D0 U293 ( .A1(n807), .A2(n846), .B(n570), .ZN(n516) );
  CKND2D0 U294 ( .A1(n694), .A2(n114), .ZN(n427) );
  NR2D0 U295 ( .A1(n445), .A2(n835), .ZN(n467) );
  OAI33D0 U296 ( .A1(n656), .A2(a[0]), .A3(n448), .B1(n488), .B2(n729), .B3(
        n761), .ZN(n489) );
  AOI32D0 U298 ( .A1(n445), .A2(n840), .A3(n816), .B1(n817), .B2(n551), .ZN(
        n553) );
  CKND2D2 U299 ( .A1(n624), .A2(n305), .ZN(d[3]) );
  INVD1 U300 ( .I(n740), .ZN(n799) );
  INVD1 U301 ( .I(n784), .ZN(n848) );
  INVD1 U302 ( .I(n677), .ZN(n862) );
  INVD1 U303 ( .I(n707), .ZN(n809) );
  INVD1 U304 ( .I(n785), .ZN(n864) );
  INVD1 U305 ( .I(n565), .ZN(n856) );
  INVD1 U306 ( .I(n582), .ZN(n813) );
  OAI222D0 U307 ( .A1(n432), .A2(n724), .B1(n590), .B2(n733), .C1(n636), .C2(
        n431), .ZN(n485) );
  INVD1 U308 ( .I(n686), .ZN(n815) );
  INVD1 U309 ( .I(n589), .ZN(n858) );
  NR2D1 U310 ( .A1(n441), .A2(n797), .ZN(n615) );
  INVD1 U311 ( .I(n756), .ZN(n822) );
  INVD1 U312 ( .I(n770), .ZN(n829) );
  INVD1 U313 ( .I(n635), .ZN(n857) );
  INVD1 U314 ( .I(n631), .ZN(n851) );
  INVD1 U315 ( .I(n557), .ZN(n821) );
  INVD1 U316 ( .I(n597), .ZN(n852) );
  ND2D1 U317 ( .A1(n796), .A2(n826), .ZN(n598) );
  ND2D1 U318 ( .A1(n821), .A2(n837), .ZN(n703) );
  AO221D0 U319 ( .A1(n801), .A2(n834), .B1(n799), .B2(n816), .C(n702), .Z(n653) );
  INVD1 U320 ( .I(n732), .ZN(n853) );
  INVD1 U321 ( .I(n636), .ZN(n855) );
  ND2D1 U322 ( .A1(n808), .A2(n795), .ZN(n707) );
  INVD1 U323 ( .I(n722), .ZN(n845) );
  INVD1 U324 ( .I(n606), .ZN(n850) );
  OAI221D0 U325 ( .A1(n740), .A2(n686), .B1(n748), .B2(n705), .C(n685), .ZN(
        n693) );
  AOI221D0 U326 ( .A1(n862), .A2(n451), .B1(n844), .B2(n720), .C(n530), .ZN(
        n533) );
  OAI222D0 U327 ( .A1(n747), .A2(n720), .B1(n770), .B2(n582), .C1(n752), .C2(
        n761), .ZN(n586) );
  NR4D0 U328 ( .A1(n711), .A2(n764), .A3(n758), .A4(n828), .ZN(n737) );
  NR4D0 U329 ( .A1(n659), .A2(n658), .A3(n657), .A4(n743), .ZN(n660) );
  NR4D0 U330 ( .A1(n577), .A2(n576), .A3(n575), .A4(n741), .ZN(n578) );
  AOI221D0 U331 ( .A1(n812), .A2(n845), .B1(n853), .B2(n818), .C(n550), .ZN(
        n581) );
  OAI221D0 U332 ( .A1(n453), .A2(n434), .B1(n776), .B2(n720), .C(n452), .ZN(
        n463) );
  NR2D1 U333 ( .A1(n626), .A2(n720), .ZN(n702) );
  INVD1 U334 ( .I(n720), .ZN(n796) );
  AOI221D0 U335 ( .A1(n475), .A2(n451), .B1(n822), .B2(n474), .C(n473), .ZN(
        n482) );
  IND4D1 U336 ( .A1(n794), .B1(n793), .B2(n792), .B3(n791), .ZN(d[0]) );
  NR4D0 U337 ( .A1(n744), .A2(n743), .A3(n742), .A4(n741), .ZN(n792) );
  AOI221D0 U338 ( .A1(n736), .A2(n816), .B1(n815), .B2(n735), .C(n734), .ZN(
        n793) );
  ND2D1 U339 ( .A1(n849), .A2(n833), .ZN(n636) );
  OAI221D0 U340 ( .A1(n449), .A2(n670), .B1(n723), .B2(n677), .C(n529), .ZN(
        n546) );
  NR2D1 U341 ( .A1(n620), .A2(n619), .ZN(n621) );
  NR4D0 U342 ( .A1(n714), .A2(n737), .A3(n713), .A4(n712), .ZN(n715) );
  INR4D0 U343 ( .A1(n760), .B1(n526), .B2(n742), .B3(n712), .ZN(n548) );
  NR3D0 U344 ( .A1(n720), .A2(n820), .A3(n731), .ZN(n575) );
  INVD1 U345 ( .I(n783), .ZN(n818) );
  ND2D1 U346 ( .A1(n831), .A2(n843), .ZN(n724) );
  NR2D1 U347 ( .A1(n708), .A2(n711), .ZN(n719) );
  NR3D0 U348 ( .A1(n513), .A2(n752), .A3(n786), .ZN(n479) );
  INVD1 U349 ( .I(n766), .ZN(n833) );
  INVD1 U350 ( .I(n749), .ZN(n808) );
  INVD1 U351 ( .I(n705), .ZN(n826) );
  INVD1 U352 ( .I(n730), .ZN(n807) );
  INVD1 U353 ( .I(n665), .ZN(n806) );
  ND2D1 U354 ( .A1(n830), .A2(n849), .ZN(n597) );
  INVD1 U355 ( .I(n769), .ZN(n834) );
  INVD1 U356 ( .I(n558), .ZN(n804) );
  INVD1 U357 ( .I(n513), .ZN(n836) );
  OAI222D0 U358 ( .A1(n425), .A2(n606), .B1(n605), .B2(n448), .C1(n604), .C2(
        n677), .ZN(n607) );
  OAI222D0 U359 ( .A1(n437), .A2(n538), .B1(n492), .B2(n753), .C1(n491), .C2(
        n756), .ZN(n496) );
  NR4D0 U360 ( .A1(n450), .A2(n840), .A3(n764), .A4(n756), .ZN(n697) );
  OAI222D0 U361 ( .A1(n636), .A2(n448), .B1(n610), .B2(n603), .C1(n444), .C2(
        n722), .ZN(n608) );
  OAI222D0 U362 ( .A1(n447), .A2(n772), .B1(n771), .B2(n770), .C1(n781), .C2(
        n433), .ZN(n779) );
  NR3D0 U363 ( .A1(n740), .A2(n444), .A3(n766), .ZN(n535) );
  OAI222D0 U364 ( .A1(n758), .A2(n626), .B1(n444), .B2(n625), .C1(n753), .C2(
        n433), .ZN(n629) );
  OAI222D0 U365 ( .A1(n764), .A2(n763), .B1(n762), .B2(n761), .C1(n449), .C2(
        n760), .ZN(n789) );
  OAI222D0 U366 ( .A1(n759), .A2(n758), .B1(n757), .B2(n756), .C1(a[0]), .C2(
        n755), .ZN(n790) );
  OAI221D0 U367 ( .A1(n456), .A2(n432), .B1(n773), .B2(n733), .C(n455), .ZN(
        n462) );
  OAI222D0 U368 ( .A1(n517), .A2(n745), .B1(n516), .B2(n752), .C1(n515), .C2(
        n764), .ZN(n521) );
  OAI222D0 U369 ( .A1(n449), .A2(n777), .B1(n114), .B2(n758), .C1(n753), .C2(
        n749), .ZN(n490) );
  OAI222D0 U370 ( .A1(n777), .A2(n786), .B1(n776), .B2(n775), .C1(n774), .C2(
        n773), .ZN(n778) );
  OAI222D0 U371 ( .A1(n426), .A2(n762), .B1(n691), .B2(n722), .C1(n690), .C2(
        n781), .ZN(n692) );
  OAI222D0 U372 ( .A1(n618), .A2(n775), .B1(n617), .B2(n724), .C1(n616), .C2(
        n756), .ZN(n619) );
  OA22D0 U373 ( .A1(n777), .A2(n745), .B1(n729), .B2(n615), .Z(n616) );
  INVD1 U374 ( .I(n768), .ZN(n841) );
  NR2XD0 U375 ( .A1(n779), .A2(n778), .ZN(n780) );
  OAI221D0 U376 ( .A1(n610), .A2(n584), .B1(n444), .B2(n775), .C(n703), .ZN(
        n531) );
  OAI222D0 U377 ( .A1(n506), .A2(n114), .B1(n820), .B2(n505), .C1(n504), .C2(
        n720), .ZN(n508) );
  ND2D1 U378 ( .A1(n447), .A2(n502), .ZN(n505) );
  INR2D1 U379 ( .A1(n762), .B1(n503), .ZN(n504) );
  OAI222D0 U380 ( .A1(n574), .A2(n775), .B1(n784), .B2(n573), .C1(n572), .C2(
        n777), .ZN(n577) );
  NR3D0 U381 ( .A1(n795), .A2(n445), .A3(n687), .ZN(n594) );
  OAI222D0 U382 ( .A1(n443), .A2(n651), .B1(n650), .B2(n785), .C1(n649), .C2(
        n784), .ZN(n652) );
  OAI221D0 U383 ( .A1(n795), .A2(n733), .B1(n706), .B2(n720), .C(n695), .ZN(
        n701) );
  AOI21D1 U384 ( .A1(n857), .A2(n449), .B(n694), .ZN(n695) );
  NR4D0 U385 ( .A1(n770), .A2(n758), .A3(n431), .A4(n444), .ZN(n741) );
  ND4D1 U386 ( .A1(n512), .A2(n511), .A3(n510), .A4(n509), .ZN(d[6]) );
  NR4D0 U387 ( .A1(n508), .A2(n507), .A3(n523), .A4(n524), .ZN(n509) );
  AOI211XD0 U388 ( .A1(n860), .A2(n497), .B(n496), .C(n495), .ZN(n511) );
  OAI221D0 U389 ( .A1(n615), .A2(n766), .B1(n752), .B2(n761), .C(n498), .ZN(
        n501) );
  NR4D0 U390 ( .A1(n459), .A2(n458), .A3(n534), .A4(n457), .ZN(n460) );
  NR4D0 U391 ( .A1(n629), .A2(n628), .A3(n850), .A4(n627), .ZN(n630) );
  NR3D0 U392 ( .A1(n740), .A2(n445), .A3(n610), .ZN(n647) );
  INVD1 U393 ( .I(n637), .ZN(n854) );
  NR4D0 U394 ( .A1(a[0]), .A2(n835), .A3(n770), .A4(n776), .ZN(n576) );
  NR3D0 U395 ( .A1(n776), .A2(n447), .A3(n445), .ZN(n668) );
  OAI221D0 U396 ( .A1(n740), .A2(n729), .B1(n450), .B2(n784), .C(n728), .ZN(
        n735) );
  AN3XD1 U397 ( .A1(n427), .A2(n428), .A3(n429), .Z(n563) );
  ND2D0 U398 ( .A1(n449), .A2(n855), .ZN(n428) );
  NR3D0 U399 ( .A1(n706), .A2(n828), .A3(n711), .ZN(n525) );
  NR3D0 U400 ( .A1(n721), .A2(n445), .A3(n840), .ZN(n658) );
  OAI222D0 U401 ( .A1(n426), .A2(n687), .B1(n486), .B2(n766), .C1(n449), .C2(
        n752), .ZN(n497) );
  INVD1 U402 ( .I(n774), .ZN(n838) );
  INVD1 U403 ( .I(n777), .ZN(n839) );
  NR4D0 U404 ( .A1(a[6]), .A2(n814), .A3(n729), .A4(n761), .ZN(n507) );
  OAI222D0 U405 ( .A1(n707), .A2(n733), .B1(a[0]), .B2(n542), .C1(n786), .C2(
        n775), .ZN(n543) );
  CKBD1 U406 ( .I(n665), .Z(n431) );
  INVD1 U407 ( .I(n817), .ZN(n432) );
  INVD1 U408 ( .I(n748), .ZN(n830) );
  CKND2D0 U409 ( .A1(n445), .A2(n800), .ZN(n584) );
  OAI33D0 U410 ( .A1(n642), .A2(n447), .A3(n770), .B1(n704), .B2(n800), .B3(
        n752), .ZN(n539) );
  ND2D0 U411 ( .A1(n800), .A2(n820), .ZN(n557) );
  INVD1 U412 ( .I(n834), .ZN(n433) );
  AOI221D0 U413 ( .A1(n806), .A2(n541), .B1(n846), .B2(n540), .C(n539), .ZN(
        n542) );
  AOI22D1 U414 ( .A1(n839), .A2(n806), .B1(n809), .B2(n838), .ZN(n472) );
  AOI22D0 U415 ( .A1(n440), .A2(n806), .B1(n803), .B2(n832), .ZN(n452) );
  AOI22D1 U416 ( .A1(n837), .A2(n750), .B1(n839), .B2(n806), .ZN(n757) );
  AOI32D0 U417 ( .A1(n447), .A2(n820), .A3(n801), .B1(n806), .B2(n454), .ZN(
        n455) );
  NR2D1 U418 ( .A1(n797), .A2(n806), .ZN(n650) );
  AOI221D1 U419 ( .A1(n843), .A2(n654), .B1(n846), .B2(n653), .C(n652), .ZN(
        n661) );
  ND2D1 U420 ( .A1(n833), .A2(n840), .ZN(n625) );
  AOI21D0 U421 ( .A1(n444), .A2(n860), .B(n819), .ZN(n771) );
  OAI222D0 U422 ( .A1(n748), .A2(n558), .B1(n642), .B2(n720), .C1(n749), .C2(
        n687), .ZN(n459) );
  OA222D0 U423 ( .A1(n749), .A2(n748), .B1(n747), .B2(n114), .C1(n751), .C2(
        n745), .Z(n759) );
  OAI32D0 U424 ( .A1(n560), .A2(n758), .A3(n748), .B1(n519), .B2(n518), .ZN(
        n520) );
  CKBD0 U425 ( .I(n611), .Z(n434) );
  OA221D0 U426 ( .A1(n464), .A2(n776), .B1(n722), .B2(n773), .C(n565), .Z(n435) );
  INVD1 U427 ( .I(n598), .ZN(n827) );
  INVD1 U428 ( .I(n656), .ZN(n837) );
  CKBD0 U429 ( .I(n800), .Z(n448) );
  OAI22D0 U430 ( .A1(n835), .A2(n711), .B1(n820), .B2(n656), .ZN(n648) );
  INVD1 U431 ( .I(n441), .ZN(n437) );
  AN4D1 U432 ( .A1(n671), .A2(n818), .A3(a[0]), .A4(n846), .Z(n523) );
  ND2D1 U433 ( .A1(n671), .A2(n860), .ZN(n775) );
  ND3D0 U434 ( .A1(n817), .A2(n671), .A3(n846), .ZN(n760) );
  ND2D1 U435 ( .A1(n671), .A2(n849), .ZN(n589) );
  ND2D1 U436 ( .A1(n843), .A2(n671), .ZN(n733) );
  OAI22D0 U437 ( .A1(n756), .A2(n425), .B1(n655), .B2(n740), .ZN(n522) );
  NR4D0 U438 ( .A1(n687), .A2(n425), .A3(n781), .A4(n820), .ZN(n657) );
  OAI22D0 U439 ( .A1(n748), .A2(n425), .B1(n766), .B2(n786), .ZN(n688) );
  OAI22D1 U440 ( .A1(n724), .A2(n426), .B1(n800), .B2(n731), .ZN(n664) );
  OA222D1 U441 ( .A1(n665), .A2(n769), .B1(a[0]), .B2(n561), .C1(n752), .C2(
        n560), .Z(n439) );
  NR4D0 U442 ( .A1(n480), .A2(n479), .A3(n713), .A4(n478), .ZN(n481) );
  AOI22D0 U443 ( .A1(n853), .A2(n528), .B1(n694), .B2(n527), .ZN(n529) );
  OAI22D0 U444 ( .A1(a[6]), .A2(n445), .B1(n446), .B2(n758), .ZN(n551) );
  OAI211D0 U445 ( .A1(n446), .A2(n783), .B(n626), .C(n751), .ZN(n540) );
  CKND2D0 U446 ( .A1(n783), .A2(n558), .ZN(n559) );
  CKND0 U447 ( .I(n748), .ZN(n440) );
  OAI222D0 U448 ( .A1(n727), .A2(n437), .B1(n725), .B2(n724), .C1(n723), .C2(
        n722), .ZN(n794) );
  AOI21D0 U449 ( .A1(n687), .A2(n766), .B(n726), .ZN(n682) );
  OAI222D0 U450 ( .A1(n729), .A2(n598), .B1(n437), .B2(n763), .C1(n614), .C2(
        n597), .ZN(n599) );
  OAI222D0 U451 ( .A1(n437), .A2(n597), .B1(n733), .B2(n678), .C1(n636), .C2(
        n761), .ZN(n550) );
  OAI222D0 U452 ( .A1(n437), .A2(n751), .B1(n691), .B2(n687), .C1(n756), .C2(
        n558), .ZN(n536) );
  CKND2D0 U453 ( .A1(n437), .A2(n426), .ZN(n528) );
  NR3D0 U454 ( .A1(n828), .A2(n450), .A3(n437), .ZN(n534) );
  CKND0 U455 ( .I(n726), .ZN(n441) );
  OA33D0 U456 ( .A1(n708), .A2(n752), .A3(n745), .B1(n707), .B2(n706), .B3(
        n433), .Z(n709) );
  OAI222D0 U457 ( .A1(n761), .A2(n433), .B1(n783), .B2(n646), .C1(n751), .C2(
        n707), .ZN(n654) );
  NR3D0 U458 ( .A1(n430), .A2(n801), .A3(n816), .ZN(n649) );
  NR2XD0 U459 ( .A1(n753), .A2(n770), .ZN(n694) );
endmodule


module aes_cipher_top ( clk, rst, ld, done, key, text_in, text_out, SE, SI, SO
 );
  input [127:0] key;
  input [127:0] text_in;
  output [127:0] text_out;
  input clk, rst, ld, SE, SI;
  output done, SO;
  wire   N12, N13, N14, N15, N16, N21, ld_r, N32, N33, N34, N35, N36, N37, N38,
         N39, N48, N49, N50, N51, N52, N53, N54, N55, N64, N65, N66, N67, N68,
         N69, N70, N71, N80, N81, N82, N83, N84, N85, N86, N87, N96, N97, N98,
         N99, N100, N101, N102, N103, N112, N113, N114, N115, N116, N117, N118,
         N119, N128, N129, N130, N131, N132, N133, N134, N135, N144, N145,
         N146, N147, N148, N149, N150, N151, N160, N161, N162, N163, N164,
         N165, N166, N167, N176, N177, N178, N179, N180, N181, N182, N183,
         N192, N193, N194, N195, N196, N197, N198, N199, N208, N209, N210,
         N211, N212, N213, N214, N215, N224, N225, N226, N227, N228, N229,
         N230, N231, N240, N241, N242, N243, N244, N245, N246, N247, N256,
         N257, N258, N259, N260, N261, N262, N263, N272, N273, N274, N275,
         N276, N277, N278, N279, N376, N377, N378, N379, N380, N381, N382,
         N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393,
         N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404,
         N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415,
         N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, N426,
         N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437,
         N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470,
         N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481,
         N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492,
         N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, n1,
         n2, n3, n6, n8, n9, n10, n12, n13, n14, n15, n16, n18, n20, n21, n22,
         n23, n24, n25, n26, n27, n31, n32, n34, n35, n37, n38, n39, n40, n42,
         n44, n45, n47, n48, n54, n55, n56, n57, n58, n59, n60, n61, n62, n66,
         n67, n68, n69, n70, n72, n75, n76, n78, n79, n80, n81, n82, n84, n85,
         n87, n88, n90, n91, n92, n93, n95, n96, n97, n98, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n126, n127,
         n128, n129, n131, n132, n133, n134, n135, n136, n139, n140, n141,
         n143, n144, n146, n147, n148, n150, n151, n152, n155, n156, n157,
         n159, n160, n163, n164, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n185, n186, n187, n188, n189, n190, n191, n192, n194, n198, n200,
         n203, n204, n205, n206, n207, n209, n211, n212, n214, n215, n216,
         n217, n219, n220, n221, n222, n223, n224, n225, n226, n228, n229,
         n230, n231, n233, n234, n235, n236, n237, n238, n239, n241, n242,
         n243, n245, n246, n248, n250, n251, n253, n254, n255, n257, n258,
         n259, n262, n263, n265, n266, n268, n269, n270, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n284, n285, n286,
         n287, n288, n289, n291, n293, n294, n296, n298, n299, n300, n302,
         n305, n306, n307, n308, n309, n311, n314, n316, n317, n318, n319,
         n321, n322, n323, n324, n325, n326, n327, n328, n330, n331, n332,
         n333, n335, n336, n337, n338, n339, n340, n341, n342, n344, n345,
         n346, n348, n349, n351, n353, n354, n356, n357, n360, n361, n362,
         n363, n364, n365, n368, n369, n371, n372, n373, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n387, n388, n389,
         n390, n391, n392, n393, n394, n396, n397, n399, n401, n402, n403,
         n405, n408, n409, n411, n412, n413, n414, n416, n417, n419, n420,
         n421, n422, n423, n424, n425, n427, n428, n429, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n442, n443, n444, n445,
         n446, n448, n449, n450, n451, n452, n453, n454, n455, n457, n458,
         n460, n461, n462, n464, n465, n466, n467, n468, n469, n470, n472,
         n474, n475, n477, n478, n479, n481, n482, n485, n488, n489, n490,
         n491, n492, n493, n494, n497, n498, n499, n500, n502, n503, n504,
         n506, n507, n508, n509, net7025, net7023, net7021, net7019, net7017,
         net7015, net7013, net7011, net7009, net7007, net7005, net7003,
         net7001, net6999, net6997, net6995, net6993, net6991, net7033,
         net7031, net7029, net7027, n196, n149, n11, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713;
  wire   [3:0] dcnt;
  wire   [127:0] text_in_r;
  wire   [31:0] w3;
  wire   [7:0] sa33;
  wire   [7:0] sa23;
  wire   [7:0] sa13;
  wire   [7:0] sa03;
  wire   [31:0] w2;
  wire   [7:0] sa32;
  wire   [7:0] sa22;
  wire   [7:0] sa12;
  wire   [7:0] sa02;
  wire   [31:0] w1;
  wire   [7:0] sa31;
  wire   [7:0] sa21;
  wire   [7:0] sa11;
  wire   [7:0] sa01;
  wire   [31:0] w0;
  wire   [7:0] sa30;
  wire   [7:0] sa20;
  wire   [7:0] sa10;
  wire   [7:0] sa00;
  wire   [7:0] sa00_sr;
  wire   [7:0] sa01_sr;
  wire   [7:0] sa02_sr;
  wire   [7:0] sa03_sr;
  wire   [7:0] sa10_sr;
  wire   [7:0] sa11_sr;
  wire   [7:0] sa12_sr;
  wire   [7:0] sa13_sr;
  wire   [7:0] sa20_sr;
  wire   [7:0] sa21_sr;
  wire   [7:0] sa22_sr;
  wire   [7:0] sa23_sr;
  wire   [7:0] sa30_sr;
  wire   [7:0] sa31_sr;
  wire   [7:0] sa32_sr;
  wire   [7:0] sa33_sr;

  aes_key_expand_128 u0 ( .clk(clk), .kld(ld), .key(key), .wo_0(w0), .wo_1(w1), 
        .wo_2(w2), .wo_3(w3) );
  aes_sbox_0 us00 ( .a(sa00), .d(sa00_sr) );
  aes_sbox_19 us01 ( .a(sa01), .d(sa01_sr) );
  aes_sbox_18 us02 ( .a(sa02), .d(sa02_sr) );
  aes_sbox_17 us03 ( .a(sa03), .d(sa03_sr) );
  aes_sbox_16 us10 ( .a(sa10), .d(sa13_sr) );
  aes_sbox_15 us11 ( .a(sa11), .d(sa10_sr) );
  aes_sbox_14 us12 ( .a(sa12), .d(sa11_sr) );
  aes_sbox_13 us13 ( .a(sa13), .d(sa12_sr) );
  aes_sbox_12 us20 ( .a(sa20), .d(sa22_sr) );
  aes_sbox_11 us21 ( .a(sa21), .d(sa23_sr) );
  aes_sbox_10 us22 ( .a(sa22), .d(sa20_sr) );
  aes_sbox_9 us23 ( .a(sa23), .d(sa21_sr) );
  aes_sbox_8 us30 ( .a(sa30), .d(sa31_sr) );
  aes_sbox_7 us31 ( .a(sa31), .d(sa32_sr) );
  aes_sbox_6 us32 ( .a(sa32), .d(sa33_sr) );
  aes_sbox_5 us33 ( .a(sa33), .d(sa30_sr) );
  EDFQD1 dcnt_reg_0_ ( .D(N13), .E(N12), .CP(clk), .Q(dcnt[0]) );
  EDFQD1 dcnt_reg_3_ ( .D(N16), .E(N12), .CP(clk), .Q(dcnt[3]) );
  EDFQD1 dcnt_reg_2_ ( .D(N15), .E(N12), .CP(clk), .Q(dcnt[2]) );
  EDFQD1 dcnt_reg_1_ ( .D(N14), .E(N12), .CP(clk), .Q(dcnt[1]) );
  DFQD1 done_reg ( .D(N21), .CP(clk), .Q(done) );
  EDFQD1 text_in_r_reg_127_ ( .D(text_in[127]), .E(ld), .CP(clk), .Q(
        text_in_r[127]) );
  EDFQD1 text_in_r_reg_126_ ( .D(text_in[126]), .E(ld), .CP(clk), .Q(
        text_in_r[126]) );
  EDFQD1 text_in_r_reg_125_ ( .D(text_in[125]), .E(ld), .CP(clk), .Q(
        text_in_r[125]) );
  EDFQD1 text_in_r_reg_124_ ( .D(text_in[124]), .E(ld), .CP(clk), .Q(
        text_in_r[124]) );
  EDFQD1 text_in_r_reg_123_ ( .D(text_in[123]), .E(ld), .CP(clk), .Q(
        text_in_r[123]) );
  EDFQD1 text_in_r_reg_122_ ( .D(text_in[122]), .E(ld), .CP(clk), .Q(
        text_in_r[122]) );
  EDFQD1 text_in_r_reg_121_ ( .D(text_in[121]), .E(ld), .CP(clk), .Q(
        text_in_r[121]) );
  EDFQD1 text_in_r_reg_120_ ( .D(text_in[120]), .E(ld), .CP(clk), .Q(
        text_in_r[120]) );
  EDFQD1 text_in_r_reg_119_ ( .D(text_in[119]), .E(ld), .CP(clk), .Q(
        text_in_r[119]) );
  EDFQD1 text_in_r_reg_118_ ( .D(text_in[118]), .E(ld), .CP(clk), .Q(
        text_in_r[118]) );
  EDFQD1 text_in_r_reg_117_ ( .D(text_in[117]), .E(ld), .CP(clk), .Q(
        text_in_r[117]) );
  EDFQD1 text_in_r_reg_116_ ( .D(text_in[116]), .E(ld), .CP(clk), .Q(
        text_in_r[116]) );
  EDFQD1 text_in_r_reg_115_ ( .D(text_in[115]), .E(ld), .CP(clk), .Q(
        text_in_r[115]) );
  EDFQD1 text_in_r_reg_114_ ( .D(text_in[114]), .E(ld), .CP(clk), .Q(
        text_in_r[114]) );
  EDFQD1 text_in_r_reg_113_ ( .D(text_in[113]), .E(ld), .CP(clk), .Q(
        text_in_r[113]) );
  EDFQD1 text_in_r_reg_112_ ( .D(text_in[112]), .E(ld), .CP(clk), .Q(
        text_in_r[112]) );
  EDFQD1 text_in_r_reg_111_ ( .D(text_in[111]), .E(ld), .CP(clk), .Q(
        text_in_r[111]) );
  EDFQD1 text_in_r_reg_110_ ( .D(text_in[110]), .E(ld), .CP(clk), .Q(
        text_in_r[110]) );
  EDFQD1 text_in_r_reg_109_ ( .D(text_in[109]), .E(ld), .CP(clk), .Q(
        text_in_r[109]) );
  EDFQD1 text_in_r_reg_108_ ( .D(text_in[108]), .E(ld), .CP(clk), .Q(
        text_in_r[108]) );
  EDFQD1 text_in_r_reg_107_ ( .D(text_in[107]), .E(ld), .CP(clk), .Q(
        text_in_r[107]) );
  EDFQD1 text_in_r_reg_106_ ( .D(text_in[106]), .E(ld), .CP(clk), .Q(
        text_in_r[106]) );
  EDFQD1 text_in_r_reg_105_ ( .D(text_in[105]), .E(ld), .CP(clk), .Q(
        text_in_r[105]) );
  EDFQD1 text_in_r_reg_104_ ( .D(text_in[104]), .E(ld), .CP(clk), .Q(
        text_in_r[104]) );
  EDFQD1 text_in_r_reg_103_ ( .D(text_in[103]), .E(ld), .CP(clk), .Q(
        text_in_r[103]) );
  EDFQD1 text_in_r_reg_102_ ( .D(text_in[102]), .E(ld), .CP(clk), .Q(
        text_in_r[102]) );
  EDFQD1 text_in_r_reg_101_ ( .D(text_in[101]), .E(ld), .CP(clk), .Q(
        text_in_r[101]) );
  EDFQD1 text_in_r_reg_100_ ( .D(text_in[100]), .E(ld), .CP(clk), .Q(
        text_in_r[100]) );
  EDFQD1 text_in_r_reg_99_ ( .D(text_in[99]), .E(ld), .CP(clk), .Q(
        text_in_r[99]) );
  EDFQD1 text_in_r_reg_98_ ( .D(text_in[98]), .E(ld), .CP(clk), .Q(
        text_in_r[98]) );
  EDFQD1 text_in_r_reg_97_ ( .D(text_in[97]), .E(ld), .CP(clk), .Q(
        text_in_r[97]) );
  EDFQD1 text_in_r_reg_96_ ( .D(text_in[96]), .E(ld), .CP(clk), .Q(
        text_in_r[96]) );
  EDFQD1 text_in_r_reg_95_ ( .D(text_in[95]), .E(ld), .CP(clk), .Q(
        text_in_r[95]) );
  EDFQD1 text_in_r_reg_94_ ( .D(text_in[94]), .E(ld), .CP(clk), .Q(
        text_in_r[94]) );
  EDFQD1 text_in_r_reg_93_ ( .D(text_in[93]), .E(ld), .CP(clk), .Q(
        text_in_r[93]) );
  EDFQD1 text_in_r_reg_92_ ( .D(text_in[92]), .E(ld), .CP(clk), .Q(
        text_in_r[92]) );
  EDFQD1 text_in_r_reg_91_ ( .D(text_in[91]), .E(ld), .CP(clk), .Q(
        text_in_r[91]) );
  EDFQD1 text_in_r_reg_90_ ( .D(text_in[90]), .E(ld), .CP(clk), .Q(
        text_in_r[90]) );
  EDFQD1 text_in_r_reg_89_ ( .D(text_in[89]), .E(ld), .CP(clk), .Q(
        text_in_r[89]) );
  EDFQD1 text_in_r_reg_88_ ( .D(text_in[88]), .E(ld), .CP(clk), .Q(
        text_in_r[88]) );
  EDFQD1 text_in_r_reg_87_ ( .D(text_in[87]), .E(ld), .CP(clk), .Q(
        text_in_r[87]) );
  EDFQD1 text_in_r_reg_86_ ( .D(text_in[86]), .E(ld), .CP(clk), .Q(
        text_in_r[86]) );
  EDFQD1 text_in_r_reg_85_ ( .D(text_in[85]), .E(ld), .CP(clk), .Q(
        text_in_r[85]) );
  EDFQD1 text_in_r_reg_84_ ( .D(text_in[84]), .E(ld), .CP(clk), .Q(
        text_in_r[84]) );
  EDFQD1 text_in_r_reg_83_ ( .D(text_in[83]), .E(ld), .CP(clk), .Q(
        text_in_r[83]) );
  EDFQD1 text_in_r_reg_82_ ( .D(text_in[82]), .E(ld), .CP(clk), .Q(
        text_in_r[82]) );
  EDFQD1 text_in_r_reg_81_ ( .D(text_in[81]), .E(ld), .CP(clk), .Q(
        text_in_r[81]) );
  EDFQD1 text_in_r_reg_80_ ( .D(text_in[80]), .E(ld), .CP(clk), .Q(
        text_in_r[80]) );
  EDFQD1 text_in_r_reg_79_ ( .D(text_in[79]), .E(ld), .CP(clk), .Q(
        text_in_r[79]) );
  EDFQD1 text_in_r_reg_78_ ( .D(text_in[78]), .E(ld), .CP(clk), .Q(
        text_in_r[78]) );
  EDFQD1 text_in_r_reg_77_ ( .D(text_in[77]), .E(ld), .CP(clk), .Q(
        text_in_r[77]) );
  EDFQD1 text_in_r_reg_76_ ( .D(text_in[76]), .E(ld), .CP(clk), .Q(
        text_in_r[76]) );
  EDFQD1 text_in_r_reg_75_ ( .D(text_in[75]), .E(ld), .CP(clk), .Q(
        text_in_r[75]) );
  EDFQD1 text_in_r_reg_74_ ( .D(text_in[74]), .E(ld), .CP(clk), .Q(
        text_in_r[74]) );
  EDFQD1 text_in_r_reg_73_ ( .D(text_in[73]), .E(ld), .CP(clk), .Q(
        text_in_r[73]) );
  EDFQD1 text_in_r_reg_72_ ( .D(text_in[72]), .E(ld), .CP(clk), .Q(
        text_in_r[72]) );
  EDFQD1 text_in_r_reg_71_ ( .D(text_in[71]), .E(ld), .CP(clk), .Q(
        text_in_r[71]) );
  EDFQD1 text_in_r_reg_70_ ( .D(text_in[70]), .E(ld), .CP(clk), .Q(
        text_in_r[70]) );
  EDFQD1 text_in_r_reg_69_ ( .D(text_in[69]), .E(ld), .CP(clk), .Q(
        text_in_r[69]) );
  EDFQD1 text_in_r_reg_68_ ( .D(text_in[68]), .E(ld), .CP(clk), .Q(
        text_in_r[68]) );
  EDFQD1 text_in_r_reg_67_ ( .D(text_in[67]), .E(ld), .CP(clk), .Q(
        text_in_r[67]) );
  EDFQD1 text_in_r_reg_66_ ( .D(text_in[66]), .E(ld), .CP(clk), .Q(
        text_in_r[66]) );
  EDFQD1 text_in_r_reg_65_ ( .D(text_in[65]), .E(ld), .CP(clk), .Q(
        text_in_r[65]) );
  EDFQD1 text_in_r_reg_64_ ( .D(text_in[64]), .E(ld), .CP(clk), .Q(
        text_in_r[64]) );
  EDFQD1 text_in_r_reg_63_ ( .D(text_in[63]), .E(ld), .CP(clk), .Q(
        text_in_r[63]) );
  EDFQD1 text_in_r_reg_62_ ( .D(text_in[62]), .E(ld), .CP(clk), .Q(
        text_in_r[62]) );
  EDFQD1 text_in_r_reg_61_ ( .D(text_in[61]), .E(ld), .CP(clk), .Q(
        text_in_r[61]) );
  EDFQD1 text_in_r_reg_60_ ( .D(text_in[60]), .E(ld), .CP(clk), .Q(
        text_in_r[60]) );
  EDFQD1 text_in_r_reg_59_ ( .D(text_in[59]), .E(ld), .CP(clk), .Q(
        text_in_r[59]) );
  EDFQD1 text_in_r_reg_58_ ( .D(text_in[58]), .E(ld), .CP(clk), .Q(
        text_in_r[58]) );
  EDFQD1 text_in_r_reg_57_ ( .D(text_in[57]), .E(ld), .CP(clk), .Q(
        text_in_r[57]) );
  EDFQD1 text_in_r_reg_56_ ( .D(text_in[56]), .E(ld), .CP(clk), .Q(
        text_in_r[56]) );
  EDFQD1 text_in_r_reg_55_ ( .D(text_in[55]), .E(ld), .CP(clk), .Q(
        text_in_r[55]) );
  EDFQD1 text_in_r_reg_54_ ( .D(text_in[54]), .E(ld), .CP(clk), .Q(
        text_in_r[54]) );
  EDFQD1 text_in_r_reg_53_ ( .D(text_in[53]), .E(ld), .CP(clk), .Q(
        text_in_r[53]) );
  EDFQD1 text_in_r_reg_52_ ( .D(text_in[52]), .E(ld), .CP(clk), .Q(
        text_in_r[52]) );
  EDFQD1 text_in_r_reg_51_ ( .D(text_in[51]), .E(ld), .CP(clk), .Q(
        text_in_r[51]) );
  EDFQD1 text_in_r_reg_50_ ( .D(text_in[50]), .E(ld), .CP(clk), .Q(
        text_in_r[50]) );
  EDFQD1 text_in_r_reg_49_ ( .D(text_in[49]), .E(ld), .CP(clk), .Q(
        text_in_r[49]) );
  EDFQD1 text_in_r_reg_48_ ( .D(text_in[48]), .E(ld), .CP(clk), .Q(
        text_in_r[48]) );
  EDFQD1 text_in_r_reg_47_ ( .D(text_in[47]), .E(ld), .CP(clk), .Q(
        text_in_r[47]) );
  EDFQD1 text_in_r_reg_46_ ( .D(text_in[46]), .E(ld), .CP(clk), .Q(
        text_in_r[46]) );
  EDFQD1 text_in_r_reg_45_ ( .D(text_in[45]), .E(ld), .CP(clk), .Q(
        text_in_r[45]) );
  EDFQD1 text_in_r_reg_44_ ( .D(text_in[44]), .E(ld), .CP(clk), .Q(
        text_in_r[44]) );
  EDFQD1 text_in_r_reg_43_ ( .D(text_in[43]), .E(ld), .CP(clk), .Q(
        text_in_r[43]) );
  EDFQD1 text_in_r_reg_42_ ( .D(text_in[42]), .E(ld), .CP(clk), .Q(
        text_in_r[42]) );
  EDFQD1 text_in_r_reg_41_ ( .D(text_in[41]), .E(ld), .CP(clk), .Q(
        text_in_r[41]) );
  EDFQD1 text_in_r_reg_40_ ( .D(text_in[40]), .E(ld), .CP(clk), .Q(
        text_in_r[40]) );
  EDFQD1 text_in_r_reg_39_ ( .D(text_in[39]), .E(ld), .CP(clk), .Q(
        text_in_r[39]) );
  EDFQD1 text_in_r_reg_38_ ( .D(text_in[38]), .E(ld), .CP(clk), .Q(
        text_in_r[38]) );
  EDFQD1 text_in_r_reg_37_ ( .D(text_in[37]), .E(ld), .CP(clk), .Q(
        text_in_r[37]) );
  EDFQD1 text_in_r_reg_36_ ( .D(text_in[36]), .E(ld), .CP(clk), .Q(
        text_in_r[36]) );
  EDFQD1 text_in_r_reg_35_ ( .D(text_in[35]), .E(ld), .CP(clk), .Q(
        text_in_r[35]) );
  EDFQD1 text_in_r_reg_34_ ( .D(text_in[34]), .E(ld), .CP(clk), .Q(
        text_in_r[34]) );
  EDFQD1 text_in_r_reg_33_ ( .D(text_in[33]), .E(ld), .CP(clk), .Q(
        text_in_r[33]) );
  EDFQD1 text_in_r_reg_32_ ( .D(text_in[32]), .E(ld), .CP(clk), .Q(
        text_in_r[32]) );
  EDFQD1 text_in_r_reg_31_ ( .D(text_in[31]), .E(ld), .CP(clk), .Q(
        text_in_r[31]) );
  EDFQD1 text_in_r_reg_30_ ( .D(text_in[30]), .E(ld), .CP(clk), .Q(
        text_in_r[30]) );
  EDFQD1 text_in_r_reg_29_ ( .D(text_in[29]), .E(ld), .CP(clk), .Q(
        text_in_r[29]) );
  EDFQD1 text_in_r_reg_28_ ( .D(text_in[28]), .E(ld), .CP(clk), .Q(
        text_in_r[28]) );
  EDFQD1 text_in_r_reg_27_ ( .D(text_in[27]), .E(ld), .CP(clk), .Q(
        text_in_r[27]) );
  EDFQD1 text_in_r_reg_26_ ( .D(text_in[26]), .E(ld), .CP(clk), .Q(
        text_in_r[26]) );
  EDFQD1 text_in_r_reg_25_ ( .D(text_in[25]), .E(ld), .CP(clk), .Q(
        text_in_r[25]) );
  EDFQD1 text_in_r_reg_24_ ( .D(text_in[24]), .E(ld), .CP(clk), .Q(
        text_in_r[24]) );
  EDFQD1 text_in_r_reg_23_ ( .D(text_in[23]), .E(ld), .CP(clk), .Q(
        text_in_r[23]) );
  EDFQD1 text_in_r_reg_22_ ( .D(text_in[22]), .E(ld), .CP(clk), .Q(
        text_in_r[22]) );
  EDFQD1 text_in_r_reg_21_ ( .D(text_in[21]), .E(ld), .CP(clk), .Q(
        text_in_r[21]) );
  EDFQD1 text_in_r_reg_20_ ( .D(text_in[20]), .E(ld), .CP(clk), .Q(
        text_in_r[20]) );
  EDFQD1 text_in_r_reg_19_ ( .D(text_in[19]), .E(ld), .CP(clk), .Q(
        text_in_r[19]) );
  EDFQD1 text_in_r_reg_18_ ( .D(text_in[18]), .E(ld), .CP(clk), .Q(
        text_in_r[18]) );
  EDFQD1 text_in_r_reg_17_ ( .D(text_in[17]), .E(ld), .CP(clk), .Q(
        text_in_r[17]) );
  EDFQD1 text_in_r_reg_16_ ( .D(text_in[16]), .E(ld), .CP(clk), .Q(
        text_in_r[16]) );
  EDFQD1 text_in_r_reg_15_ ( .D(text_in[15]), .E(ld), .CP(clk), .Q(
        text_in_r[15]) );
  EDFQD1 text_in_r_reg_14_ ( .D(text_in[14]), .E(ld), .CP(clk), .Q(
        text_in_r[14]) );
  EDFQD1 text_in_r_reg_13_ ( .D(text_in[13]), .E(ld), .CP(clk), .Q(
        text_in_r[13]) );
  EDFQD1 text_in_r_reg_12_ ( .D(text_in[12]), .E(ld), .CP(clk), .Q(
        text_in_r[12]) );
  EDFQD1 text_in_r_reg_11_ ( .D(text_in[11]), .E(ld), .CP(clk), .Q(
        text_in_r[11]) );
  EDFQD1 text_in_r_reg_10_ ( .D(text_in[10]), .E(ld), .CP(clk), .Q(
        text_in_r[10]) );
  EDFQD1 text_in_r_reg_9_ ( .D(text_in[9]), .E(ld), .CP(clk), .Q(text_in_r[9])
         );
  EDFQD1 text_in_r_reg_8_ ( .D(text_in[8]), .E(ld), .CP(clk), .Q(text_in_r[8])
         );
  EDFQD1 text_in_r_reg_7_ ( .D(text_in[7]), .E(ld), .CP(clk), .Q(text_in_r[7])
         );
  EDFQD1 text_in_r_reg_6_ ( .D(text_in[6]), .E(ld), .CP(clk), .Q(text_in_r[6])
         );
  EDFQD1 text_in_r_reg_5_ ( .D(text_in[5]), .E(ld), .CP(clk), .Q(text_in_r[5])
         );
  EDFQD1 text_in_r_reg_4_ ( .D(text_in[4]), .E(ld), .CP(clk), .Q(text_in_r[4])
         );
  EDFQD1 text_in_r_reg_3_ ( .D(text_in[3]), .E(ld), .CP(clk), .Q(text_in_r[3])
         );
  EDFQD1 text_in_r_reg_2_ ( .D(text_in[2]), .E(ld), .CP(clk), .Q(text_in_r[2])
         );
  EDFQD1 text_in_r_reg_1_ ( .D(text_in[1]), .E(ld), .CP(clk), .Q(text_in_r[1])
         );
  EDFQD1 text_in_r_reg_0_ ( .D(text_in[0]), .E(ld), .CP(clk), .Q(text_in_r[0])
         );
  DFQD1 ld_r_reg ( .D(ld), .CP(clk), .Q(ld_r) );
  DFQD1 sa32_reg_4_ ( .D(N100), .CP(clk), .Q(sa32[4]) );
  DFQD1 sa20_reg_0_ ( .D(N240), .CP(clk), .Q(sa20[0]) );
  DFQD1 sa22_reg_7_ ( .D(N119), .CP(clk), .Q(sa22[7]) );
  DFQD1 sa21_reg_7_ ( .D(N183), .CP(clk), .Q(sa21[7]) );
  DFQD1 sa03_reg_7_ ( .D(N87), .CP(clk), .Q(sa03[7]) );
  DFQD1 sa13_reg_1_ ( .D(N65), .CP(clk), .Q(sa13[1]) );
  DFQD1 sa23_reg_2_ ( .D(N50), .CP(clk), .Q(sa23[2]) );
  DFQD1 sa03_reg_4_ ( .D(N84), .CP(clk), .Q(sa03[4]) );
  DFQD1 sa13_reg_3_ ( .D(N67), .CP(clk), .Q(sa13[3]) );
  DFQD1 sa03_reg_5_ ( .D(N85), .CP(clk), .Q(sa03[5]) );
  DFQD1 sa13_reg_4_ ( .D(N68), .CP(clk), .Q(sa13[4]) );
  DFQD1 sa13_reg_7_ ( .D(N71), .CP(clk), .Q(sa13[7]) );
  DFQD1 sa32_reg_0_ ( .D(N96), .CP(clk), .Q(sa32[0]) );
  DFQD1 sa12_reg_5_ ( .D(N133), .CP(clk), .Q(sa12[5]) );
  DFQD1 sa12_reg_0_ ( .D(N128), .CP(clk), .Q(sa12[0]) );
  DFQD1 sa31_reg_3_ ( .D(N163), .CP(clk), .Q(sa31[3]) );
  DFQD1 sa21_reg_4_ ( .D(N180), .CP(clk), .Q(sa21[4]) );
  DFQD1 sa21_reg_5_ ( .D(N181), .CP(clk), .Q(sa21[5]) );
  DFQD1 sa10_reg_4_ ( .D(N260), .CP(clk), .Q(sa10[4]) );
  DFQD1 sa20_reg_4_ ( .D(N244), .CP(clk), .Q(sa20[4]) );
  DFQD1 sa30_reg_4_ ( .D(N228), .CP(clk), .Q(sa30[4]) );
  DFQD1 sa20_reg_5_ ( .D(N245), .CP(clk), .Q(sa20[5]) );
  DFQD1 sa30_reg_6_ ( .D(N230), .CP(clk), .Q(sa30[6]) );
  DFQD1 sa00_reg_7_ ( .D(N279), .CP(clk), .Q(sa00[7]) );
  DFQD1 text_out_reg_127_ ( .D(N376), .CP(clk), .Q(text_out[127]) );
  DFQD1 text_out_reg_126_ ( .D(N377), .CP(clk), .Q(text_out[126]) );
  DFQD1 text_out_reg_125_ ( .D(N378), .CP(clk), .Q(text_out[125]) );
  DFQD1 text_out_reg_124_ ( .D(N379), .CP(clk), .Q(text_out[124]) );
  DFQD1 text_out_reg_123_ ( .D(N380), .CP(clk), .Q(text_out[123]) );
  DFQD1 text_out_reg_122_ ( .D(N381), .CP(clk), .Q(text_out[122]) );
  DFQD1 text_out_reg_121_ ( .D(N382), .CP(clk), .Q(text_out[121]) );
  DFQD1 text_out_reg_120_ ( .D(N383), .CP(clk), .Q(text_out[120]) );
  DFQD1 text_out_reg_95_ ( .D(N384), .CP(clk), .Q(text_out[95]) );
  DFQD1 text_out_reg_94_ ( .D(N385), .CP(clk), .Q(text_out[94]) );
  DFQD1 text_out_reg_93_ ( .D(N386), .CP(clk), .Q(text_out[93]) );
  DFQD1 text_out_reg_92_ ( .D(N387), .CP(clk), .Q(text_out[92]) );
  DFQD1 text_out_reg_91_ ( .D(N388), .CP(clk), .Q(text_out[91]) );
  DFQD1 text_out_reg_90_ ( .D(N389), .CP(clk), .Q(text_out[90]) );
  DFQD1 text_out_reg_89_ ( .D(N390), .CP(clk), .Q(text_out[89]) );
  DFQD1 text_out_reg_88_ ( .D(N391), .CP(clk), .Q(text_out[88]) );
  DFQD1 text_out_reg_63_ ( .D(N392), .CP(clk), .Q(text_out[63]) );
  DFQD1 text_out_reg_62_ ( .D(N393), .CP(clk), .Q(text_out[62]) );
  DFQD1 text_out_reg_61_ ( .D(N394), .CP(clk), .Q(text_out[61]) );
  DFQD1 text_out_reg_60_ ( .D(N395), .CP(clk), .Q(text_out[60]) );
  DFQD1 text_out_reg_59_ ( .D(N396), .CP(clk), .Q(text_out[59]) );
  DFQD1 text_out_reg_58_ ( .D(N397), .CP(clk), .Q(text_out[58]) );
  DFQD1 text_out_reg_57_ ( .D(N398), .CP(clk), .Q(text_out[57]) );
  DFQD1 text_out_reg_56_ ( .D(N399), .CP(clk), .Q(text_out[56]) );
  DFQD1 text_out_reg_31_ ( .D(N400), .CP(clk), .Q(text_out[31]) );
  DFQD1 text_out_reg_30_ ( .D(N401), .CP(clk), .Q(text_out[30]) );
  DFQD1 text_out_reg_29_ ( .D(N402), .CP(clk), .Q(text_out[29]) );
  DFQD1 text_out_reg_28_ ( .D(N403), .CP(clk), .Q(text_out[28]) );
  DFQD1 text_out_reg_27_ ( .D(N404), .CP(clk), .Q(text_out[27]) );
  DFQD1 text_out_reg_26_ ( .D(N405), .CP(clk), .Q(text_out[26]) );
  DFQD1 text_out_reg_25_ ( .D(N406), .CP(clk), .Q(text_out[25]) );
  DFQD1 text_out_reg_24_ ( .D(N407), .CP(clk), .Q(text_out[24]) );
  DFQD1 text_out_reg_119_ ( .D(N408), .CP(clk), .Q(text_out[119]) );
  DFQD1 text_out_reg_118_ ( .D(N409), .CP(clk), .Q(text_out[118]) );
  DFQD1 text_out_reg_117_ ( .D(N410), .CP(clk), .Q(text_out[117]) );
  DFQD1 text_out_reg_116_ ( .D(N411), .CP(clk), .Q(text_out[116]) );
  DFQD1 text_out_reg_115_ ( .D(N412), .CP(clk), .Q(text_out[115]) );
  DFQD1 text_out_reg_114_ ( .D(N413), .CP(clk), .Q(text_out[114]) );
  DFQD1 text_out_reg_113_ ( .D(N414), .CP(clk), .Q(text_out[113]) );
  DFQD1 text_out_reg_112_ ( .D(N415), .CP(clk), .Q(text_out[112]) );
  DFQD1 text_out_reg_87_ ( .D(N416), .CP(clk), .Q(text_out[87]) );
  DFQD1 text_out_reg_86_ ( .D(N417), .CP(clk), .Q(text_out[86]) );
  DFQD1 text_out_reg_85_ ( .D(N418), .CP(clk), .Q(text_out[85]) );
  DFQD1 text_out_reg_84_ ( .D(N419), .CP(clk), .Q(text_out[84]) );
  DFQD1 text_out_reg_83_ ( .D(N420), .CP(clk), .Q(text_out[83]) );
  DFQD1 text_out_reg_82_ ( .D(N421), .CP(clk), .Q(text_out[82]) );
  DFQD1 text_out_reg_81_ ( .D(N422), .CP(clk), .Q(text_out[81]) );
  DFQD1 text_out_reg_80_ ( .D(N423), .CP(clk), .Q(text_out[80]) );
  DFQD1 text_out_reg_55_ ( .D(N424), .CP(clk), .Q(text_out[55]) );
  DFQD1 text_out_reg_54_ ( .D(N425), .CP(clk), .Q(text_out[54]) );
  DFQD1 text_out_reg_53_ ( .D(N426), .CP(clk), .Q(text_out[53]) );
  DFQD1 text_out_reg_52_ ( .D(N427), .CP(clk), .Q(text_out[52]) );
  DFQD1 text_out_reg_51_ ( .D(N428), .CP(clk), .Q(text_out[51]) );
  DFQD1 text_out_reg_50_ ( .D(N429), .CP(clk), .Q(text_out[50]) );
  DFQD1 text_out_reg_49_ ( .D(N430), .CP(clk), .Q(text_out[49]) );
  DFQD1 text_out_reg_48_ ( .D(N431), .CP(clk), .Q(text_out[48]) );
  DFQD1 text_out_reg_23_ ( .D(N432), .CP(clk), .Q(text_out[23]) );
  DFQD1 text_out_reg_22_ ( .D(N433), .CP(clk), .Q(text_out[22]) );
  DFQD1 text_out_reg_21_ ( .D(N434), .CP(clk), .Q(text_out[21]) );
  DFQD1 text_out_reg_20_ ( .D(N435), .CP(clk), .Q(text_out[20]) );
  DFQD1 text_out_reg_19_ ( .D(N436), .CP(clk), .Q(text_out[19]) );
  DFQD1 text_out_reg_18_ ( .D(N437), .CP(clk), .Q(text_out[18]) );
  DFQD1 text_out_reg_17_ ( .D(N438), .CP(clk), .Q(text_out[17]) );
  DFQD1 text_out_reg_16_ ( .D(N439), .CP(clk), .Q(text_out[16]) );
  DFQD1 text_out_reg_111_ ( .D(N440), .CP(clk), .Q(text_out[111]) );
  DFQD1 text_out_reg_110_ ( .D(N441), .CP(clk), .Q(text_out[110]) );
  DFQD1 text_out_reg_109_ ( .D(N442), .CP(clk), .Q(text_out[109]) );
  DFQD1 text_out_reg_108_ ( .D(N443), .CP(clk), .Q(text_out[108]) );
  DFQD1 text_out_reg_107_ ( .D(N444), .CP(clk), .Q(text_out[107]) );
  DFQD1 text_out_reg_106_ ( .D(N445), .CP(clk), .Q(text_out[106]) );
  DFQD1 text_out_reg_105_ ( .D(N446), .CP(clk), .Q(text_out[105]) );
  DFQD1 text_out_reg_104_ ( .D(N447), .CP(clk), .Q(text_out[104]) );
  DFQD1 text_out_reg_79_ ( .D(N448), .CP(clk), .Q(text_out[79]) );
  DFQD1 text_out_reg_78_ ( .D(N449), .CP(clk), .Q(text_out[78]) );
  DFQD1 text_out_reg_77_ ( .D(N450), .CP(clk), .Q(text_out[77]) );
  DFQD1 text_out_reg_76_ ( .D(N451), .CP(clk), .Q(text_out[76]) );
  DFQD1 text_out_reg_75_ ( .D(N452), .CP(clk), .Q(text_out[75]) );
  DFQD1 text_out_reg_74_ ( .D(N453), .CP(clk), .Q(text_out[74]) );
  DFQD1 text_out_reg_73_ ( .D(N454), .CP(clk), .Q(text_out[73]) );
  DFQD1 text_out_reg_72_ ( .D(N455), .CP(clk), .Q(text_out[72]) );
  DFQD1 text_out_reg_47_ ( .D(N456), .CP(clk), .Q(text_out[47]) );
  DFQD1 text_out_reg_46_ ( .D(N457), .CP(clk), .Q(text_out[46]) );
  DFQD1 text_out_reg_45_ ( .D(N458), .CP(clk), .Q(text_out[45]) );
  DFQD1 text_out_reg_44_ ( .D(N459), .CP(clk), .Q(text_out[44]) );
  DFQD1 text_out_reg_43_ ( .D(N460), .CP(clk), .Q(text_out[43]) );
  DFQD1 text_out_reg_42_ ( .D(N461), .CP(clk), .Q(text_out[42]) );
  DFQD1 text_out_reg_41_ ( .D(N462), .CP(clk), .Q(text_out[41]) );
  DFQD1 text_out_reg_40_ ( .D(N463), .CP(clk), .Q(text_out[40]) );
  DFQD1 text_out_reg_15_ ( .D(N464), .CP(clk), .Q(text_out[15]) );
  DFQD1 text_out_reg_14_ ( .D(N465), .CP(clk), .Q(text_out[14]) );
  DFQD1 text_out_reg_13_ ( .D(N466), .CP(clk), .Q(text_out[13]) );
  DFQD1 text_out_reg_12_ ( .D(N467), .CP(clk), .Q(text_out[12]) );
  DFQD1 text_out_reg_11_ ( .D(N468), .CP(clk), .Q(text_out[11]) );
  DFQD1 text_out_reg_10_ ( .D(N469), .CP(clk), .Q(text_out[10]) );
  DFQD1 text_out_reg_9_ ( .D(N470), .CP(clk), .Q(text_out[9]) );
  DFQD1 text_out_reg_8_ ( .D(N471), .CP(clk), .Q(text_out[8]) );
  DFQD1 text_out_reg_103_ ( .D(N472), .CP(clk), .Q(text_out[103]) );
  DFQD1 text_out_reg_102_ ( .D(N473), .CP(clk), .Q(text_out[102]) );
  DFQD1 text_out_reg_101_ ( .D(N474), .CP(clk), .Q(text_out[101]) );
  DFQD1 text_out_reg_100_ ( .D(N475), .CP(clk), .Q(text_out[100]) );
  DFQD1 text_out_reg_99_ ( .D(N476), .CP(clk), .Q(text_out[99]) );
  DFQD1 text_out_reg_98_ ( .D(N477), .CP(clk), .Q(text_out[98]) );
  DFQD1 text_out_reg_97_ ( .D(N478), .CP(clk), .Q(text_out[97]) );
  DFQD1 text_out_reg_96_ ( .D(N479), .CP(clk), .Q(text_out[96]) );
  DFQD1 text_out_reg_71_ ( .D(N480), .CP(clk), .Q(text_out[71]) );
  DFQD1 text_out_reg_70_ ( .D(N481), .CP(clk), .Q(text_out[70]) );
  DFQD1 text_out_reg_69_ ( .D(N482), .CP(clk), .Q(text_out[69]) );
  DFQD1 text_out_reg_68_ ( .D(N483), .CP(clk), .Q(text_out[68]) );
  DFQD1 text_out_reg_67_ ( .D(N484), .CP(clk), .Q(text_out[67]) );
  DFQD1 text_out_reg_66_ ( .D(N485), .CP(clk), .Q(text_out[66]) );
  DFQD1 text_out_reg_65_ ( .D(N486), .CP(clk), .Q(text_out[65]) );
  DFQD1 text_out_reg_64_ ( .D(N487), .CP(clk), .Q(text_out[64]) );
  DFQD1 text_out_reg_39_ ( .D(N488), .CP(clk), .Q(text_out[39]) );
  DFQD1 text_out_reg_38_ ( .D(N489), .CP(clk), .Q(text_out[38]) );
  DFQD1 text_out_reg_37_ ( .D(N490), .CP(clk), .Q(text_out[37]) );
  DFQD1 text_out_reg_36_ ( .D(N491), .CP(clk), .Q(text_out[36]) );
  DFQD1 text_out_reg_35_ ( .D(N492), .CP(clk), .Q(text_out[35]) );
  DFQD1 text_out_reg_34_ ( .D(N493), .CP(clk), .Q(text_out[34]) );
  DFQD1 text_out_reg_33_ ( .D(N494), .CP(clk), .Q(text_out[33]) );
  DFQD1 text_out_reg_32_ ( .D(N495), .CP(clk), .Q(text_out[32]) );
  DFQD1 text_out_reg_7_ ( .D(N496), .CP(clk), .Q(text_out[7]) );
  DFQD1 text_out_reg_6_ ( .D(N497), .CP(clk), .Q(text_out[6]) );
  DFQD1 text_out_reg_5_ ( .D(N498), .CP(clk), .Q(text_out[5]) );
  DFQD1 text_out_reg_4_ ( .D(N499), .CP(clk), .Q(text_out[4]) );
  DFQD1 text_out_reg_3_ ( .D(N500), .CP(clk), .Q(text_out[3]) );
  DFQD1 text_out_reg_2_ ( .D(N501), .CP(clk), .Q(text_out[2]) );
  DFQD1 text_out_reg_1_ ( .D(N502), .CP(clk), .Q(text_out[1]) );
  DFQD1 text_out_reg_0_ ( .D(N503), .CP(clk), .Q(text_out[0]) );
  XNR2D1 U6 ( .A1(text_in_r[35]), .A2(w2[3]), .ZN(n95) );
  MOAI22D1 U7 ( .A1(n101), .A2(net7009), .B1(net7009), .B2(n102), .ZN(N98) );
  XNR2D1 U8 ( .A1(text_in_r[34]), .A2(w2[2]), .ZN(n101) );
  XNR2D1 U12 ( .A1(text_in_r[33]), .A2(w2[1]), .ZN(n105) );
  XNR2D1 U45 ( .A1(text_in_r[22]), .A2(w3[22]), .ZN(n147) );
  MOAI22D1 U62 ( .A1(n169), .A2(net7009), .B1(n170), .B2(net7009), .ZN(N64) );
  XNR2D1 U64 ( .A1(text_in_r[16]), .A2(w3[16]), .ZN(n169) );
  XNR2D1 U68 ( .A1(text_in_r[15]), .A2(w3[15]), .ZN(n172) );
  XNR2D1 U72 ( .A1(text_in_r[14]), .A2(w3[14]), .ZN(n175) );
  XNR2D1 U79 ( .A1(text_in_r[12]), .A2(w3[12]), .ZN(n181) );
  CKXOR2D1 U92 ( .A1(w3[5]), .A2(n584), .Z(N498) );
  CKXOR2D1 U93 ( .A1(w3[6]), .A2(sa33_sr[6]), .Z(N497) );
  CKXOR2D1 U95 ( .A1(w2[0]), .A2(n630), .Z(N495) );
  CKXOR2D1 U123 ( .A1(w0[6]), .A2(n601), .Z(N473) );
  CKXOR2D1 U131 ( .A1(w3[14]), .A2(sa23_sr[6]), .Z(N465) );
  CKXOR2D1 U132 ( .A1(w3[15]), .A2(n613), .Z(N464) );
  CKXOR2D1 U133 ( .A1(w2[8]), .A2(sa22_sr[0]), .Z(N463) );
  CKXOR2D1 U135 ( .A1(w2[10]), .A2(sa22_sr[2]), .Z(N461) );
  CKXOR2D1 U138 ( .A1(w2[13]), .A2(sa22_sr[5]), .Z(N458) );
  CKXOR2D1 U139 ( .A1(w2[14]), .A2(sa22_sr[6]), .Z(N457) );
  CKXOR2D1 U141 ( .A1(w1[8]), .A2(n548), .Z(N455) );
  CKXOR2D1 U143 ( .A1(w1[10]), .A2(sa21_sr[2]), .Z(N453) );
  CKXOR2D1 U147 ( .A1(w1[14]), .A2(n571), .Z(N449) );
  CKXOR2D1 U151 ( .A1(w0[10]), .A2(sa20_sr[2]), .Z(N445) );
  CKXOR2D1 U153 ( .A1(w0[12]), .A2(n624), .Z(N443) );
  CKXOR2D1 U154 ( .A1(w0[13]), .A2(sa20_sr[5]), .Z(N442) );
  CKXOR2D1 U155 ( .A1(w0[14]), .A2(sa20_sr[6]), .Z(N441) );
  CKXOR2D1 U163 ( .A1(w3[22]), .A2(sa13_sr[6]), .Z(N433) );
  CKXOR2D1 U170 ( .A1(w2[21]), .A2(sa12_sr[5]), .Z(N426) );
  CKXOR2D1 U173 ( .A1(w1[16]), .A2(sa11_sr[0]), .Z(N423) );
  CKXOR2D1 U175 ( .A1(w1[18]), .A2(n675), .Z(N421) );
  CKXOR2D1 U178 ( .A1(w1[21]), .A2(sa11_sr[5]), .Z(N418) );
  CKXOR2D1 U179 ( .A1(w1[22]), .A2(sa11_sr[6]), .Z(N417) );
  CKXOR2D1 U181 ( .A1(w0[16]), .A2(n574), .Z(N415) );
  CKXOR2D1 U183 ( .A1(w0[18]), .A2(sa10_sr[2]), .Z(N413) );
  CKXOR2D1 U186 ( .A1(w0[21]), .A2(sa10_sr[5]), .Z(N410) );
  CKXOR2D1 U194 ( .A1(w3[29]), .A2(sa03_sr[5]), .Z(N402) );
  CKXOR2D1 U195 ( .A1(w3[30]), .A2(sa03_sr[6]), .Z(N401) );
  CKXOR2D1 U197 ( .A1(w2[24]), .A2(n591), .Z(N399) );
  CKXOR2D1 U199 ( .A1(w2[26]), .A2(sa02_sr[2]), .Z(N397) );
  CKXOR2D1 U200 ( .A1(w2[27]), .A2(sa02_sr[3]), .Z(N396) );
  CKXOR2D1 U211 ( .A1(w1[26]), .A2(sa01_sr[2]), .Z(N389) );
  CKXOR2D1 U216 ( .A1(w1[31]), .A2(n566), .Z(N384) );
  CKXOR2D1 U219 ( .A1(w0[26]), .A2(n606), .Z(N381) );
  CKXOR2D1 U222 ( .A1(sa33_sr[5]), .A2(sa03_sr[5]), .Z(n152) );
  CKXOR2D1 U223 ( .A1(sa23_sr[6]), .A2(sa13_sr[6]), .Z(n119) );
  CKXOR2D1 U226 ( .A1(w0[29]), .A2(sa00_sr[5]), .Z(N378) );
  CKXOR2D1 U227 ( .A1(w0[30]), .A2(sa00_sr[6]), .Z(N377) );
  CKXOR2D1 U228 ( .A1(w0[31]), .A2(n554), .Z(N376) );
  CKXOR2D1 U230 ( .A1(sa03_sr[4]), .A2(sa33_sr[4]), .Z(n156) );
  CKXOR2D1 U231 ( .A1(sa23_sr[5]), .A2(sa13_sr[5]), .Z(n123) );
  CKXOR2D1 U243 ( .A1(sa03_sr[2]), .A2(sa33_sr[2]), .Z(n164) );
  CKXOR2D1 U244 ( .A1(text_in_r[3]), .A2(n712), .Z(n205) );
  CKXOR2D1 U247 ( .A1(sa23_sr[2]), .A2(sa13_sr[2]), .Z(n136) );
  CKXOR2D1 U257 ( .A1(sa23_sr[0]), .A2(n82), .Z(n144) );
  XNR2D1 U262 ( .A1(text_in_r[127]), .A2(w0[31]), .ZN(n215) );
  CKXOR2D1 U266 ( .A1(text_in_r[126]), .A2(n76), .Z(n219) );
  CKXOR2D1 U270 ( .A1(text_in_r[125]), .A2(n75), .Z(n223) );
  CKXOR2D1 U280 ( .A1(text_in_r[122]), .A2(n72), .Z(n236) );
  CKXOR2D1 U295 ( .A1(text_in_r[116]), .A2(n68), .Z(n255) );
  XNR2D1 U312 ( .A1(text_in_r[111]), .A2(w0[15]), .ZN(n274) );
  XNR2D1 U316 ( .A1(text_in_r[110]), .A2(w0[14]), .ZN(n277) );
  XNR2D1 U320 ( .A1(text_in_r[109]), .A2(w0[13]), .ZN(n280) );
  MOAI22D1 U324 ( .A1(n286), .A2(net7009), .B1(net7009), .B2(n287), .ZN(N243)
         );
  XNR2D1 U330 ( .A1(text_in_r[106]), .A2(w0[10]), .ZN(n289) );
  CKXOR2D1 U338 ( .A1(sa30_sr[6]), .A2(sa00_sr[6]), .Z(n251) );
  CKXOR2D1 U342 ( .A1(sa30_sr[5]), .A2(sa00_sr[5]), .Z(n254) );
  CKXOR2D1 U343 ( .A1(sa20_sr[6]), .A2(sa10_sr[6]), .Z(n221) );
  CKXOR2D1 U344 ( .A1(text_in_r[102]), .A2(n60), .Z(n299) );
  CKXOR2D1 U346 ( .A1(sa30_sr[4]), .A2(sa00_sr[4]), .Z(n258) );
  CKXOR2D1 U347 ( .A1(sa20_sr[5]), .A2(sa10_sr[5]), .Z(n225) );
  CKXOR2D1 U353 ( .A1(sa30_sr[3]), .A2(sa00_sr[3]), .Z(n262) );
  CKXOR2D1 U359 ( .A1(sa30_sr[2]), .A2(sa00_sr[2]), .Z(n266) );
  CKXOR2D1 U360 ( .A1(text_in_r[99]), .A2(n57), .Z(n307) );
  CKXOR2D1 U362 ( .A1(sa00_sr[1]), .A2(sa30_sr[1]), .Z(n269) );
  CKXOR2D1 U369 ( .A1(sa00_sr[0]), .A2(sa30_sr[0]), .Z(n273) );
  XNR2D1 U378 ( .A1(text_in_r[95]), .A2(w1[31]), .ZN(n317) );
  CKXOR2D1 U382 ( .A1(text_in_r[94]), .A2(n54), .Z(n321) );
  XNR2D1 U417 ( .A1(text_in_r[83]), .A2(w1[19]), .ZN(n363) );
  XNR2D1 U430 ( .A1(text_in_r[79]), .A2(w1[15]), .ZN(n377) );
  XNR2D1 U434 ( .A1(text_in_r[78]), .A2(w1[14]), .ZN(n380) );
  XNR2D1 U438 ( .A1(text_in_r[77]), .A2(w1[13]), .ZN(n383) );
  CKXOR2D1 U444 ( .A1(text_in_r[75]), .A2(n42), .Z(n389) );
  XNR2D1 U448 ( .A1(text_in_r[74]), .A2(w1[10]), .ZN(n392) );
  CKXOR2D1 U456 ( .A1(sa31_sr[6]), .A2(sa01_sr[6]), .Z(n354) );
  CKXOR2D1 U460 ( .A1(sa31_sr[5]), .A2(sa01_sr[5]), .Z(n357) );
  CKXOR2D1 U461 ( .A1(sa21_sr[6]), .A2(sa11_sr[6]), .Z(n323) );
  CKXOR2D1 U462 ( .A1(text_in_r[70]), .A2(n38), .Z(n402) );
  CKXOR2D1 U464 ( .A1(sa01_sr[4]), .A2(sa31_sr[4]), .Z(n361) );
  CKXOR2D1 U465 ( .A1(sa21_sr[5]), .A2(sa11_sr[5]), .Z(n327) );
  CKXOR2D1 U471 ( .A1(sa01_sr[3]), .A2(sa31_sr[3]), .Z(n365) );
  XNR2D1 U476 ( .A1(sa21_sr[3]), .A2(sa11_sr[3]), .ZN(n336) );
  CKXOR2D1 U477 ( .A1(sa31_sr[2]), .A2(sa01_sr[2]), .Z(n369) );
  CKXOR2D1 U482 ( .A1(text_in_r[66]), .A2(n34), .Z(n413) );
  CKXOR2D1 U487 ( .A1(sa01_sr[0]), .A2(sa31_sr[0]), .Z(n376) );
  XNR2D1 U497 ( .A1(text_in_r[63]), .A2(w2[31]), .ZN(n423) );
  XNR2D1 U501 ( .A1(text_in_r[62]), .A2(w2[30]), .ZN(n427) );
  CKXOR2D1 U507 ( .A1(text_in_r[61]), .A2(n32), .Z(n432) );
  CKXOR2D1 U510 ( .A1(text_in_r[60]), .A2(n31), .Z(n436) );
  XNR2D1 U517 ( .A1(text_in_r[58]), .A2(w2[26]), .ZN(n444) );
  CKXOR2D1 U526 ( .A1(text_in_r[55]), .A2(n27), .Z(n454) );
  CKXOR2D1 U535 ( .A1(text_in_r[52]), .A2(n24), .Z(n462) );
  XNR2D1 U539 ( .A1(sa22_sr[2]), .A2(sa12_sr[2]), .ZN(n104) );
  CKXOR2D1 U540 ( .A1(text_in_r[51]), .A2(n23), .Z(n467) );
  XNR2D1 U561 ( .A1(text_in_r[47]), .A2(w2[15]), .ZN(n478) );
  XNR2D1 U565 ( .A1(text_in_r[46]), .A2(w2[14]), .ZN(n481) );
  CKXOR2D1 U575 ( .A1(text_in_r[43]), .A2(n18), .Z(n490) );
  CKXOR2D1 U579 ( .A1(sa32_sr[2]), .A2(sa02_sr[2]), .Z(n100) );
  XNR2D1 U580 ( .A1(text_in_r[42]), .A2(w2[10]), .ZN(n493) );
  CKXOR2D1 U588 ( .A1(text_in_r[40]), .A2(n16), .Z(n499) );
  CKXOR2D1 U590 ( .A1(sa32_sr[6]), .A2(sa02_sr[6]), .Z(n458) );
  CKXOR2D1 U594 ( .A1(sa32_sr[5]), .A2(sa02_sr[5]), .Z(n461) );
  CKXOR2D1 U595 ( .A1(sa22_sr[6]), .A2(sa12_sr[6]), .Z(n429) );
  CKXOR2D1 U596 ( .A1(text_in_r[38]), .A2(n14), .Z(n503) );
  CKXOR2D1 U598 ( .A1(sa02_sr[4]), .A2(sa32_sr[4]), .Z(n465) );
  CKXOR2D1 U599 ( .A1(sa22_sr[5]), .A2(sa12_sr[5]), .Z(n434) );
  CKXOR2D1 U605 ( .A1(sa02_sr[3]), .A2(sa32_sr[3]), .Z(n469) );
  CKXOR2D1 U607 ( .A1(text_in_r[36]), .A2(n12), .Z(n507) );
  XOR4D0 U707 ( .A1(n127), .A2(n144), .A3(n526), .A4(w3[24]), .Z(n143) );
  XOR4D0 U715 ( .A1(n115), .A2(n167), .A3(sa13_sr[1]), .A4(n192), .Z(n191) );
  XOR4D0 U718 ( .A1(n119), .A2(n152), .A3(sa03_sr[6]), .A4(n10), .Z(n198) );
  XOR4D0 U719 ( .A1(n123), .A2(n9), .A3(sa03_sr[5]), .A4(n156), .Z(n200) );
  XOR4D0 U721 ( .A1(n144), .A2(n203), .A3(sa03_sr[0]), .A4(w3[0]), .Z(n214) );
  XOR4D0 U727 ( .A1(n225), .A2(n251), .A3(sa20_sr[6]), .A4(n69), .Z(n250) );
  XOR4D0 U728 ( .A1(n230), .A2(n254), .A3(sa20_sr[5]), .A4(w0[21]), .Z(n253)
         );
  XOR4D0 U729 ( .A1(n266), .A2(n242), .A3(sa20_sr[2]), .A4(w0[18]), .Z(n265)
         );
  XOR4D0 U733 ( .A1(n84), .A2(n269), .A3(n217), .A4(n294), .Z(n293) );
  XOR4D0 U737 ( .A1(n225), .A2(n258), .A3(sa00_sr[5]), .A4(n59), .Z(n302) );
  XOR4D0 U741 ( .A1(n544), .A2(n336), .A3(sa01_sr[2]), .A4(n337), .Z(n335) );
  XOR4D0 U750 ( .A1(n319), .A2(n365), .A3(n547), .A4(n391), .Z(n390) );
  XOR4D0 U754 ( .A1(n323), .A2(n357), .A3(sa01_sr[6]), .A4(n38), .Z(n403) );
  XOR4D0 U755 ( .A1(n327), .A2(sa01_sr[5]), .A3(n361), .A4(n37), .Z(n405) );
  XOR4D0 U768 ( .A1(n469), .A2(n425), .A3(sa12_sr[3]), .A4(n492), .Z(n491) );
  XOR4D0 U769 ( .A1(n103), .A2(n425), .A3(n639), .A4(n498), .Z(n497) );
  XOR4D0 U771 ( .A1(n438), .A2(n458), .A3(n573), .A4(n15), .Z(n502) );
  XOR4D0 U772 ( .A1(n429), .A2(n461), .A3(sa02_sr[6]), .A4(n14), .Z(n504) );
  DFQD4 sa12_reg_1_ ( .D(N129), .CP(clk), .Q(sa12[1]) );
  DFQD4 sa32_reg_1_ ( .D(N97), .CP(clk), .Q(sa32[1]) );
  DFQD4 sa21_reg_2_ ( .D(N178), .CP(clk), .Q(sa21[2]) );
  DFQD4 sa00_reg_2_ ( .D(N274), .CP(clk), .Q(sa00[2]) );
  DFQD4 sa11_reg_2_ ( .D(N194), .CP(clk), .Q(sa11[2]) );
  DFQD1 sa13_reg_0_ ( .D(N64), .CP(clk), .Q(sa13[0]) );
  DFQD1 sa13_reg_5_ ( .D(N69), .CP(clk), .Q(sa13[5]) );
  DFQD1 sa00_reg_5_ ( .D(N277), .CP(clk), .Q(sa00[5]) );
  DFQD1 sa20_reg_7_ ( .D(N247), .CP(clk), .Q(sa20[7]) );
  DFQD1 sa01_reg_7_ ( .D(N215), .CP(clk), .Q(sa01[7]) );
  DFQD1 sa23_reg_7_ ( .D(N55), .CP(clk), .Q(sa23[7]) );
  DFQD1 sa31_reg_7_ ( .D(N167), .CP(clk), .Q(sa31[7]) );
  DFQD1 sa12_reg_7_ ( .D(N135), .CP(clk), .Q(sa12[7]) );
  DFQD1 sa33_reg_7_ ( .D(N39), .CP(clk), .Q(sa33[7]) );
  DFQD1 sa02_reg_7_ ( .D(N151), .CP(clk), .Q(sa02[7]) );
  DFQD1 sa22_reg_4_ ( .D(N116), .CP(clk), .Q(sa22[4]) );
  DFQD1 sa23_reg_0_ ( .D(N48), .CP(clk), .Q(sa23[0]) );
  DFQD1 sa11_reg_0_ ( .D(N192), .CP(clk), .Q(sa11[0]) );
  DFQD1 sa02_reg_0_ ( .D(N144), .CP(clk), .Q(sa02[0]) );
  DFQD1 sa23_reg_5_ ( .D(N53), .CP(clk), .Q(sa23[5]) );
  DFQD1 sa22_reg_5_ ( .D(N117), .CP(clk), .Q(sa22[5]) );
  DFQD1 sa31_reg_2_ ( .D(N162), .CP(clk), .Q(sa31[2]) );
  DFQD1 sa30_reg_2_ ( .D(N226), .CP(clk), .Q(sa30[2]) );
  DFQD1 sa12_reg_3_ ( .D(N131), .CP(clk), .Q(sa12[3]) );
  DFQD1 sa11_reg_3_ ( .D(N195), .CP(clk), .Q(sa11[3]) );
  DFQD1 sa30_reg_3_ ( .D(N227), .CP(clk), .Q(sa30[3]) );
  DFQD1 sa00_reg_3_ ( .D(N275), .CP(clk), .Q(sa00[3]) );
  DFQD1 sa10_reg_3_ ( .D(N259), .CP(clk), .Q(sa10[3]) );
  DFQD1 sa01_reg_3_ ( .D(N211), .CP(clk), .Q(sa01[3]) );
  DFQD1 sa20_reg_1_ ( .D(N241), .CP(clk), .Q(sa20[1]) );
  DFQD1 sa30_reg_7_ ( .D(N231), .CP(clk), .Q(sa30[7]) );
  DFQD1 sa32_reg_7_ ( .D(N103), .CP(clk), .Q(sa32[7]) );
  DFQD1 sa01_reg_4_ ( .D(N212), .CP(clk), .Q(sa01[4]) );
  DFQD1 sa10_reg_5_ ( .D(N261), .CP(clk), .Q(sa10[5]) );
  DFQD1 sa23_reg_3_ ( .D(N51), .CP(clk), .Q(sa23[3]) );
  DFQD1 sa30_reg_1_ ( .D(N225), .CP(clk), .Q(sa30[1]) );
  DFQD1 sa30_reg_0_ ( .D(N224), .CP(clk), .Q(sa30[0]) );
  DFQD1 sa01_reg_6_ ( .D(N214), .CP(clk), .Q(sa01[6]) );
  DFQD1 sa32_reg_2_ ( .D(N98), .CP(clk), .Q(sa32[2]) );
  DFQD1 sa02_reg_2_ ( .D(N146), .CP(clk), .Q(sa02[2]) );
  DFQD1 sa20_reg_2_ ( .D(N242), .CP(clk), .Q(sa20[2]) );
  DFQD1 sa01_reg_5_ ( .D(N213), .CP(clk), .Q(sa01[5]) );
  DFQD1 sa00_reg_0_ ( .D(N272), .CP(clk), .Q(sa00[0]) );
  DFQD1 sa22_reg_0_ ( .D(N112), .CP(clk), .Q(sa22[0]) );
  DFQD1 sa22_reg_2_ ( .D(N114), .CP(clk), .Q(sa22[2]) );
  DFQD1 sa32_reg_3_ ( .D(N99), .CP(clk), .Q(sa32[3]) );
  DFQD1 sa03_reg_1_ ( .D(N81), .CP(clk), .Q(sa03[1]) );
  DFQD1 sa00_reg_1_ ( .D(N273), .CP(clk), .Q(sa00[1]) );
  DFQD1 sa12_reg_6_ ( .D(N134), .CP(clk), .Q(sa12[6]) );
  DFQD1 sa33_reg_1_ ( .D(N33), .CP(clk), .Q(sa33[1]) );
  DFQD1 sa20_reg_6_ ( .D(N246), .CP(clk), .Q(sa20[6]) );
  DFQD1 sa23_reg_6_ ( .D(N54), .CP(clk), .Q(sa23[6]) );
  DFQD1 sa13_reg_2_ ( .D(N66), .CP(clk), .Q(sa13[2]) );
  DFQD1 sa12_reg_2_ ( .D(N130), .CP(clk), .Q(sa12[2]) );
  DFQD1 sa31_reg_0_ ( .D(N160), .CP(clk), .Q(sa31[0]) );
  DFQD4 sa02_reg_1_ ( .D(N145), .CP(clk), .Q(sa02[1]) );
  DFQD4 sa10_reg_0_ ( .D(N256), .CP(clk), .Q(sa10[0]) );
  DFQD4 sa03_reg_2_ ( .D(N82), .CP(clk), .Q(sa03[2]) );
  DFQD1 sa10_reg_2_ ( .D(N258), .CP(clk), .Q(sa10[2]) );
  DFQD4 sa02_reg_5_ ( .D(N149), .CP(clk), .Q(sa02[5]) );
  DFQD2 sa13_reg_6_ ( .D(N70), .CP(clk), .Q(sa13[6]) );
  CKXOR2D1 U208 ( .A1(sa33_sr[6]), .A2(sa03_sr[6]), .Z(n149) );
  DFQD1 sa33_reg_5_ ( .D(N37), .CP(clk), .Q(sa33[5]) );
  DFQD2 sa21_reg_1_ ( .D(N177), .CP(clk), .Q(sa21[1]) );
  DFQD1 sa11_reg_6_ ( .D(N198), .CP(clk), .Q(sa11[6]) );
  DFQD1 sa33_reg_2_ ( .D(N34), .CP(clk), .Q(sa33[2]) );
  DFQD1 sa10_reg_1_ ( .D(N257), .CP(clk), .Q(sa10[1]) );
  DFQD1 sa11_reg_7_ ( .D(N199), .CP(clk), .Q(sa11[7]) );
  DFQD1 sa31_reg_4_ ( .D(N164), .CP(clk), .Q(sa31[4]) );
  DFQD4 sa33_reg_0_ ( .D(N32), .CP(clk), .Q(sa33[0]) );
  DFQD1 sa10_reg_6_ ( .D(N262), .CP(clk), .Q(sa10[6]) );
  DFQD1 sa31_reg_5_ ( .D(N165), .CP(clk), .Q(sa31[5]) );
  DFQD1 sa31_reg_1_ ( .D(N161), .CP(clk), .Q(sa31[1]) );
  DFQD1 sa11_reg_1_ ( .D(N193), .CP(clk), .Q(sa11[1]) );
  DFQD2 sa31_reg_6_ ( .D(N166), .CP(clk), .Q(sa31[6]) );
  DFQD1 sa01_reg_1_ ( .D(N209), .CP(clk), .Q(sa01[1]) );
  DFQD2 sa33_reg_6_ ( .D(N38), .CP(clk), .Q(sa33[6]) );
  DFQD4 sa03_reg_3_ ( .D(N83), .CP(clk), .Q(sa03[3]) );
  DFQD2 sa32_reg_5_ ( .D(N101), .CP(clk), .Q(sa32[5]) );
  DFQD1 sa02_reg_3_ ( .D(N147), .CP(clk), .Q(sa02[3]) );
  DFQD1 sa11_reg_4_ ( .D(N196), .CP(clk), .Q(sa11[4]) );
  DFQD2 sa21_reg_6_ ( .D(N182), .CP(clk), .Q(sa21[6]) );
  DFQD4 sa33_reg_3_ ( .D(N35), .CP(clk), .Q(sa33[3]) );
  DFQD1 sa30_reg_5_ ( .D(N229), .CP(clk), .Q(sa30[5]) );
  DFQD1 sa22_reg_1_ ( .D(N113), .CP(clk), .Q(sa22[1]) );
  DFQD1 sa03_reg_0_ ( .D(N80), .CP(clk), .Q(sa03[0]) );
  DFQD1 sa22_reg_6_ ( .D(N118), .CP(clk), .Q(sa22[6]) );
  DFQD1 sa20_reg_3_ ( .D(N243), .CP(clk), .Q(sa20[3]) );
  DFQD1 sa11_reg_5_ ( .D(N197), .CP(clk), .Q(sa11[5]) );
  DFQD1 sa21_reg_0_ ( .D(N176), .CP(clk), .Q(sa21[0]) );
  DFQD1 sa02_reg_6_ ( .D(N150), .CP(clk), .Q(sa02[6]) );
  DFQD1 sa03_reg_6_ ( .D(N86), .CP(clk), .Q(sa03[6]) );
  DFQD1 sa23_reg_4_ ( .D(N52), .CP(clk), .Q(sa23[4]) );
  DFQD1 sa12_reg_4_ ( .D(N132), .CP(clk), .Q(sa12[4]) );
  DFQD1 sa00_reg_4_ ( .D(N276), .CP(clk), .Q(sa00[4]) );
  DFQD2 sa01_reg_2_ ( .D(N210), .CP(clk), .Q(sa01[2]) );
  DFQD1 sa00_reg_6_ ( .D(N278), .CP(clk), .Q(sa00[6]) );
  DFQD1 sa01_reg_0_ ( .D(N208), .CP(clk), .Q(sa01[0]) );
  DFQD2 sa32_reg_6_ ( .D(N102), .CP(clk), .Q(sa32[6]) );
  DFQD2 sa22_reg_3_ ( .D(N115), .CP(clk), .Q(sa22[3]) );
  DFQD2 sa21_reg_3_ ( .D(N179), .CP(clk), .Q(sa21[3]) );
  DFQD2 sa23_reg_1_ ( .D(N49), .CP(clk), .Q(sa23[1]) );
  DFQD1 sa33_reg_4_ ( .D(N36), .CP(clk), .Q(sa33[4]) );
  DFQD2 sa10_reg_7_ ( .D(N263), .CP(clk), .Q(sa10[7]) );
  DFQD2 sa02_reg_4_ ( .D(N148), .CP(clk), .Q(sa02[4]) );
  INVD1 U774 ( .I(sa13_sr[4]), .ZN(n567) );
  XOR4D2 U775 ( .A1(n123), .A2(n149), .A3(sa23_sr[6]), .A4(w3[22]), .Z(n148)
         );
  CKXOR2D0 U776 ( .A1(w1[30]), .A2(sa01_sr[6]), .Z(N385) );
  XNR3D4 U777 ( .A1(n464), .A2(n465), .A3(n466), .ZN(n638) );
  XOR3D2 U778 ( .A1(n439), .A2(n469), .A3(n509), .Z(n508) );
  INVD0 U779 ( .I(sa10_sr[1]), .ZN(n84) );
  XOR4D2 U780 ( .A1(n434), .A2(n465), .A3(sa02_sr[5]), .A4(n13), .Z(n506) );
  XOR4D0 U781 ( .A1(n425), .A2(n465), .A3(n90), .A4(n489), .Z(n488) );
  MOAI22D1 U782 ( .A1(n316), .A2(net7021), .B1(n510), .B2(net7013), .ZN(N224)
         );
  XOR2D2 U783 ( .A1(text_in_r[96]), .A2(w0[0]), .Z(n510) );
  MOAI22D1 U784 ( .A1(n512), .A2(n511), .B1(n513), .B2(net7007), .ZN(N228) );
  INVD16 U785 ( .I(net7013), .ZN(n511) );
  XOR2D2 U786 ( .A1(text_in_r[100]), .A2(n58), .Z(n512) );
  XNR3D1 U787 ( .A1(n262), .A2(n305), .A3(n306), .ZN(n513) );
  CKND0 U788 ( .I(sa32_sr[1]), .ZN(n514) );
  INVD1 U789 ( .I(n514), .ZN(n515) );
  XOR3D1 U790 ( .A1(sa33_sr[4]), .A2(w3[13]), .A3(n92), .Z(n180) );
  MOAI22D2 U791 ( .A1(n436), .A2(net7009), .B1(n437), .B2(net7009), .ZN(N148)
         );
  XOR3D1 U792 ( .A1(n622), .A2(n225), .A3(n226), .Z(n224) );
  XOR3D1 U793 ( .A1(w0[31]), .A2(sa10_sr[7]), .A3(sa10_sr[6]), .Z(n659) );
  XOR4D2 U794 ( .A1(n408), .A2(n349), .A3(n635), .A4(w1[0]), .Z(n419) );
  MOAI22D1 U795 ( .A1(net7017), .A2(n485), .B1(n516), .B2(net7023), .ZN(N117)
         );
  XOR2D2 U796 ( .A1(text_in_r[45]), .A2(w2[13]), .Z(n516) );
  XOR4D2 U797 ( .A1(n559), .A2(n369), .A3(sa21_sr[2]), .A4(w1[18]), .Z(n368)
         );
  OAI22D2 U798 ( .A1(n450), .A2(net7005), .B1(net7017), .B2(n451), .ZN(N144)
         );
  XNR3D0 U799 ( .A1(w1[14]), .A2(sa31_sr[5]), .A3(sa21_sr[5]), .ZN(n382) );
  INVD1 U800 ( .I(sa03_sr[4]), .ZN(n557) );
  XOR4D0 U801 ( .A1(n522), .A2(n152), .A3(sa23_sr[5]), .A4(w3[21]), .Z(n151)
         );
  MOAI22D1 U802 ( .A1(net7025), .A2(n151), .B1(n517), .B2(net7017), .ZN(N69)
         );
  INVD16 U803 ( .I(n150), .ZN(n517) );
  XOR3D1 U804 ( .A1(n558), .A2(n123), .A3(n124), .Z(n122) );
  XOR4D0 U805 ( .A1(n115), .A2(n119), .A3(n81), .A4(w3[23]), .Z(n146) );
  MOAI22D1 U806 ( .A1(n502), .A2(net7017), .B1(n518), .B2(net7011), .ZN(N103)
         );
  XNR2D1 U807 ( .A1(text_in_r[39]), .A2(n15), .ZN(n518) );
  CKXOR2D0 U808 ( .A1(w3[11]), .A2(sa23_sr[3]), .Z(N468) );
  XOR3D4 U809 ( .A1(w3[19]), .A2(sa23_sr[3]), .A3(n136), .Z(n664) );
  XOR3D2 U810 ( .A1(w3[12]), .A2(sa23_sr[3]), .A3(n570), .Z(n183) );
  XOR2D4 U811 ( .A1(sa23_sr[7]), .A2(sa33_sr[7]), .Z(n115) );
  MOAI22D1 U812 ( .A1(net7025), .A2(n146), .B1(n519), .B2(net7023), .ZN(N71)
         );
  XOR2D2 U813 ( .A1(text_in_r[23]), .A2(w3[23]), .Z(n519) );
  MOAI22D2 U814 ( .A1(n147), .A2(net7009), .B1(net7009), .B2(n148), .ZN(N70)
         );
  CKBD1 U815 ( .I(sa30_sr[0]), .Z(n520) );
  MOAI22D1 U816 ( .A1(n272), .A2(net7023), .B1(n521), .B2(net7015), .ZN(N256)
         );
  XNR2D1 U817 ( .A1(text_in_r[112]), .A2(n66), .ZN(n521) );
  XOR3D2 U818 ( .A1(sa03_sr[3]), .A2(n711), .A3(n132), .Z(n207) );
  XOR2D0 U819 ( .A1(w3[27]), .A2(sa03_sr[3]), .Z(N404) );
  CKXOR2D1 U820 ( .A1(sa33_sr[3]), .A2(sa03_sr[3]), .Z(n160) );
  XOR4D0 U821 ( .A1(n629), .A2(n112), .A3(n591), .A4(w2[0]), .Z(n111) );
  CKXOR2D0 U822 ( .A1(w2[6]), .A2(sa32_sr[6]), .Z(N489) );
  XOR2D2 U823 ( .A1(sa22_sr[0]), .A2(sa12_sr[0]), .Z(n112) );
  OAI22D2 U824 ( .A1(n307), .A2(net6999), .B1(net7021), .B2(n308), .ZN(N227)
         );
  XOR3D2 U825 ( .A1(n266), .A2(n305), .A3(n309), .Z(n308) );
  CKXOR2D1 U826 ( .A1(n545), .A2(sa33_sr[1]), .Z(n683) );
  INVD1 U827 ( .I(n656), .ZN(n545) );
  XNR2D1 U828 ( .A1(sa23_sr[4]), .A2(sa13_sr[4]), .ZN(n522) );
  XNR2D1 U829 ( .A1(sa23_sr[4]), .A2(sa13_sr[4]), .ZN(n128) );
  XOR3D1 U830 ( .A1(w3[20]), .A2(sa23_sr[4]), .A3(n132), .Z(n157) );
  CKXOR2D0 U831 ( .A1(w0[5]), .A2(sa30_sr[5]), .Z(N474) );
  XOR3D4 U832 ( .A1(w1[1]), .A2(sa01_sr[1]), .A3(n345), .Z(n417) );
  CKND0 U833 ( .I(sa21_sr[1]), .ZN(n523) );
  INVD1 U834 ( .I(n523), .ZN(n524) );
  MOAI22D2 U835 ( .A1(n190), .A2(net7009), .B1(n191), .B2(net7009), .ZN(N49)
         );
  CKND0 U836 ( .I(sa33_sr[0]), .ZN(n525) );
  INVD1 U837 ( .I(n525), .ZN(n526) );
  XOR3D2 U838 ( .A1(w0[28]), .A2(sa10_sr[3]), .A3(sa30_sr[4]), .Z(n231) );
  XOR3D2 U839 ( .A1(sa21_sr[1]), .A2(w1[17]), .A3(n349), .Z(n373) );
  MOAI22D1 U840 ( .A1(net7017), .A2(n477), .B1(n527), .B2(net7011), .ZN(N128)
         );
  XNR2D1 U841 ( .A1(text_in_r[48]), .A2(n20), .ZN(n527) );
  MOAI22D1 U842 ( .A1(net7021), .A2(n302), .B1(n528), .B2(net7013), .ZN(N229)
         );
  XNR2D1 U843 ( .A1(text_in_r[101]), .A2(n59), .ZN(n528) );
  OAI22D2 U844 ( .A1(n474), .A2(net7017), .B1(n611), .B2(net7007), .ZN(N129)
         );
  CKND0 U845 ( .I(sa31_sr[0]), .ZN(n529) );
  INVD1 U846 ( .I(n529), .ZN(n530) );
  CKND0 U847 ( .I(w3[1]), .ZN(n710) );
  CKXOR2D0 U848 ( .A1(w3[1]), .A2(sa33_sr[1]), .Z(N502) );
  XOR3D2 U849 ( .A1(w3[1]), .A2(n545), .A3(n140), .Z(n212) );
  OAI22D2 U850 ( .A1(n299), .A2(net6999), .B1(net7021), .B2(n300), .ZN(N230)
         );
  MOAI22D2 U851 ( .A1(n389), .A2(net7009), .B1(net7009), .B2(n390), .ZN(N179)
         );
  XOR3D4 U852 ( .A1(n376), .A2(n408), .A3(n417), .Z(n416) );
  XOR3D4 U853 ( .A1(n360), .A2(n372), .A3(n373), .Z(n371) );
  OAI22D2 U854 ( .A1(n134), .A2(net6991), .B1(net7025), .B2(n135), .ZN(N82) );
  XNR3D1 U855 ( .A1(n545), .A2(n136), .A3(n665), .ZN(n135) );
  MOAI22D2 U856 ( .A1(n181), .A2(net7009), .B1(n182), .B2(net7009), .ZN(N52)
         );
  MOAI22D2 U857 ( .A1(n490), .A2(net7009), .B1(net7009), .B2(n491), .ZN(N115)
         );
  CKND0 U858 ( .I(sa33_sr[4]), .ZN(n531) );
  INVD1 U859 ( .I(n531), .ZN(n532) );
  CKND0 U860 ( .I(sa12_sr[0]), .ZN(n533) );
  INVD1 U861 ( .I(n533), .ZN(n534) );
  CKND0 U862 ( .I(sa21_sr[3]), .ZN(n535) );
  INVD1 U863 ( .I(n535), .ZN(n536) );
  XOR2D2 U864 ( .A1(sa10_sr[7]), .A2(sa00_sr[7]), .Z(n229) );
  XOR2D2 U865 ( .A1(sa20_sr[7]), .A2(sa10_sr[7]), .Z(n257) );
  XNR2D2 U866 ( .A1(sa02_sr[1]), .A2(sa32_sr[1]), .ZN(n103) );
  XOR3D1 U867 ( .A1(w2[29]), .A2(sa32_sr[5]), .A3(n90), .Z(n435) );
  CKXOR2D1 U868 ( .A1(sa31_sr[1]), .A2(sa01_sr[1]), .Z(n372) );
  CKXOR2D1 U869 ( .A1(sa03_sr[0]), .A2(sa33_sr[0]), .Z(n171) );
  CKXOR2D1 U870 ( .A1(sa32_sr[7]), .A2(sa22_sr[7]), .Z(n425) );
  CKXOR2D1 U871 ( .A1(sa30_sr[7]), .A2(sa00_sr[7]), .Z(n305) );
  CKBD1 U872 ( .I(sa10_sr[0]), .Z(n574) );
  INVD1 U873 ( .I(sa20_sr[3]), .ZN(n676) );
  XNR3D0 U874 ( .A1(w1[30]), .A2(sa31_sr[6]), .A3(sa11_sr[5]), .ZN(n324) );
  INVD1 U875 ( .I(w2[1]), .ZN(n546) );
  CKBD1 U876 ( .I(sa11_sr[2]), .Z(n675) );
  CKXOR2D1 U877 ( .A1(text_in_r[88]), .A2(w1[24]), .Z(n588) );
  CKXOR2D1 U878 ( .A1(text_in_r[84]), .A2(w1[20]), .Z(n556) );
  XOR3D1 U879 ( .A1(w1[26]), .A2(sa31_sr[2]), .A3(n87), .Z(n341) );
  CKXOR2D1 U880 ( .A1(text_in_r[0]), .A2(w3[0]), .Z(n640) );
  MOAI22D1 U881 ( .A1(n462), .A2(net7005), .B1(n637), .B2(n638), .ZN(N132) );
  INVD1 U882 ( .I(net7017), .ZN(n637) );
  CKXOR2D1 U883 ( .A1(text_in_r[68]), .A2(w1[4]), .Z(n620) );
  XOR4D0 U884 ( .A1(n319), .A2(n323), .A3(n78), .A4(w1[23]), .Z(n351) );
  XOR3D1 U885 ( .A1(n434), .A2(n564), .A3(n435), .Z(n433) );
  CKXOR2D1 U886 ( .A1(text_in_r[114]), .A2(w0[18]), .Z(n645) );
  XOR3D1 U887 ( .A1(w2[30]), .A2(sa32_sr[6]), .A3(sa12_sr[5]), .Z(n662) );
  CKXOR2D1 U888 ( .A1(text_in_r[18]), .A2(w3[18]), .Z(n631) );
  CKXOR2D1 U889 ( .A1(text_in_r[121]), .A2(w0[25]), .Z(n653) );
  CKXOR2D1 U890 ( .A1(text_in_r[25]), .A2(w3[25]), .Z(n655) );
  CKXOR2D1 U891 ( .A1(text_in_r[120]), .A2(w0[24]), .Z(n647) );
  OAI22D1 U892 ( .A1(n325), .A2(net7001), .B1(net7021), .B2(n326), .ZN(N213)
         );
  XOR3D1 U893 ( .A1(n626), .A2(n327), .A3(n328), .Z(n326) );
  CKXOR2D1 U894 ( .A1(text_in_r[97]), .A2(n55), .Z(n541) );
  CKXOR2D1 U895 ( .A1(text_in_r[105]), .A2(w0[9]), .Z(n654) );
  CKXOR2D1 U896 ( .A1(text_in_r[8]), .A2(w3[8]), .Z(n644) );
  XOR4D0 U897 ( .A1(n127), .A2(n149), .A3(n613), .A4(n11), .Z(n196) );
  XNR3D0 U898 ( .A1(w0[15]), .A2(sa30_sr[7]), .A3(n601), .ZN(n276) );
  XOR3D1 U899 ( .A1(w0[11]), .A2(sa30_sr[2]), .A3(sa20_sr[2]), .Z(n288) );
  XOR3D1 U900 ( .A1(w2[14]), .A2(sa32_sr[5]), .A3(sa22_sr[5]), .Z(n669) );
  CKXOR2D1 U901 ( .A1(text_in_r[82]), .A2(w1[18]), .Z(n561) );
  OAI22D1 U902 ( .A1(n236), .A2(net6995), .B1(net7023), .B2(n237), .ZN(N274)
         );
  XOR3D1 U903 ( .A1(n651), .A2(n238), .A3(n239), .Z(n237) );
  CKXOR2D1 U904 ( .A1(text_in_r[49]), .A2(n21), .Z(n611) );
  CKXOR2D1 U905 ( .A1(text_in_r[108]), .A2(w0[12]), .Z(n603) );
  XOR3D1 U906 ( .A1(n369), .A2(n408), .A3(n412), .Z(n411) );
  CKXOR2D1 U907 ( .A1(text_in_r[32]), .A2(w2[0]), .Z(n652) );
  CKXOR2D1 U908 ( .A1(text_in_r[19]), .A2(w3[19]), .Z(n594) );
  XOR3D1 U909 ( .A1(w3[10]), .A2(sa33_sr[1]), .A3(n91), .Z(n189) );
  CKXOR2D1 U910 ( .A1(text_in_r[17]), .A2(w3[17]), .Z(n604) );
  OAI22D1 U911 ( .A1(n377), .A2(net7003), .B1(net7019), .B2(n378), .ZN(N183)
         );
  OAI22D1 U912 ( .A1(n507), .A2(net6991), .B1(net7011), .B2(n508), .ZN(N100)
         );
  XOR4D1 U913 ( .A1(sa22_sr[5]), .A2(n461), .A3(n439), .A4(n25), .Z(n460) );
  XOR4D1 U914 ( .A1(n691), .A2(sa02_sr[3]), .A3(n439), .A4(n440), .Z(n437) );
  XOR3D1 U915 ( .A1(sa01_sr[1]), .A2(n340), .A3(n341), .Z(n339) );
  CKXOR2D1 U916 ( .A1(sa11_sr[2]), .A2(sa21_sr[2]), .Z(n340) );
  XOR4D0 U917 ( .A1(n238), .A2(n269), .A3(n606), .A4(n56), .Z(n311) );
  CKND0 U918 ( .I(sa31_sr[3]), .ZN(n537) );
  INVD1 U919 ( .I(n537), .ZN(n538) );
  XOR4D0 U920 ( .A1(n115), .A2(n171), .A3(n82), .A4(w3[8]), .Z(n194) );
  XOR3D1 U921 ( .A1(sa03_sr[6]), .A2(n115), .A3(n116), .Z(n114) );
  MOAI22D1 U922 ( .A1(n289), .A2(net6997), .B1(net7005), .B2(n539), .ZN(N242)
         );
  XNR3D0 U923 ( .A1(sa10_sr[2]), .A2(n266), .A3(n291), .ZN(n539) );
  INVD1 U924 ( .I(n92), .ZN(n540) );
  XOR4D1 U925 ( .A1(n127), .A2(n522), .A3(sa03_sr[3]), .A4(n129), .Z(n126) );
  XOR3D4 U926 ( .A1(w0[3]), .A2(sa00_sr[3]), .A3(n234), .Z(n309) );
  OAI22D2 U927 ( .A1(net7025), .A2(n615), .B1(n541), .B2(net6993), .ZN(N225)
         );
  XOR4D1 U928 ( .A1(n229), .A2(n579), .A3(n242), .A4(n243), .Z(n241) );
  CKND0 U929 ( .I(sa23_sr[4]), .ZN(n92) );
  CKXOR2D0 U930 ( .A1(w3[13]), .A2(sa23_sr[5]), .Z(N466) );
  XNR3D0 U931 ( .A1(w1[13]), .A2(sa31_sr[4]), .A3(sa21_sr[4]), .ZN(n385) );
  XOR4D1 U932 ( .A1(n229), .A2(n234), .A3(n606), .A4(n235), .Z(n233) );
  XOR4D1 U933 ( .A1(n217), .A2(n258), .A3(n681), .A4(n285), .Z(n284) );
  CKXOR2D1 U934 ( .A1(text_in_r[11]), .A2(w3[11]), .Z(n542) );
  CKBD0 U935 ( .I(sa12_sr[2]), .Z(n543) );
  CKXOR2D1 U936 ( .A1(sa11_sr[7]), .A2(sa01_sr[7]), .Z(n544) );
  CKXOR2D1 U937 ( .A1(sa11_sr[7]), .A2(sa01_sr[7]), .Z(n331) );
  XOR3D1 U938 ( .A1(n571), .A2(n544), .A3(n379), .Z(n378) );
  XOR4D0 U939 ( .A1(n229), .A2(n251), .A3(sa20_sr[7]), .A4(n61), .Z(n298) );
  XOR4D0 U940 ( .A1(n217), .A2(n273), .A3(n574), .A4(n62), .Z(n296) );
  CKXOR2D1 U941 ( .A1(sa31_sr[7]), .A2(sa01_sr[7]), .Z(n408) );
  INVD1 U942 ( .I(n656), .ZN(n657) );
  CKXOR2D0 U943 ( .A1(w3[18]), .A2(sa13_sr[2]), .Z(N437) );
  XOR3D1 U944 ( .A1(sa32_sr[1]), .A2(w2[10]), .A3(n614), .Z(n667) );
  CKXOR2D0 U945 ( .A1(w2[18]), .A2(n543), .Z(N429) );
  XOR3D4 U946 ( .A1(n257), .A2(n269), .A3(n270), .Z(n268) );
  XOR3D2 U947 ( .A1(sa02_sr[1]), .A2(n546), .A3(n98), .Z(n670) );
  CKBD0 U948 ( .I(sa11_sr[3]), .Z(n547) );
  CKBD0 U949 ( .I(sa21_sr[0]), .Z(n548) );
  XNR2D1 U950 ( .A1(sa21_sr[0]), .A2(sa11_sr[0]), .ZN(n349) );
  CKBD1 U951 ( .I(sa32_sr[3]), .Z(n549) );
  CKND0 U952 ( .I(n361), .ZN(n550) );
  INVD1 U953 ( .I(n550), .ZN(n551) );
  MOAI22D1 U954 ( .A1(net7021), .A2(n298), .B1(n552), .B2(net7013), .ZN(N231)
         );
  XNR2D1 U955 ( .A1(text_in_r[103]), .A2(n61), .ZN(n552) );
  CKND0 U956 ( .I(sa00_sr[7]), .ZN(n553) );
  INVD1 U957 ( .I(n553), .ZN(n554) );
  XOR3D1 U958 ( .A1(w0[26]), .A2(sa30_sr[2]), .A3(n84), .Z(n239) );
  MOAI22D1 U959 ( .A1(n555), .A2(net7023), .B1(n556), .B2(net7023), .ZN(N196)
         );
  XOR3D1 U960 ( .A1(n551), .A2(n360), .A3(n362), .Z(n555) );
  INVD1 U961 ( .I(n557), .ZN(n558) );
  CKXOR2D0 U962 ( .A1(w2[29]), .A2(sa02_sr[5]), .Z(N394) );
  XNR2D1 U963 ( .A1(sa21_sr[1]), .A2(sa11_sr[1]), .ZN(n559) );
  XNR2D1 U964 ( .A1(sa21_sr[1]), .A2(sa11_sr[1]), .ZN(n345) );
  XOR4D0 U965 ( .A1(n160), .A2(n115), .A3(n616), .A4(n186), .Z(n185) );
  CKXOR2D1 U966 ( .A1(sa12_sr[7]), .A2(sa22_sr[7]), .Z(n464) );
  CKBD0 U967 ( .I(sa03_sr[2]), .Z(n560) );
  XOR3D1 U968 ( .A1(w0[27]), .A2(sa30_sr[3]), .A3(sa10_sr[2]), .Z(n235) );
  XOR2D4 U969 ( .A1(sa20_sr[2]), .A2(sa10_sr[2]), .Z(n238) );
  XOR3D1 U970 ( .A1(w2[9]), .A2(sa32_sr[0]), .A3(sa22_sr[0]), .Z(n498) );
  INVD1 U971 ( .I(sa32_sr[0]), .ZN(n93) );
  MOAI22D1 U972 ( .A1(n368), .A2(net7019), .B1(n561), .B2(net7019), .ZN(N194)
         );
  XNR3D4 U973 ( .A1(w1[4]), .A2(n625), .A3(n332), .ZN(n409) );
  XOR4D0 U974 ( .A1(n217), .A2(n221), .A3(n553), .A4(w0[23]), .Z(n248) );
  XOR4D2 U975 ( .A1(n434), .A2(n458), .A3(sa22_sr[6]), .A4(n26), .Z(n457) );
  XOR4D0 U976 ( .A1(n88), .A2(n361), .A3(n319), .A4(n388), .Z(n387) );
  CKND0 U977 ( .I(sa10_sr[3]), .ZN(n677) );
  OAI22D2 U978 ( .A1(n499), .A2(net7009), .B1(n500), .B2(net7017), .ZN(N112)
         );
  XOR3D1 U979 ( .A1(sa13_sr[0]), .A2(w3[25]), .A3(sa33_sr[1]), .Z(n141) );
  MOAI22D1 U980 ( .A1(net7023), .A2(n250), .B1(n562), .B2(net7025), .ZN(N262)
         );
  XNR2D1 U981 ( .A1(text_in_r[118]), .A2(n69), .ZN(n562) );
  XOR3D1 U982 ( .A1(sa13_sr[2]), .A2(n164), .A3(n189), .Z(n188) );
  XOR3D4 U983 ( .A1(w1[19]), .A2(sa21_sr[3]), .A3(n340), .Z(n660) );
  XNR3D0 U984 ( .A1(w3[15]), .A2(sa33_sr[7]), .A3(sa33_sr[6]), .ZN(n174) );
  CKXOR2D1 U985 ( .A1(sa33_sr[7]), .A2(sa03_sr[7]), .Z(n203) );
  CKND1 U986 ( .I(sa33_sr[3]), .ZN(n569) );
  XOR4D2 U987 ( .A1(n107), .A2(n425), .A3(n534), .A4(n16), .Z(n500) );
  XNR3D4 U988 ( .A1(n107), .A2(n108), .A3(n670), .ZN(n106) );
  XOR2D4 U989 ( .A1(n93), .A2(n79), .Z(n107) );
  XOR2D2 U990 ( .A1(sa23_sr[7]), .A2(sa13_sr[7]), .Z(n155) );
  MOAI22D1 U991 ( .A1(net7021), .A2(n353), .B1(n563), .B2(net7013), .ZN(N198)
         );
  XNR2D1 U992 ( .A1(text_in_r[86]), .A2(n47), .ZN(n563) );
  CKBD0 U993 ( .I(sa02_sr[4]), .Z(n564) );
  XNR3D0 U994 ( .A1(w1[10]), .A2(sa31_sr[1]), .A3(sa21_sr[1]), .ZN(n394) );
  CKBD0 U995 ( .I(sa12_sr[6]), .Z(n565) );
  INVD1 U996 ( .I(n78), .ZN(n566) );
  CKXOR2D0 U997 ( .A1(w3[21]), .A2(sa13_sr[5]), .Z(N434) );
  XOR3D0 U998 ( .A1(sa13_sr[5]), .A2(n152), .A3(n180), .Z(n179) );
  XOR4D2 U999 ( .A1(n221), .A2(n254), .A3(sa00_sr[6]), .A4(n60), .Z(n300) );
  INVD1 U1000 ( .I(n567), .ZN(n568) );
  INVD1 U1001 ( .I(n569), .ZN(n570) );
  CKBD0 U1002 ( .I(sa21_sr[6]), .Z(n571) );
  CKND0 U1003 ( .I(sa22_sr[7]), .ZN(n572) );
  INVD1 U1004 ( .I(n572), .ZN(n573) );
  XOR3D2 U1005 ( .A1(w2[11]), .A2(sa32_sr[2]), .A3(sa22_sr[2]), .Z(n492) );
  CKND1 U1006 ( .I(n98), .ZN(n628) );
  XNR3D4 U1007 ( .A1(n360), .A2(n365), .A3(n660), .ZN(n364) );
  XOR4D0 U1008 ( .A1(n319), .A2(n376), .A3(sa11_sr[0]), .A4(n40), .Z(n399) );
  XNR3D4 U1009 ( .A1(n155), .A2(n160), .A3(n664), .ZN(n159) );
  XNR2D1 U1010 ( .A1(sa22_sr[3]), .A2(sa12_sr[3]), .ZN(n575) );
  XNR2D1 U1011 ( .A1(sa22_sr[3]), .A2(sa12_sr[3]), .ZN(n97) );
  XNR3D4 U1012 ( .A1(w0[19]), .A2(n646), .A3(n238), .ZN(n263) );
  MOAI22D1 U1013 ( .A1(net7025), .A2(n196), .B1(n576), .B2(net7015), .ZN(N39)
         );
  XNR2D1 U1014 ( .A1(text_in_r[7]), .A2(n11), .ZN(n576) );
  XOR2D0 U1015 ( .A1(w1[7]), .A2(sa31_sr[7]), .Z(N480) );
  XNR3D0 U1016 ( .A1(sa31_sr[7]), .A2(w1[15]), .A3(sa31_sr[6]), .ZN(n379) );
  XOR3D1 U1017 ( .A1(w2[4]), .A2(sa02_sr[4]), .A3(n98), .Z(n509) );
  XOR4D1 U1018 ( .A1(n331), .A2(n635), .A3(n559), .A4(n346), .Z(n344) );
  XOR2D2 U1019 ( .A1(sa11_sr[7]), .A2(sa21_sr[7]), .Z(n360) );
  CKND0 U1020 ( .I(sa22_sr[4]), .ZN(n598) );
  XOR3D2 U1021 ( .A1(w3[4]), .A2(n558), .A3(n128), .Z(n204) );
  XNR2D1 U1022 ( .A1(sa20_sr[1]), .A2(sa10_sr[1]), .ZN(n242) );
  XOR3D0 U1023 ( .A1(sa32_sr[4]), .A2(w2[13]), .A3(n599), .Z(n668) );
  MOAI22D1 U1024 ( .A1(net7021), .A2(n351), .B1(n577), .B2(net7013), .ZN(N199)
         );
  XNR2D1 U1025 ( .A1(text_in_r[87]), .A2(n48), .ZN(n577) );
  XOR3D2 U1026 ( .A1(w3[11]), .A2(sa33_sr[2]), .A3(sa23_sr[2]), .Z(n186) );
  CKXOR2D0 U1027 ( .A1(w3[8]), .A2(sa23_sr[0]), .Z(N471) );
  CKXOR2D0 U1028 ( .A1(w1[13]), .A2(sa21_sr[5]), .Z(N450) );
  MOAI22D1 U1029 ( .A1(n411), .A2(net7019), .B1(n578), .B2(net7013), .ZN(N163)
         );
  XNR2D1 U1030 ( .A1(text_in_r[67]), .A2(n35), .ZN(n578) );
  XOR2D0 U1031 ( .A1(w1[11]), .A2(n536), .Z(N452) );
  XOR2D0 U1032 ( .A1(w2[19]), .A2(sa12_sr[3]), .Z(N428) );
  ND2D0 U1033 ( .A1(sa20_sr[3]), .A2(sa10_sr[3]), .ZN(n678) );
  CKBD0 U1034 ( .I(sa00_sr[0]), .Z(n579) );
  XNR3D4 U1035 ( .A1(n614), .A2(n21), .A3(n103), .ZN(n475) );
  MOAI22D1 U1036 ( .A1(n375), .A2(net7019), .B1(n580), .B2(net7013), .ZN(N192)
         );
  XNR2D1 U1037 ( .A1(text_in_r[80]), .A2(n44), .ZN(n580) );
  XNR3D0 U1038 ( .A1(sa30_sr[1]), .A2(w0[10]), .A3(sa20_sr[1]), .ZN(n291) );
  CKBD0 U1039 ( .I(sa02_sr[6]), .Z(n581) );
  XOR4D0 U1040 ( .A1(n127), .A2(n132), .A3(n560), .A4(n133), .Z(n131) );
  INVD1 U1041 ( .I(n81), .ZN(n582) );
  CKND0 U1042 ( .I(sa33_sr[5]), .ZN(n583) );
  INVD1 U1043 ( .I(n583), .ZN(n584) );
  CKND1 U1044 ( .I(sa13_sr[3]), .ZN(n616) );
  CKXOR2D0 U1045 ( .A1(text_in_r[20]), .A2(w3[20]), .Z(n649) );
  XOR3D0 U1046 ( .A1(sa10_sr[6]), .A2(n251), .A3(n279), .Z(n278) );
  INVD0 U1047 ( .I(n625), .ZN(n626) );
  MOAI22D1 U1048 ( .A1(n401), .A2(net7019), .B1(n585), .B2(net7013), .ZN(N167)
         );
  XNR2D1 U1049 ( .A1(text_in_r[71]), .A2(n39), .ZN(n585) );
  CKXOR2D0 U1050 ( .A1(w1[29]), .A2(sa01_sr[5]), .Z(N386) );
  XOR3D0 U1051 ( .A1(sa01_sr[5]), .A2(n323), .A3(n324), .Z(n322) );
  MOAI22D1 U1052 ( .A1(net7021), .A2(n586), .B1(n587), .B2(net7015), .ZN(N36)
         );
  XOR3D4 U1053 ( .A1(n160), .A2(n203), .A3(n204), .Z(n586) );
  XNR2D1 U1054 ( .A1(text_in_r[4]), .A2(n8), .ZN(n587) );
  XNR3D1 U1055 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n618) );
  MOAI22D1 U1056 ( .A1(n348), .A2(net7021), .B1(n588), .B2(net7013), .ZN(N208)
         );
  XOR3D0 U1057 ( .A1(w1[31]), .A2(sa11_sr[6]), .A3(sa11_sr[7]), .Z(n658) );
  MOAI22D1 U1058 ( .A1(net7017), .A2(n457), .B1(n589), .B2(net7011), .ZN(N134)
         );
  XNR2D1 U1059 ( .A1(text_in_r[54]), .A2(n26), .ZN(n589) );
  XOR3D0 U1060 ( .A1(sa23_sr[1]), .A2(w3[17]), .A3(n144), .Z(n168) );
  CKXOR2D0 U1061 ( .A1(w2[30]), .A2(n581), .Z(N393) );
  MOAI22D1 U1062 ( .A1(net7023), .A2(n198), .B1(n590), .B2(net7025), .ZN(N38)
         );
  XNR2D1 U1063 ( .A1(text_in_r[6]), .A2(n10), .ZN(n590) );
  CKND0 U1064 ( .I(n79), .ZN(n591) );
  CKND2 U1065 ( .I(sa02_sr[0]), .ZN(n79) );
  CKXOR2D0 U1066 ( .A1(w2[22]), .A2(n565), .Z(N425) );
  XOR3D1 U1067 ( .A1(n155), .A2(n683), .A3(n168), .Z(n166) );
  MOAI22D1 U1068 ( .A1(net7021), .A2(n296), .B1(n592), .B2(net7013), .ZN(N240)
         );
  XNR2D1 U1069 ( .A1(text_in_r[104]), .A2(n62), .ZN(n592) );
  CKXOR2D0 U1070 ( .A1(w0[24]), .A2(n579), .Z(N383) );
  CKBD0 U1071 ( .I(sa23_sr[2]), .Z(n593) );
  MOAI22D1 U1072 ( .A1(net7025), .A2(n159), .B1(n594), .B2(net7015), .ZN(N67)
         );
  CKND0 U1073 ( .I(sa30_sr[1]), .ZN(n595) );
  INVD1 U1074 ( .I(n595), .ZN(n596) );
  MOAI22D1 U1075 ( .A1(net7023), .A2(n248), .B1(n597), .B2(net7015), .ZN(N263)
         );
  XNR2D1 U1076 ( .A1(text_in_r[119]), .A2(n70), .ZN(n597) );
  CKXOR2D0 U1077 ( .A1(w0[22]), .A2(sa10_sr[6]), .Z(N409) );
  INVD1 U1078 ( .I(n598), .ZN(n599) );
  CKXOR2D0 U1079 ( .A1(w1[27]), .A2(sa01_sr[3]), .Z(N388) );
  XOR3D4 U1080 ( .A1(n464), .A2(n469), .A3(n470), .Z(n468) );
  CKND1 U1081 ( .I(sa01_sr[4]), .ZN(n625) );
  CKND0 U1082 ( .I(sa30_sr[6]), .ZN(n600) );
  INVD1 U1083 ( .I(n600), .ZN(n601) );
  CKND0 U1084 ( .I(n90), .ZN(n602) );
  XOR3D2 U1085 ( .A1(w2[25]), .A2(sa12_sr[0]), .A3(sa32_sr[1]), .Z(n449) );
  XOR4D2 U1086 ( .A1(n112), .A2(n438), .A3(n93), .A4(w2[24]), .Z(n451) );
  MOAI22D1 U1087 ( .A1(n284), .A2(net7021), .B1(n603), .B2(net7015), .ZN(N244)
         );
  XOR3D2 U1088 ( .A1(w3[9]), .A2(sa33_sr[0]), .A3(sa23_sr[0]), .Z(n192) );
  CKXOR2D0 U1089 ( .A1(w3[0]), .A2(n526), .Z(N503) );
  MOAI22D1 U1090 ( .A1(net7025), .A2(n166), .B1(n604), .B2(net7015), .ZN(N65)
         );
  CKND0 U1091 ( .I(sa00_sr[2]), .ZN(n605) );
  INVD1 U1092 ( .I(n605), .ZN(n606) );
  XOR3D2 U1093 ( .A1(w2[3]), .A2(sa02_sr[3]), .A3(n100), .Z(n663) );
  CKND0 U1094 ( .I(sa02_sr[1]), .ZN(n607) );
  INVD1 U1095 ( .I(n607), .ZN(n608) );
  XOR2D0 U1096 ( .A1(n711), .A2(n570), .Z(N500) );
  XOR3D2 U1097 ( .A1(w3[27]), .A2(sa13_sr[2]), .A3(sa33_sr[3]), .Z(n133) );
  CKBD0 U1098 ( .I(n568), .Z(n609) );
  XOR4D1 U1099 ( .A1(n331), .A2(sa01_sr[3]), .A3(n332), .A4(n333), .Z(n330) );
  CKND0 U1100 ( .I(n91), .ZN(n610) );
  XOR3D2 U1101 ( .A1(w2[12]), .A2(sa32_sr[3]), .A3(sa22_sr[3]), .Z(n489) );
  XOR3D2 U1102 ( .A1(w2[27]), .A2(sa12_sr[2]), .A3(n549), .Z(n443) );
  CKXOR2D0 U1103 ( .A1(w2[15]), .A2(n573), .Z(N456) );
  XOR4D2 U1104 ( .A1(n360), .A2(n376), .A3(n548), .A4(n44), .Z(n375) );
  CKND0 U1105 ( .I(sa23_sr[7]), .ZN(n612) );
  INVD1 U1106 ( .I(n612), .ZN(n613) );
  BUFFD2 U1107 ( .I(sa22_sr[1]), .Z(n614) );
  XOR4D2 U1108 ( .A1(n155), .A2(n171), .A3(sa23_sr[0]), .A4(w3[16]), .Z(n170)
         );
  XOR3D4 U1109 ( .A1(n273), .A2(n305), .A3(n314), .Z(n615) );
  OAI22D2 U1110 ( .A1(n432), .A2(net7005), .B1(net7019), .B2(n433), .ZN(N149)
         );
  INVD1 U1111 ( .I(n616), .ZN(n617) );
  MOAI22D1 U1112 ( .A1(n255), .A2(net6997), .B1(net7007), .B2(n618), .ZN(N260)
         );
  CKND0 U1113 ( .I(sa23_sr[1]), .ZN(n91) );
  MOAI22D1 U1114 ( .A1(n619), .A2(net7021), .B1(n620), .B2(net7011), .ZN(N164)
         );
  XOR3D1 U1115 ( .A1(n365), .A2(n408), .A3(n409), .Z(n619) );
  XOR3D2 U1116 ( .A1(w0[9]), .A2(sa20_sr[0]), .A3(n520), .Z(n294) );
  CKXOR2D0 U1117 ( .A1(w0[0]), .A2(n520), .Z(N479) );
  CKBD1 U1118 ( .I(sa12_sr[1]), .Z(n639) );
  CKND0 U1119 ( .I(sa00_sr[4]), .ZN(n621) );
  INVD1 U1120 ( .I(n621), .ZN(n622) );
  CKND0 U1121 ( .I(sa20_sr[4]), .ZN(n623) );
  INVD1 U1122 ( .I(n623), .ZN(n624) );
  MOAI22D1 U1123 ( .A1(net7023), .A2(n268), .B1(n627), .B2(net7015), .ZN(N257)
         );
  XNR2D1 U1124 ( .A1(text_in_r[113]), .A2(n67), .ZN(n627) );
  INVD1 U1125 ( .I(n628), .ZN(n629) );
  CKXOR2D1 U1126 ( .A1(sa32_sr[7]), .A2(n80), .Z(n98) );
  XOR4D0 U1127 ( .A1(n575), .A2(n438), .A3(sa02_sr[2]), .A4(n443), .Z(n442) );
  XOR3D4 U1128 ( .A1(w2[20]), .A2(sa22_sr[4]), .A3(n97), .Z(n466) );
  CKND0 U1129 ( .I(n93), .ZN(n630) );
  XOR3D1 U1130 ( .A1(n156), .A2(n155), .A3(n157), .Z(n672) );
  CKXOR2D0 U1131 ( .A1(w2[5]), .A2(sa32_sr[5]), .Z(N490) );
  CKXOR2D0 U1132 ( .A1(w0[27]), .A2(sa00_sr[3]), .Z(N380) );
  XNR2D1 U1133 ( .A1(sa23_sr[1]), .A2(sa13_sr[1]), .ZN(n140) );
  XOR4D2 U1134 ( .A1(n107), .A2(n464), .A3(sa22_sr[0]), .A4(n20), .Z(n477) );
  MOAI22D1 U1135 ( .A1(net7025), .A2(n163), .B1(n631), .B2(net7015), .ZN(N66)
         );
  XOR3D1 U1136 ( .A1(w0[12]), .A2(sa30_sr[3]), .A3(sa20_sr[3]), .Z(n285) );
  CKXOR2D0 U1137 ( .A1(w2[12]), .A2(n599), .Z(N459) );
  MOAI22D1 U1138 ( .A1(n200), .A2(net7023), .B1(n632), .B2(net7015), .ZN(N37)
         );
  XNR2D1 U1139 ( .A1(text_in_r[5]), .A2(n9), .ZN(n632) );
  CKND0 U1140 ( .I(n88), .ZN(n633) );
  CKND0 U1141 ( .I(sa11_sr[4]), .ZN(n88) );
  XOR2D2 U1142 ( .A1(sa13_sr[7]), .A2(sa03_sr[7]), .Z(n127) );
  CKND0 U1143 ( .I(sa01_sr[0]), .ZN(n634) );
  INVD1 U1144 ( .I(n634), .ZN(n635) );
  MOAI22D1 U1145 ( .A1(net7019), .A2(n399), .B1(n636), .B2(net7013), .ZN(N176)
         );
  XNR2D1 U1146 ( .A1(text_in_r[72]), .A2(n40), .ZN(n636) );
  MOAI22D1 U1147 ( .A1(n214), .A2(net7023), .B1(n640), .B2(net7013), .ZN(N32)
         );
  MOAI22D1 U1148 ( .A1(net7019), .A2(n371), .B1(n641), .B2(net7013), .ZN(N193)
         );
  XNR2D1 U1149 ( .A1(text_in_r[81]), .A2(n45), .ZN(n641) );
  MOAI22D1 U1150 ( .A1(n642), .A2(net7005), .B1(net7005), .B2(n643), .ZN(N259)
         );
  XNR2D1 U1151 ( .A1(text_in_r[115]), .A2(w0[19]), .ZN(n642) );
  XNR3D1 U1152 ( .A1(n257), .A2(n262), .A3(n263), .ZN(n643) );
  MOAI22D1 U1153 ( .A1(net7025), .A2(n194), .B1(n644), .B2(net7015), .ZN(N48)
         );
  MOAI22D1 U1154 ( .A1(net7023), .A2(n265), .B1(n645), .B2(net7013), .ZN(N258)
         );
  OAI22D2 U1155 ( .A1(n363), .A2(net7001), .B1(net7019), .B2(n364), .ZN(N195)
         );
  MOAI22D1 U1156 ( .A1(n185), .A2(net7025), .B1(n542), .B2(net7015), .ZN(N51)
         );
  XOR4D2 U1157 ( .A1(n108), .A2(n100), .A3(sa22_sr[2]), .A4(n22), .Z(n472) );
  XOR3D4 U1158 ( .A1(n112), .A2(n464), .A3(n475), .Z(n474) );
  OAI22D2 U1159 ( .A1(n467), .A2(net7007), .B1(net7017), .B2(n468), .ZN(N131)
         );
  INVD1 U1160 ( .I(n676), .ZN(n646) );
  XOR3D2 U1161 ( .A1(w3[28]), .A2(sa33_sr[4]), .A3(n617), .Z(n129) );
  MOAI22D1 U1162 ( .A1(net7023), .A2(n245), .B1(n647), .B2(net7013), .ZN(N272)
         );
  INVD1 U1163 ( .I(w3[7]), .ZN(n11) );
  INVD1 U1164 ( .I(net7015), .ZN(net6993) );
  CKBD1 U1165 ( .I(net7033), .Z(net7025) );
  XOR3D0 U1166 ( .A1(sa13_sr[6]), .A2(n149), .A3(n177), .Z(n176) );
  MOAI22D1 U1167 ( .A1(n211), .A2(net7023), .B1(n648), .B2(net7015), .ZN(N33)
         );
  XNR2D1 U1168 ( .A1(text_in_r[1]), .A2(n710), .ZN(n648) );
  CKXOR2D0 U1169 ( .A1(w2[23]), .A2(sa12_sr[7]), .Z(N424) );
  XOR4D2 U1170 ( .A1(n257), .A2(n273), .A3(sa20_sr[0]), .A4(n66), .Z(n272) );
  XOR3D2 U1171 ( .A1(w0[25]), .A2(sa30_sr[1]), .A3(n574), .Z(n243) );
  XOR3D4 U1172 ( .A1(n164), .A2(n203), .A3(n207), .Z(n206) );
  XOR3D2 U1173 ( .A1(w1[12]), .A2(sa31_sr[3]), .A3(sa21_sr[3]), .Z(n388) );
  XOR3D2 U1174 ( .A1(w1[27]), .A2(sa31_sr[3]), .A3(n675), .Z(n337) );
  OAI22D2 U1175 ( .A1(n205), .A2(net6995), .B1(n206), .B2(net7023), .ZN(N35)
         );
  XOR2D0 U1176 ( .A1(w1[5]), .A2(sa31_sr[5]), .Z(N482) );
  MOAI22D1 U1177 ( .A1(n672), .A2(net7025), .B1(n649), .B2(net7015), .ZN(N68)
         );
  XOR4D2 U1178 ( .A1(n327), .A2(n354), .A3(n571), .A4(n47), .Z(n353) );
  XOR2D0 U1179 ( .A1(w2[25]), .A2(n608), .Z(N398) );
  XOR3D0 U1180 ( .A1(w2[15]), .A2(sa32_sr[7]), .A3(sa32_sr[6]), .Z(n666) );
  CKND0 U1181 ( .I(sa00_sr[1]), .ZN(n650) );
  INVD1 U1182 ( .I(n650), .ZN(n651) );
  XOR2D2 U1183 ( .A1(sa31_sr[7]), .A2(sa21_sr[7]), .Z(n319) );
  XOR3D2 U1184 ( .A1(w0[1]), .A2(n651), .A3(n242), .Z(n314) );
  CKXOR2D0 U1185 ( .A1(w0[25]), .A2(n651), .Z(N382) );
  MOAI22D1 U1186 ( .A1(n111), .A2(net7025), .B1(n652), .B2(net7017), .ZN(N96)
         );
  XOR3D2 U1187 ( .A1(w2[28]), .A2(sa32_sr[4]), .A3(sa12_sr[3]), .Z(n440) );
  MOAI22D1 U1188 ( .A1(n241), .A2(net7023), .B1(n653), .B2(net7015), .ZN(N273)
         );
  XOR2D0 U1189 ( .A1(w1[19]), .A2(n547), .Z(N420) );
  XOR3D2 U1190 ( .A1(w1[28]), .A2(sa31_sr[4]), .A3(sa11_sr[3]), .Z(n333) );
  XNR2D0 U1191 ( .A1(text_in_r[29]), .A2(w3[29]), .ZN(n121) );
  XNR3D4 U1192 ( .A1(n575), .A2(n629), .A3(n663), .ZN(n96) );
  MOAI22D1 U1193 ( .A1(n293), .A2(net7021), .B1(n654), .B2(net7013), .ZN(N241)
         );
  CKXOR2D0 U1194 ( .A1(w2[31]), .A2(sa02_sr[7]), .Z(N392) );
  XOR3D2 U1195 ( .A1(w3[26]), .A2(n674), .A3(sa13_sr[1]), .Z(n665) );
  XNR2D0 U1196 ( .A1(text_in_r[26]), .A2(w3[26]), .ZN(n134) );
  CKXOR2D0 U1197 ( .A1(w3[26]), .A2(n560), .Z(N405) );
  OAI22D2 U1198 ( .A1(n95), .A2(net6999), .B1(net7025), .B2(n96), .ZN(N99) );
  XOR3D2 U1199 ( .A1(w1[9]), .A2(sa31_sr[0]), .A3(sa21_sr[0]), .Z(n397) );
  CKXOR2D0 U1200 ( .A1(w3[16]), .A2(sa13_sr[0]), .Z(N439) );
  CKND2 U1201 ( .I(sa13_sr[0]), .ZN(n82) );
  XOR2D0 U1202 ( .A1(w1[2]), .A2(sa31_sr[2]), .Z(N485) );
  XOR3D2 U1203 ( .A1(w1[11]), .A2(sa31_sr[2]), .A3(sa21_sr[2]), .Z(n391) );
  MOAI22D1 U1204 ( .A1(net7025), .A2(n139), .B1(n655), .B2(net7017), .ZN(N81)
         );
  XOR2D0 U1205 ( .A1(w0[2]), .A2(sa30_sr[2]), .Z(N477) );
  XOR3D4 U1206 ( .A1(n171), .A2(n203), .A3(n212), .Z(n211) );
  XOR2D0 U1207 ( .A1(w0[7]), .A2(sa30_sr[7]), .Z(N472) );
  XOR2D2 U1208 ( .A1(sa30_sr[7]), .A2(sa20_sr[7]), .Z(n217) );
  CKND1 U1209 ( .I(sa03_sr[1]), .ZN(n656) );
  XOR3D2 U1210 ( .A1(w1[25]), .A2(sa31_sr[1]), .A3(sa11_sr[0]), .Z(n346) );
  CKXOR2D0 U1211 ( .A1(w3[10]), .A2(n593), .Z(N469) );
  XNR3D0 U1212 ( .A1(w2[26]), .A2(sa32_sr[2]), .A3(n639), .ZN(n446) );
  XOR2D0 U1213 ( .A1(w2[2]), .A2(sa32_sr[2]), .Z(N493) );
  XOR4D0 U1214 ( .A1(n217), .A2(sa10_sr[3]), .A3(n262), .A4(n288), .Z(n287) );
  XOR3D0 U1215 ( .A1(sa00_sr[5]), .A2(n221), .A3(n222), .Z(n220) );
  XOR3D1 U1216 ( .A1(sa20_sr[6]), .A2(n229), .A3(n276), .Z(n275) );
  XNR3D0 U1217 ( .A1(sa02_sr[5]), .A2(n429), .A3(n662), .ZN(n428) );
  XOR3D0 U1218 ( .A1(sa12_sr[7]), .A2(w2[31]), .A3(n565), .Z(n661) );
  CKND1 U1219 ( .I(sa02_sr[7]), .ZN(n80) );
  CKND0 U1220 ( .I(sa01_sr[7]), .ZN(n78) );
  XNR3D0 U1221 ( .A1(sa01_sr[6]), .A2(n319), .A3(n658), .ZN(n318) );
  XOR4D0 U1222 ( .A1(n246), .A2(n305), .A3(sa00_sr[0]), .A4(w0[0]), .Z(n316)
         );
  XOR4D0 U1223 ( .A1(n229), .A2(n246), .A3(n520), .A4(w0[24]), .Z(n245) );
  XNR3D0 U1224 ( .A1(sa00_sr[6]), .A2(n217), .A3(n659), .ZN(n216) );
  CKND0 U1225 ( .I(w3[6]), .ZN(n10) );
  XNR3D0 U1226 ( .A1(w0[14]), .A2(sa30_sr[5]), .A3(sa20_sr[5]), .ZN(n279) );
  XNR3D0 U1227 ( .A1(n581), .A2(n425), .A3(n661), .ZN(n424) );
  XOR3D0 U1228 ( .A1(sa11_sr[6]), .A2(n354), .A3(n382), .Z(n381) );
  XOR4D0 U1229 ( .A1(n127), .A2(n140), .A3(n673), .A4(n141), .Z(n139) );
  XNR3D0 U1230 ( .A1(w3[14]), .A2(sa33_sr[5]), .A3(sa23_sr[5]), .ZN(n177) );
  XOR4D0 U1231 ( .A1(n544), .A2(n349), .A3(n530), .A4(w1[24]), .Z(n348) );
  XOR4D0 U1232 ( .A1(n425), .A2(n429), .A3(n80), .A4(w2[23]), .Z(n455) );
  XNR3D0 U1233 ( .A1(sa22_sr[6]), .A2(n691), .A3(n666), .ZN(n479) );
  XNR3D0 U1234 ( .A1(n543), .A2(n100), .A3(n667), .ZN(n494) );
  XNR3D1 U1235 ( .A1(sa12_sr[5]), .A2(n461), .A3(n668), .ZN(n485) );
  XNR3D0 U1236 ( .A1(n565), .A2(n458), .A3(n669), .ZN(n482) );
  XOR4D0 U1237 ( .A1(n544), .A2(n354), .A3(sa21_sr[7]), .A4(n39), .Z(n401) );
  XOR4D0 U1238 ( .A1(n319), .A2(n372), .A3(n87), .A4(n397), .Z(n396) );
  XOR2D0 U1239 ( .A1(text_in_r[24]), .A2(w3[24]), .Z(n684) );
  XOR2D0 U1240 ( .A1(text_in_r[27]), .A2(w3[27]), .Z(n671) );
  XOR2D0 U1241 ( .A1(text_in_r[28]), .A2(w3[28]), .Z(n696) );
  XOR4D1 U1242 ( .A1(n115), .A2(n609), .A3(n156), .A4(n183), .Z(n182) );
  XOR4D0 U1243 ( .A1(w2[2]), .A2(n104), .A3(sa02_sr[2]), .A4(n103), .Z(n102)
         );
  XOR3D0 U1244 ( .A1(sa03_sr[5]), .A2(n119), .A3(n120), .Z(n118) );
  XNR3D0 U1245 ( .A1(sa30_sr[6]), .A2(w0[30]), .A3(sa10_sr[5]), .ZN(n222) );
  XOR2D0 U1246 ( .A1(w0[3]), .A2(sa30_sr[3]), .Z(N476) );
  CKBD1 U1247 ( .I(n438), .Z(n691) );
  CKXOR2D1 U1248 ( .A1(sa12_sr[7]), .A2(sa02_sr[7]), .Z(n438) );
  CKXOR2D1 U1249 ( .A1(n85), .A2(sa20_sr[4]), .Z(n230) );
  XNR2D1 U1250 ( .A1(sa21_sr[4]), .A2(sa11_sr[4]), .ZN(n332) );
  CKXOR2D1 U1251 ( .A1(sa12_sr[1]), .A2(sa22_sr[1]), .Z(n108) );
  XNR2D1 U1252 ( .A1(sa20_sr[0]), .A2(sa10_sr[0]), .ZN(n246) );
  XNR2D1 U1253 ( .A1(sa23_sr[3]), .A2(sa13_sr[3]), .ZN(n132) );
  INVD1 U1254 ( .I(net7013), .ZN(net6999) );
  INVD1 U1255 ( .I(net7011), .ZN(net7007) );
  INVD1 U1256 ( .I(net7013), .ZN(net7003) );
  INVD1 U1257 ( .I(net7015), .ZN(net6997) );
  INVD1 U1258 ( .I(net7011), .ZN(net7009) );
  INVD1 U1259 ( .I(net7015), .ZN(net6995) );
  INVD1 U1260 ( .I(net7017), .ZN(net6991) );
  INVD1 U1261 ( .I(net7011), .ZN(net7005) );
  INVD1 U1262 ( .I(net7013), .ZN(net7001) );
  INVD1 U1263 ( .I(n712), .ZN(n711) );
  CKBD1 U1264 ( .I(net7027), .Z(net7011) );
  CKBD1 U1265 ( .I(net7029), .Z(net7017) );
  CKBD1 U1266 ( .I(net7031), .Z(net7019) );
  CKBD1 U1267 ( .I(net7033), .Z(net7023) );
  CKBD1 U1268 ( .I(net7027), .Z(net7013) );
  CKBD1 U1269 ( .I(net7029), .Z(net7015) );
  CKBD1 U1270 ( .I(net7031), .Z(net7021) );
  INVD1 U1271 ( .I(n453), .ZN(n3) );
  INVD1 U1272 ( .I(w3[3]), .ZN(n712) );
  OAI211D1 U1273 ( .A1(dcnt[3]), .A2(n2), .B(n713), .C(rst), .ZN(n420) );
  INVD1 U1274 ( .I(n421), .ZN(n2) );
  ND3D1 U1275 ( .A1(n420), .A2(n713), .A3(rst), .ZN(N12) );
  INVD1 U1276 ( .I(w1[16]), .ZN(n44) );
  INVD1 U1277 ( .I(w0[5]), .ZN(n59) );
  XNR2D1 U1278 ( .A1(text_in_r[56]), .A2(w2[24]), .ZN(n450) );
  INVD1 U1279 ( .I(w0[16]), .ZN(n66) );
  INVD1 U1280 ( .I(w1[22]), .ZN(n47) );
  INVD1 U1281 ( .I(w0[6]), .ZN(n60) );
  XNR2D1 U1282 ( .A1(text_in_r[93]), .A2(w1[29]), .ZN(n325) );
  XNR2D1 U1283 ( .A1(text_in_r[90]), .A2(w1[26]), .ZN(n338) );
  INVD1 U1284 ( .I(w0[8]), .ZN(n62) );
  INVD1 U1285 ( .I(w2[7]), .ZN(n15) );
  INVD1 U1286 ( .I(w0[22]), .ZN(n69) );
  NR2D1 U1287 ( .A1(n3), .A2(dcnt[2]), .ZN(n421) );
  OAI31D1 U1288 ( .A1(n420), .A2(n421), .A3(n1), .B(n422), .ZN(N16) );
  INVD1 U1289 ( .I(dcnt[3]), .ZN(n1) );
  NR4D0 U1290 ( .A1(n342), .A2(dcnt[2]), .A3(ld), .A4(dcnt[3]), .ZN(N21) );
  IND2D1 U1291 ( .A1(dcnt[1]), .B1(dcnt[0]), .ZN(n342) );
  INVD1 U1292 ( .I(w2[8]), .ZN(n16) );
  INVD1 U1293 ( .I(w1[7]), .ZN(n39) );
  CKXOR2D1 U1294 ( .A1(text_in_r[92]), .A2(w1[28]), .Z(n700) );
  INVD1 U1295 ( .I(w1[8]), .ZN(n40) );
  INVD1 U1296 ( .I(w0[23]), .ZN(n70) );
  OAI22D1 U1297 ( .A1(n454), .A2(net7007), .B1(n455), .B2(net7017), .ZN(N135)
         );
  INVD1 U1298 ( .I(w2[23]), .ZN(n27) );
  INVD1 U1299 ( .I(w1[23]), .ZN(n48) );
  INVD1 U1300 ( .I(w2[16]), .ZN(n20) );
  INVD1 U1301 ( .I(w0[7]), .ZN(n61) );
  OAI22D1 U1302 ( .A1(n402), .A2(net7003), .B1(n403), .B2(net7019), .ZN(N166)
         );
  INVD1 U1303 ( .I(w1[6]), .ZN(n38) );
  OAI22D1 U1304 ( .A1(n503), .A2(net7009), .B1(net7015), .B2(n504), .ZN(N102)
         );
  INVD1 U1305 ( .I(w2[6]), .ZN(n14) );
  INVD1 U1306 ( .I(w2[22]), .ZN(n26) );
  OAI22D1 U1307 ( .A1(n223), .A2(net6995), .B1(net7023), .B2(n224), .ZN(N277)
         );
  INVD1 U1308 ( .I(w0[29]), .ZN(n75) );
  INVD1 U1309 ( .I(w0[26]), .ZN(n72) );
  OAI22D1 U1310 ( .A1(n444), .A2(net7005), .B1(net7019), .B2(n445), .ZN(N146)
         );
  OAI22D1 U1311 ( .A1(n121), .A2(net6991), .B1(net7025), .B2(n122), .ZN(N85)
         );
  OAI22D1 U1312 ( .A1(n178), .A2(net6993), .B1(net7025), .B2(n179), .ZN(N53)
         );
  OAI22D1 U1313 ( .A1(n105), .A2(net6991), .B1(net7025), .B2(n106), .ZN(N97)
         );
  OAI22D1 U1314 ( .A1(n187), .A2(net6993), .B1(net7025), .B2(n188), .ZN(N50)
         );
  INVD1 U1315 ( .I(w2[19]), .ZN(n23) );
  INVD1 U1316 ( .I(w2[20]), .ZN(n24) );
  OAI22D1 U1317 ( .A1(n427), .A2(net7005), .B1(net7019), .B2(n428), .ZN(N150)
         );
  INVD1 U1318 ( .I(w2[29]), .ZN(n32) );
  OAI22D1 U1319 ( .A1(n423), .A2(net7005), .B1(net7019), .B2(n424), .ZN(N151)
         );
  OAI22D1 U1320 ( .A1(n321), .A2(net6999), .B1(net7021), .B2(n322), .ZN(N214)
         );
  INVD1 U1321 ( .I(w1[30]), .ZN(n54) );
  OAI22D1 U1322 ( .A1(n317), .A2(net6999), .B1(net7021), .B2(n318), .ZN(N215)
         );
  OAI22D1 U1323 ( .A1(n274), .A2(net6997), .B1(net7023), .B2(n275), .ZN(N247)
         );
  OAI22D1 U1324 ( .A1(n219), .A2(net6995), .B1(net7023), .B2(n220), .ZN(N278)
         );
  INVD1 U1325 ( .I(w0[30]), .ZN(n76) );
  INVD1 U1326 ( .I(w0[17]), .ZN(n67) );
  OAI22D1 U1327 ( .A1(n215), .A2(net6995), .B1(net7023), .B2(n216), .ZN(N279)
         );
  OAI22D1 U1328 ( .A1(n383), .A2(net7003), .B1(net7019), .B2(n384), .ZN(N181)
         );
  XOR3D1 U1329 ( .A1(sa11_sr[5]), .A2(n357), .A3(n385), .Z(n384) );
  OAI22D1 U1330 ( .A1(n478), .A2(net7007), .B1(net7017), .B2(n479), .ZN(N119)
         );
  INVD1 U1331 ( .I(w2[4]), .ZN(n12) );
  OAI22D1 U1332 ( .A1(n413), .A2(net7005), .B1(net7019), .B2(n414), .ZN(N162)
         );
  OAI22D1 U1333 ( .A1(n392), .A2(net7003), .B1(net7019), .B2(n393), .ZN(N178)
         );
  INVD1 U1334 ( .I(w1[3]), .ZN(n35) );
  INVD1 U1335 ( .I(w0[1]), .ZN(n55) );
  INVD1 U1336 ( .I(w0[3]), .ZN(n57) );
  INVD1 U1337 ( .I(w1[17]), .ZN(n45) );
  INVD1 U1338 ( .I(w2[17]), .ZN(n21) );
  INVD1 U1339 ( .I(w3[4]), .ZN(n8) );
  INVD1 U1340 ( .I(w0[4]), .ZN(n58) );
  XNR2D1 U1341 ( .A1(text_in_r[107]), .A2(w0[11]), .ZN(n286) );
  CKXOR2D1 U1342 ( .A1(text_in_r[85]), .A2(w1[21]), .Z(n687) );
  INVD1 U1343 ( .I(w2[11]), .ZN(n18) );
  CKXOR2D1 U1344 ( .A1(text_in_r[41]), .A2(w2[9]), .Z(n698) );
  CKXOR2D1 U1345 ( .A1(text_in_r[59]), .A2(w2[27]), .Z(n682) );
  CKXOR2D1 U1346 ( .A1(text_in_r[57]), .A2(w2[25]), .Z(n702) );
  CKXOR2D1 U1347 ( .A1(text_in_r[124]), .A2(w0[28]), .Z(n701) );
  CKXOR2D1 U1348 ( .A1(text_in_r[117]), .A2(w0[21]), .Z(n699) );
  CKXOR2D1 U1349 ( .A1(text_in_r[44]), .A2(w2[12]), .Z(n693) );
  CKXOR2D1 U1350 ( .A1(text_in_r[91]), .A2(w1[27]), .Z(n689) );
  NR2D1 U1351 ( .A1(dcnt[1]), .A2(dcnt[0]), .ZN(n453) );
  INVD1 U1352 ( .I(w2[21]), .ZN(n25) );
  CKXOR2D1 U1353 ( .A1(text_in_r[73]), .A2(w1[9]), .Z(n697) );
  CKXOR2D1 U1354 ( .A1(text_in_r[89]), .A2(w1[25]), .Z(n708) );
  INVD1 U1355 ( .I(w2[18]), .ZN(n22) );
  CKXOR2D1 U1356 ( .A1(text_in_r[76]), .A2(w1[12]), .Z(n686) );
  CKXOR2D1 U1357 ( .A1(text_in_r[64]), .A2(w1[0]), .Z(n688) );
  INVD1 U1358 ( .I(w0[2]), .ZN(n56) );
  CKXOR2D1 U1359 ( .A1(text_in_r[123]), .A2(w0[27]), .Z(n704) );
  INVD1 U1360 ( .I(w2[5]), .ZN(n13) );
  INVD1 U1361 ( .I(w1[5]), .ZN(n37) );
  CKXOR2D1 U1362 ( .A1(text_in_r[65]), .A2(w1[1]), .Z(n709) );
  ND2D1 U1363 ( .A1(ld), .A2(rst), .ZN(n422) );
  OAI21D1 U1364 ( .A1(n452), .A2(n420), .B(n422), .ZN(N14) );
  AOI21D1 U1365 ( .A1(dcnt[1]), .A2(dcnt[0]), .B(n453), .ZN(n452) );
  OAI21D1 U1366 ( .A1(dcnt[0]), .A2(n420), .B(n422), .ZN(N13) );
  XOR3D1 U1367 ( .A1(sa01_sr[3]), .A2(w1[3]), .A3(n336), .Z(n412) );
  OAI22D1 U1368 ( .A1(n117), .A2(net6991), .B1(net7025), .B2(n118), .ZN(N86)
         );
  INVD1 U1369 ( .I(w0[20]), .ZN(n68) );
  XOR3D1 U1370 ( .A1(w0[4]), .A2(n622), .A3(n230), .Z(n306) );
  XOR3D1 U1371 ( .A1(w1[29]), .A2(sa31_sr[5]), .A3(n88), .Z(n328) );
  XOR3D1 U1372 ( .A1(w0[17]), .A2(sa20_sr[1]), .A3(n246), .Z(n270) );
  OAI22D1 U1373 ( .A1(n280), .A2(net6997), .B1(net7021), .B2(n281), .ZN(N245)
         );
  XOR3D1 U1374 ( .A1(sa10_sr[5]), .A2(n254), .A3(n282), .Z(n281) );
  XNR3D0 U1375 ( .A1(w0[13]), .A2(sa30_sr[4]), .A3(n624), .ZN(n282) );
  OAI22D1 U1376 ( .A1(n175), .A2(net6993), .B1(net7025), .B2(n176), .ZN(N54)
         );
  OAI22D1 U1377 ( .A1(n481), .A2(net7007), .B1(net7017), .B2(n482), .ZN(N118)
         );
  OAI22D1 U1378 ( .A1(n277), .A2(net6997), .B1(net7023), .B2(n278), .ZN(N246)
         );
  OAI22D1 U1379 ( .A1(n380), .A2(net7003), .B1(net7019), .B2(n381), .ZN(N182)
         );
  XOR3D1 U1380 ( .A1(w0[29]), .A2(sa30_sr[5]), .A3(n681), .Z(n226) );
  NR2D1 U1381 ( .A1(n431), .A2(n420), .ZN(N15) );
  AOI21D1 U1382 ( .A1(dcnt[2]), .A2(n3), .B(n421), .ZN(n431) );
  INVD1 U1383 ( .I(ld), .ZN(n713) );
  CKBD1 U1384 ( .I(ld_r), .Z(net7033) );
  CKBD1 U1385 ( .I(ld_r), .Z(net7031) );
  CKBD1 U1386 ( .I(ld_r), .Z(net7029) );
  CKBD1 U1387 ( .I(ld_r), .Z(net7027) );
  INVD1 U1388 ( .I(w1[11]), .ZN(n42) );
  INVD1 U1389 ( .I(w2[28]), .ZN(n31) );
  XNR2D1 U1390 ( .A1(w2[4]), .A2(n690), .ZN(N491) );
  CKXOR2D0 U1391 ( .A1(w3[7]), .A2(sa33_sr[7]), .Z(N496) );
  XOR3D1 U1392 ( .A1(n372), .A2(n695), .A3(n340), .Z(n414) );
  CKXOR2D0 U1393 ( .A1(w1[6]), .A2(sa31_sr[6]), .Z(N481) );
  BUFFD1 U1394 ( .I(sa03_sr[0]), .Z(n673) );
  CKBD1 U1395 ( .I(sa33_sr[2]), .Z(n674) );
  CKXOR2D0 U1396 ( .A1(w1[17]), .A2(sa11_sr[1]), .Z(N422) );
  CKND1 U1397 ( .I(sa11_sr[1]), .ZN(n87) );
  XOR3D1 U1398 ( .A1(n675), .A2(n369), .A3(n394), .Z(n393) );
  XOR2D0 U1399 ( .A1(w2[16]), .A2(n534), .Z(N431) );
  OAI22D1 U1400 ( .A1(n113), .A2(net6991), .B1(net7025), .B2(n114), .ZN(N87)
         );
  OAI22D1 U1401 ( .A1(n172), .A2(net6993), .B1(net7025), .B2(n173), .ZN(N55)
         );
  CKXOR2D0 U1402 ( .A1(w1[15]), .A2(sa21_sr[7]), .Z(N448) );
  XOR2D0 U1403 ( .A1(w3[24]), .A2(n673), .Z(N407) );
  XOR4D0 U1404 ( .A1(n136), .A2(n167), .A3(n560), .A4(n6), .Z(n209) );
  XOR4D0 U1405 ( .A1(n164), .A2(n593), .A3(n140), .A4(w3[18]), .Z(n163) );
  XOR3D1 U1406 ( .A1(sa23_sr[6]), .A2(n127), .A3(n174), .Z(n173) );
  CKND2D1 U1407 ( .A1(n676), .A2(n677), .ZN(n679) );
  ND2D1 U1408 ( .A1(n678), .A2(n679), .ZN(n234) );
  CKXOR2D0 U1409 ( .A1(w3[23]), .A2(sa13_sr[7]), .Z(N432) );
  XOR4D0 U1410 ( .A1(w1[21]), .A2(n357), .A3(sa21_sr[5]), .A4(n332), .Z(n356)
         );
  CKXOR2D0 U1411 ( .A1(w1[0]), .A2(n530), .Z(N487) );
  CKND0 U1412 ( .I(n85), .ZN(n680) );
  INVD1 U1413 ( .I(n680), .ZN(n681) );
  CKND1 U1414 ( .I(sa10_sr[4]), .ZN(n85) );
  OAI22D1 U1415 ( .A1(n493), .A2(net7007), .B1(net7017), .B2(n494), .ZN(N114)
         );
  XOR2D0 U1416 ( .A1(w0[19]), .A2(sa10_sr[3]), .Z(N412) );
  XNR2D0 U1417 ( .A1(text_in_r[9]), .A2(w3[9]), .ZN(n190) );
  MOAI22D1 U1418 ( .A1(n442), .A2(net7019), .B1(n682), .B2(net7011), .ZN(N147)
         );
  CKXOR2D1 U1419 ( .A1(n657), .A2(sa33_sr[1]), .Z(n167) );
  CKXOR2D0 U1420 ( .A1(w1[24]), .A2(n635), .Z(N391) );
  CKXOR2D0 U1421 ( .A1(w3[2]), .A2(n674), .Z(N501) );
  CKND0 U1422 ( .I(w3[2]), .ZN(n6) );
  MOAI22D1 U1423 ( .A1(net7025), .A2(n143), .B1(n684), .B2(net7017), .ZN(N80)
         );
  XOR2D0 U1424 ( .A1(w3[31]), .A2(n582), .Z(N400) );
  CKND0 U1425 ( .I(sa03_sr[7]), .ZN(n81) );
  CKXOR2D0 U1426 ( .A1(w3[19]), .A2(n617), .Z(N436) );
  XOR2D0 U1427 ( .A1(w0[8]), .A2(sa20_sr[0]), .Z(N447) );
  MOAI22D1 U1428 ( .A1(n506), .A2(net7013), .B1(n685), .B2(net7011), .ZN(N101)
         );
  XNR2D1 U1429 ( .A1(text_in_r[37]), .A2(n13), .ZN(n685) );
  XOR4D1 U1430 ( .A1(n79), .A2(n438), .A3(n108), .A4(n449), .Z(n448) );
  MOAI22D1 U1431 ( .A1(n387), .A2(net7019), .B1(n686), .B2(net7013), .ZN(N180)
         );
  MOAI22D1 U1432 ( .A1(net7021), .A2(n356), .B1(n687), .B2(net7019), .ZN(N197)
         );
  MOAI22D1 U1433 ( .A1(net7019), .A2(n419), .B1(n688), .B2(net7017), .ZN(N160)
         );
  MOAI22D1 U1434 ( .A1(n335), .A2(net7021), .B1(n689), .B2(net7015), .ZN(N211)
         );
  CKND0 U1435 ( .I(sa32_sr[4]), .ZN(n690) );
  XOR2D0 U1436 ( .A1(w0[11]), .A2(n646), .Z(N444) );
  MOAI22D1 U1437 ( .A1(n131), .A2(net7025), .B1(n671), .B2(net7021), .ZN(N83)
         );
  INVD1 U1438 ( .I(w3[5]), .ZN(n9) );
  XOR2D0 U1439 ( .A1(w1[20]), .A2(n633), .Z(N419) );
  MOAI22D1 U1440 ( .A1(n405), .A2(net7019), .B1(n692), .B2(net7013), .ZN(N165)
         );
  XNR2D1 U1441 ( .A1(text_in_r[69]), .A2(n37), .ZN(n692) );
  CKXOR2D0 U1442 ( .A1(w1[12]), .A2(sa21_sr[4]), .Z(N451) );
  XOR4D0 U1443 ( .A1(n230), .A2(n229), .A3(sa00_sr[3]), .A4(n231), .Z(n228) );
  XOR2D0 U1444 ( .A1(w1[3]), .A2(n538), .Z(N484) );
  MOAI22D1 U1445 ( .A1(n488), .A2(net7017), .B1(n693), .B2(net7011), .ZN(N116)
         );
  CKND0 U1446 ( .I(n84), .ZN(n694) );
  XOR2D0 U1447 ( .A1(w0[28]), .A2(n622), .Z(N379) );
  CKXOR2D0 U1448 ( .A1(w0[23]), .A2(sa10_sr[7]), .Z(N408) );
  XOR2D0 U1449 ( .A1(n34), .A2(sa01_sr[2]), .Z(n695) );
  INVD1 U1450 ( .I(w1[2]), .ZN(n34) );
  MOAI22D1 U1451 ( .A1(n126), .A2(net7025), .B1(n696), .B2(net7017), .ZN(N84)
         );
  CKXOR2D1 U1452 ( .A1(sa22_sr[4]), .A2(sa12_sr[4]), .Z(n439) );
  MOAI22D1 U1453 ( .A1(n396), .A2(net7019), .B1(n697), .B2(net7013), .ZN(N177)
         );
  XOR2D0 U1454 ( .A1(w2[3]), .A2(n549), .Z(N492) );
  XOR2D0 U1455 ( .A1(w2[17]), .A2(n639), .Z(N430) );
  MOAI22D1 U1456 ( .A1(n497), .A2(net7017), .B1(n698), .B2(net7023), .ZN(N113)
         );
  XOR2D0 U1457 ( .A1(w1[28]), .A2(n626), .Z(N387) );
  MOAI22D1 U1458 ( .A1(n253), .A2(net7023), .B1(n699), .B2(net7021), .ZN(N261)
         );
  XNR2D0 U1459 ( .A1(text_in_r[21]), .A2(w3[21]), .ZN(n150) );
  MOAI22D1 U1460 ( .A1(n330), .A2(net7021), .B1(n700), .B2(net7013), .ZN(N212)
         );
  XOR2D0 U1461 ( .A1(w2[7]), .A2(sa32_sr[7]), .Z(N488) );
  MOAI22D1 U1462 ( .A1(n228), .A2(net7023), .B1(n701), .B2(net7021), .ZN(N276)
         );
  CKXOR2D0 U1463 ( .A1(w3[28]), .A2(n558), .Z(N403) );
  MOAI22D1 U1464 ( .A1(n448), .A2(net7019), .B1(n702), .B2(net7011), .ZN(N145)
         );
  CKXOR2D0 U1465 ( .A1(w1[23]), .A2(sa11_sr[7]), .Z(N416) );
  XOR2D0 U1466 ( .A1(w1[9]), .A2(n524), .Z(N454) );
  CKXOR2D0 U1467 ( .A1(w3[4]), .A2(n532), .Z(N499) );
  MOAI22D1 U1468 ( .A1(n209), .A2(net7023), .B1(n703), .B2(net7019), .ZN(N34)
         );
  XNR2D1 U1469 ( .A1(text_in_r[2]), .A2(n6), .ZN(n703) );
  MOAI22D1 U1470 ( .A1(n233), .A2(net7023), .B1(n704), .B2(net7015), .ZN(N275)
         );
  MOAI22D1 U1471 ( .A1(net7021), .A2(n311), .B1(n705), .B2(net7025), .ZN(N226)
         );
  XNR2D1 U1472 ( .A1(text_in_r[98]), .A2(n56), .ZN(n705) );
  OAI22D1 U1473 ( .A1(n338), .A2(net7001), .B1(net7021), .B2(n339), .ZN(N210)
         );
  CKXOR2D0 U1474 ( .A1(w0[15]), .A2(sa20_sr[7]), .Z(N440) );
  XNR2D0 U1475 ( .A1(text_in_r[31]), .A2(w3[31]), .ZN(n113) );
  XNR3D0 U1476 ( .A1(w3[31]), .A2(sa13_sr[6]), .A3(sa13_sr[7]), .ZN(n116) );
  CKXOR2D0 U1477 ( .A1(w2[28]), .A2(n564), .Z(N395) );
  CKXOR2D0 U1478 ( .A1(w3[9]), .A2(n610), .Z(N470) );
  MOAI22D1 U1479 ( .A1(net7017), .A2(n472), .B1(n706), .B2(net7011), .ZN(N130)
         );
  XNR2D1 U1480 ( .A1(text_in_r[50]), .A2(n22), .ZN(n706) );
  CKXOR2D0 U1481 ( .A1(w3[17]), .A2(sa13_sr[1]), .Z(N438) );
  XNR2D0 U1482 ( .A1(text_in_r[13]), .A2(w3[13]), .ZN(n178) );
  CKND0 U1483 ( .I(sa12_sr[4]), .ZN(n90) );
  MOAI22D1 U1484 ( .A1(n460), .A2(net7017), .B1(n707), .B2(net7023), .ZN(N133)
         );
  XNR2D1 U1485 ( .A1(text_in_r[53]), .A2(n25), .ZN(n707) );
  XNR2D0 U1486 ( .A1(text_in_r[10]), .A2(w3[10]), .ZN(n187) );
  MOAI22D1 U1487 ( .A1(net7021), .A2(n344), .B1(n708), .B2(net7031), .ZN(N209)
         );
  CKXOR2D0 U1488 ( .A1(w2[20]), .A2(n602), .Z(N427) );
  XOR2D0 U1489 ( .A1(w2[11]), .A2(sa22_sr[3]), .Z(N460) );
  XOR3D1 U1490 ( .A1(sa22_sr[3]), .A2(w2[19]), .A3(n104), .Z(n470) );
  CKXOR2D0 U1491 ( .A1(w3[12]), .A2(n540), .Z(N467) );
  XOR3D1 U1492 ( .A1(w0[20]), .A2(n624), .A3(n234), .Z(n259) );
  XOR2D0 U1493 ( .A1(w0[4]), .A2(sa30_sr[4]), .Z(N475) );
  CKXOR2D0 U1494 ( .A1(w0[20]), .A2(n680), .Z(N411) );
  MOAI22D1 U1495 ( .A1(n416), .A2(net7019), .B1(n709), .B2(net7033), .ZN(N161)
         );
  CKXOR2D0 U1496 ( .A1(w0[1]), .A2(n596), .Z(N478) );
  CKXOR2D0 U1497 ( .A1(w0[17]), .A2(n694), .Z(N414) );
  XOR3D1 U1498 ( .A1(sa21_sr[4]), .A2(w1[20]), .A3(n336), .Z(n362) );
  XNR2D0 U1499 ( .A1(text_in_r[30]), .A2(w3[30]), .ZN(n117) );
  XNR3D0 U1500 ( .A1(w3[30]), .A2(sa33_sr[6]), .A3(sa13_sr[5]), .ZN(n120) );
  XNR3D0 U1501 ( .A1(w3[29]), .A2(sa33_sr[5]), .A3(n568), .ZN(n124) );
  CKXOR2D0 U1502 ( .A1(w3[20]), .A2(n609), .Z(N435) );
  CKXOR2D0 U1503 ( .A1(w2[9]), .A2(n614), .Z(N462) );
  CKXOR2D0 U1504 ( .A1(w3[25]), .A2(n545), .Z(N406) );
  CKXOR2D0 U1505 ( .A1(w1[25]), .A2(sa01_sr[1]), .Z(N390) );
  XOR2D0 U1506 ( .A1(w1[4]), .A2(sa31_sr[4]), .Z(N483) );
  CKXOR2D0 U1507 ( .A1(w0[9]), .A2(sa20_sr[1]), .Z(N446) );
  XOR2D0 U1508 ( .A1(w1[1]), .A2(sa31_sr[1]), .Z(N486) );
  XOR2D0 U1509 ( .A1(w2[1]), .A2(n515), .Z(N494) );
  XNR3D0 U1510 ( .A1(n608), .A2(n104), .A3(n446), .ZN(n445) );
endmodule


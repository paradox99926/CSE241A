/*
###############################################################
#  Design:            usb_phy
###############################################################
*/
module usb_phy (
	clk, 
	rst, 
	phy_tx_mode, 
	usb_rst, 
	txdp, 
	txdn, 
	txoe, 
	rxd, 
	rxdp, 
	rxdn, 
	DataOut_i, 
	TxValid_i, 
	TxReady_o, 
	RxValid_o, 
	RxActive_o, 
	RxError_o, 
	DataIn_o, 
	LineState_o);
   input clk;
   input rst;
   input phy_tx_mode;
   output usb_rst;
   output txdp;
   output txdn;
   output txoe;
   input rxd;
   input rxdp;
   input rxdn;
   input [7:0] DataOut_i;
   input TxValid_i;
   output TxReady_o;
   output RxValid_o;
   output RxActive_o;
   output RxError_o;
   output [7:0] DataIn_o;
   output [1:0] LineState_o;

   // Internal wires
   wire FE_OFN1_fs_ce;
   wire FE_DBTN0_i_tx_phy_state_1_;
   wire fs_ce;
   wire N26;
   wire i_tx_phy_txoe_r2;
   wire i_tx_phy_append_eop_sync4;
   wire i_tx_phy_append_eop_sync3;
   wire i_tx_phy_append_eop_sync1;
   wire i_tx_phy_append_eop;
   wire i_tx_phy_append_eop_sync2;
   wire i_tx_phy_txoe_r1;
   wire i_tx_phy_sd_nrzi_o;
   wire i_tx_phy_sd_bs_o;
   wire i_tx_phy_sft_done_r;
   wire i_tx_phy_sft_done;
   wire i_tx_phy_N88;
   wire i_tx_phy_N87;
   wire i_tx_phy_sd_raw_o;
   wire i_tx_phy_data_done;
   wire i_tx_phy_tx_ip_sync;
   wire i_tx_phy_tx_ip;
   wire i_tx_phy_ld_data;
   wire i_tx_phy_N18;
   wire i_rx_phy_N166;
   wire i_rx_phy_se0_r;
   wire i_rx_phy_N165;
   wire i_rx_phy_rx_valid1;
   wire i_rx_phy_N136;
   wire i_rx_phy_shift_en;
   wire i_rx_phy_sd_nrzi;
   wire i_rx_phy_sd_r;
   wire i_rx_phy_rx_valid_r;
   wire i_rx_phy_fs_ce_r2;
   wire i_rx_phy_fs_ce_r1;
   wire i_rx_phy_fs_ce_d;
   wire i_rx_phy_N32;
   wire i_rx_phy_N31;
   wire i_rx_phy_rxd_r;
   wire i_rx_phy_se0_s;
   wire i_rx_phy_rxdn_s;
   wire i_rx_phy_N29;
   wire i_rx_phy_rxdn_s_r;
   wire i_rx_phy_N28;
   wire i_rx_phy_rxdn_s0;
   wire i_rx_phy_rxdp_s;
   wire i_rx_phy_N27;
   wire i_rx_phy_rxdp_s_r;
   wire i_rx_phy_N26;
   wire i_rx_phy_rxdp_s0;
   wire i_rx_phy_rxd_s;
   wire i_rx_phy_rxd_s1;
   wire i_rx_phy_rxd_s0;
   wire i_rx_phy_N20;
   wire i_rx_phy_rx_en;
   wire i_rx_phy_byte_err;
   wire i_rx_phy_bit_stuff_err;
   wire i_rx_phy_sync_err;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire [4:0] rst_cnt;
   wire [2:0] i_tx_phy_state;
   wire [2:0] i_tx_phy_one_cnt;
   wire [7:0] i_tx_phy_hold_reg;
   wire [7:0] i_tx_phy_hold_reg_d;
   wire [2:0] i_tx_phy_bit_cnt;
   wire [2:0] i_rx_phy_bit_cnt;
   wire [2:0] i_rx_phy_one_cnt;
   wire [2:0] i_rx_phy_fs_state;
   wire [1:0] i_rx_phy_dpll_state;

   in01f04 FE_OFC1_fs_ce (.o(FE_OFN1_fs_ce),
	.a(fs_ce));
   in01f03 FE_DBTC0_i_tx_phy_state_1_ (.o(FE_DBTN0_i_tx_phy_state_1_),
	.a(i_tx_phy_state[1]));
   ms00f80 i_rx_phy_rxdn_s0_reg (.o(i_rx_phy_rxdn_s0),
	.ck(clk),
	.d(rxdn));
   ms00f80 i_rx_phy_rxdn_s1_reg (.o(LineState_o[1]),
	.ck(clk),
	.d(i_rx_phy_rxdn_s0));
   ms00f80 i_rx_phy_rxdn_s_r_reg (.o(i_rx_phy_rxdn_s_r),
	.ck(clk),
	.d(i_rx_phy_N28));
   ms00f80 i_rx_phy_rxdn_s_reg (.o(i_rx_phy_rxdn_s),
	.ck(clk),
	.d(i_rx_phy_N29));
   ms00f80 i_rx_phy_rxdp_s0_reg (.o(i_rx_phy_rxdp_s0),
	.ck(clk),
	.d(rxdp));
   ms00f80 i_rx_phy_rxdp_s1_reg (.o(LineState_o[0]),
	.ck(clk),
	.d(i_rx_phy_rxdp_s0));
   ms00f80 i_rx_phy_rxdp_s_r_reg (.o(i_rx_phy_rxdp_s_r),
	.ck(clk),
	.d(i_rx_phy_N26));
   ms00f80 i_rx_phy_rxdp_s_reg (.o(i_rx_phy_rxdp_s),
	.ck(clk),
	.d(i_rx_phy_N27));
   ms00f80 i_rx_phy_se0_r_reg (.o(i_rx_phy_se0_r),
	.ck(clk),
	.d(n592));
   ms00f80 i_rx_phy_rxd_s0_reg (.o(i_rx_phy_rxd_s0),
	.ck(clk),
	.d(rxd));
   ms00f80 i_rx_phy_rxd_s1_reg (.o(i_rx_phy_rxd_s1),
	.ck(clk),
	.d(i_rx_phy_rxd_s0));
   ms00f80 i_rx_phy_rxd_s_reg (.o(i_rx_phy_rxd_s),
	.ck(clk),
	.d(n147));
   ms00f80 i_rx_phy_rxd_r_reg (.o(i_rx_phy_rxd_r),
	.ck(clk),
	.d(i_rx_phy_rxd_s));
   ms00f80 i_rx_phy_rx_en_reg (.o(i_rx_phy_rx_en),
	.ck(clk),
	.d(txoe));
   ms00f80 i_rx_phy_dpll_state_reg_1_ (.o(i_rx_phy_dpll_state[1]),
	.ck(clk),
	.d(i_rx_phy_N32));
   ms00f80 i_rx_phy_fs_ce_r1_reg (.o(i_rx_phy_fs_ce_r1),
	.ck(clk),
	.d(i_rx_phy_fs_ce_d));
   ms00f80 i_rx_phy_fs_ce_r2_reg (.o(i_rx_phy_fs_ce_r2),
	.ck(clk),
	.d(i_rx_phy_fs_ce_r1));
   ms00f80 i_rx_phy_fs_ce_reg (.o(fs_ce),
	.ck(clk),
	.d(i_rx_phy_fs_ce_r2));
   ms00f80 i_rx_phy_sd_r_reg (.o(i_rx_phy_sd_r),
	.ck(clk),
	.d(n146));
   ms00f80 i_rx_phy_se0_s_reg (.o(i_rx_phy_se0_s),
	.ck(clk),
	.d(n145));
   ms00f80 rst_cnt_reg_0_ (.o(rst_cnt[0]),
	.ck(clk),
	.d(n144));
   ms00f80 rst_cnt_reg_4_ (.o(rst_cnt[4]),
	.ck(clk),
	.d(n143));
   ms00f80 rst_cnt_reg_3_ (.o(rst_cnt[3]),
	.ck(clk),
	.d(n142));
   ms00f80 rst_cnt_reg_2_ (.o(rst_cnt[2]),
	.ck(clk),
	.d(n141));
   ms00f80 rst_cnt_reg_1_ (.o(rst_cnt[1]),
	.ck(clk),
	.d(n140));
   ms00f80 usb_rst_reg (.o(usb_rst),
	.ck(clk),
	.d(N26));
   ms00f80 i_tx_phy_append_eop_sync1_reg (.o(i_tx_phy_append_eop_sync1),
	.ck(clk),
	.d(n139));
   ms00f80 i_tx_phy_append_eop_sync2_reg (.o(i_tx_phy_append_eop_sync2),
	.ck(clk),
	.d(n138));
   ms00f80 i_tx_phy_append_eop_sync3_reg (.o(i_tx_phy_append_eop_sync3),
	.ck(clk),
	.d(n137));
   ms00f80 i_tx_phy_append_eop_sync4_reg (.o(i_tx_phy_append_eop_sync4),
	.ck(clk),
	.d(n136));
   ms00f80 i_tx_phy_tx_ip_reg (.o(i_tx_phy_tx_ip),
	.ck(clk),
	.d(n135));
   ms00f80 i_tx_phy_tx_ip_sync_reg (.o(i_tx_phy_tx_ip_sync),
	.ck(clk),
	.d(n134));
   ms00f80 i_tx_phy_txoe_r1_reg (.o(i_tx_phy_txoe_r1),
	.ck(clk),
	.d(n133));
   ms00f80 i_tx_phy_txoe_r2_reg (.o(i_tx_phy_txoe_r2),
	.ck(clk),
	.d(n132));
   ms00f80 i_tx_phy_txoe_reg (.o(txoe),
	.ck(clk),
	.d(n131));
   ms00f80 i_tx_phy_data_done_reg (.o(i_tx_phy_data_done),
	.ck(clk),
	.d(n130));
   ms00f80 i_tx_phy_state_reg_0_ (.o(i_tx_phy_state[0]),
	.ck(clk),
	.d(n129));
   ms00f80 i_tx_phy_state_reg_2_ (.o(i_tx_phy_state[2]),
	.ck(clk),
	.d(n128));
   ms00f80 i_tx_phy_state_reg_1_ (.o(i_tx_phy_state[1]),
	.ck(clk),
	.d(n127));
   ms00f80 i_tx_phy_ld_data_reg (.o(i_tx_phy_ld_data),
	.ck(clk),
	.d(n591));
   ms00f80 i_tx_phy_hold_reg_reg_7_ (.o(i_tx_phy_hold_reg[7]),
	.ck(clk),
	.d(n126));
   ms00f80 i_tx_phy_hold_reg_d_reg_7_ (.o(i_tx_phy_hold_reg_d[7]),
	.ck(clk),
	.d(i_tx_phy_hold_reg[7]));
   ms00f80 i_tx_phy_hold_reg_reg_6_ (.o(i_tx_phy_hold_reg[6]),
	.ck(clk),
	.d(n125));
   ms00f80 i_tx_phy_hold_reg_d_reg_6_ (.o(i_tx_phy_hold_reg_d[6]),
	.ck(clk),
	.d(i_tx_phy_hold_reg[6]));
   ms00f80 i_tx_phy_hold_reg_reg_5_ (.o(i_tx_phy_hold_reg[5]),
	.ck(clk),
	.d(n124));
   ms00f80 i_tx_phy_hold_reg_d_reg_5_ (.o(i_tx_phy_hold_reg_d[5]),
	.ck(clk),
	.d(i_tx_phy_hold_reg[5]));
   ms00f80 i_tx_phy_hold_reg_reg_4_ (.o(i_tx_phy_hold_reg[4]),
	.ck(clk),
	.d(n123));
   ms00f80 i_tx_phy_hold_reg_d_reg_4_ (.o(i_tx_phy_hold_reg_d[4]),
	.ck(clk),
	.d(i_tx_phy_hold_reg[4]));
   ms00f80 i_tx_phy_hold_reg_reg_3_ (.o(i_tx_phy_hold_reg[3]),
	.ck(clk),
	.d(n122));
   ms00f80 i_tx_phy_hold_reg_d_reg_3_ (.o(i_tx_phy_hold_reg_d[3]),
	.ck(clk),
	.d(i_tx_phy_hold_reg[3]));
   ms00f80 i_tx_phy_hold_reg_reg_2_ (.o(i_tx_phy_hold_reg[2]),
	.ck(clk),
	.d(n121));
   ms00f80 i_tx_phy_hold_reg_d_reg_2_ (.o(i_tx_phy_hold_reg_d[2]),
	.ck(clk),
	.d(i_tx_phy_hold_reg[2]));
   ms00f80 i_tx_phy_hold_reg_reg_1_ (.o(i_tx_phy_hold_reg[1]),
	.ck(clk),
	.d(n120));
   ms00f80 i_tx_phy_hold_reg_d_reg_1_ (.o(i_tx_phy_hold_reg_d[1]),
	.ck(clk),
	.d(i_tx_phy_hold_reg[1]));
   ms00f80 i_tx_phy_hold_reg_reg_0_ (.o(i_tx_phy_hold_reg[0]),
	.ck(clk),
	.d(n119));
   ms00f80 i_tx_phy_hold_reg_d_reg_0_ (.o(i_tx_phy_hold_reg_d[0]),
	.ck(clk),
	.d(i_tx_phy_hold_reg[0]));
   ms00f80 i_tx_phy_sd_raw_o_reg (.o(i_tx_phy_sd_raw_o),
	.ck(clk),
	.d(i_tx_phy_N87));
   ms00f80 i_tx_phy_one_cnt_reg_0_ (.o(i_tx_phy_one_cnt[0]),
	.ck(clk),
	.d(n118));
   ms00f80 i_tx_phy_one_cnt_reg_1_ (.o(i_tx_phy_one_cnt[1]),
	.ck(clk),
	.d(n117));
   ms00f80 i_tx_phy_one_cnt_reg_2_ (.o(i_tx_phy_one_cnt[2]),
	.ck(clk),
	.d(n116));
   ms00f80 i_tx_phy_bit_cnt_reg_0_ (.o(i_tx_phy_bit_cnt[0]),
	.ck(clk),
	.d(n115));
   ms00f80 i_tx_phy_bit_cnt_reg_1_ (.o(i_tx_phy_bit_cnt[1]),
	.ck(clk),
	.d(n114));
   ms00f80 i_tx_phy_bit_cnt_reg_2_ (.o(i_tx_phy_bit_cnt[2]),
	.ck(clk),
	.d(n113));
   ms00f80 i_tx_phy_sft_done_r_reg (.o(i_tx_phy_sft_done_r),
	.ck(clk),
	.d(i_tx_phy_sft_done));
   ms00f80 i_tx_phy_TxReady_o_reg (.o(TxReady_o),
	.ck(clk),
	.d(i_tx_phy_N18));
   ms00f80 i_tx_phy_append_eop_reg (.o(i_tx_phy_append_eop),
	.ck(clk),
	.d(n112));
   ms00f80 i_tx_phy_sd_bs_o_reg (.o(i_tx_phy_sd_bs_o),
	.ck(clk),
	.d(n111));
   ms00f80 i_tx_phy_sd_nrzi_o_reg (.o(i_tx_phy_sd_nrzi_o),
	.ck(clk),
	.d(n110));
   ms00f80 i_tx_phy_txdn_reg (.o(txdn),
	.ck(clk),
	.d(n109));
   ms00f80 i_tx_phy_txdp_reg (.o(txdp),
	.ck(clk),
	.d(n108));
   ms00f80 i_rx_phy_dpll_state_reg_0_ (.o(i_rx_phy_dpll_state[0]),
	.ck(clk),
	.d(i_rx_phy_N31));
   ms00f80 i_rx_phy_fs_state_reg_0_ (.o(i_rx_phy_fs_state[0]),
	.ck(clk),
	.d(n107));
   ms00f80 i_rx_phy_fs_state_reg_2_ (.o(i_rx_phy_fs_state[2]),
	.ck(clk),
	.d(n106));
   ms00f80 i_rx_phy_fs_state_reg_1_ (.o(i_rx_phy_fs_state[1]),
	.ck(clk),
	.d(n105));
   ms00f80 i_rx_phy_rx_active_reg (.o(RxActive_o),
	.ck(clk),
	.d(n104));
   ms00f80 i_rx_phy_shift_en_reg (.o(i_rx_phy_shift_en),
	.ck(clk),
	.d(n103));
   ms00f80 i_rx_phy_sd_nrzi_reg (.o(i_rx_phy_sd_nrzi),
	.ck(clk),
	.d(n102));
   ms00f80 i_rx_phy_one_cnt_reg_0_ (.o(i_rx_phy_one_cnt[0]),
	.ck(clk),
	.d(n101));
   ms00f80 i_rx_phy_one_cnt_reg_1_ (.o(i_rx_phy_one_cnt[1]),
	.ck(clk),
	.d(n100));
   ms00f80 i_rx_phy_one_cnt_reg_2_ (.o(i_rx_phy_one_cnt[2]),
	.ck(clk),
	.d(n99));
   ms00f80 i_rx_phy_bit_stuff_err_reg (.o(i_rx_phy_bit_stuff_err),
	.ck(clk),
	.d(i_rx_phy_N136));
   ms00f80 i_rx_phy_hold_reg_reg_7_ (.o(DataIn_o[7]),
	.ck(clk),
	.d(n98));
   ms00f80 i_rx_phy_hold_reg_reg_6_ (.o(DataIn_o[6]),
	.ck(clk),
	.d(n97));
   ms00f80 i_rx_phy_hold_reg_reg_5_ (.o(DataIn_o[5]),
	.ck(clk),
	.d(n96));
   ms00f80 i_rx_phy_hold_reg_reg_4_ (.o(DataIn_o[4]),
	.ck(clk),
	.d(n95));
   ms00f80 i_rx_phy_hold_reg_reg_3_ (.o(DataIn_o[3]),
	.ck(clk),
	.d(n94));
   ms00f80 i_rx_phy_hold_reg_reg_2_ (.o(DataIn_o[2]),
	.ck(clk),
	.d(n93));
   ms00f80 i_rx_phy_hold_reg_reg_1_ (.o(DataIn_o[1]),
	.ck(clk),
	.d(n92));
   ms00f80 i_rx_phy_hold_reg_reg_0_ (.o(DataIn_o[0]),
	.ck(clk),
	.d(n91));
   ms00f80 i_rx_phy_bit_cnt_reg_0_ (.o(i_rx_phy_bit_cnt[0]),
	.ck(clk),
	.d(n90));
   ms00f80 i_rx_phy_bit_cnt_reg_1_ (.o(i_rx_phy_bit_cnt[1]),
	.ck(clk),
	.d(n89));
   ms00f80 i_rx_phy_bit_cnt_reg_2_ (.o(i_rx_phy_bit_cnt[2]),
	.ck(clk),
	.d(n88));
   ms00f80 i_rx_phy_byte_err_reg (.o(i_rx_phy_byte_err),
	.ck(clk),
	.d(i_rx_phy_N166));
   ms00f80 i_rx_phy_rx_valid1_reg (.o(i_rx_phy_rx_valid1),
	.ck(clk),
	.d(n87));
   ms00f80 i_rx_phy_rx_valid_reg (.o(RxValid_o),
	.ck(clk),
	.d(i_rx_phy_N165));
   ms00f80 i_rx_phy_rx_valid_r_reg (.o(i_rx_phy_rx_valid_r),
	.ck(clk),
	.d(n86));
   ms00f80 i_rx_phy_sync_err_reg (.o(i_rx_phy_sync_err),
	.ck(clk),
	.d(i_rx_phy_N20));
   ms00f80 i_tx_phy_sft_done_reg (.o(i_tx_phy_sft_done),
	.ck(clk),
	.d(i_tx_phy_N88));
   no02m02 U407 (.o(i_rx_phy_N20),
	.a(n439),
	.b(n438));
   na02m01 U408 (.o(n538),
	.a(i_rx_phy_sd_nrzi),
	.b(n562));
   ao12f01 U409 (.o(n493),
	.a(n496),
	.b(n489),
	.c(n488));
   na03m01 U410 (.o(n380),
	.a(i_rx_phy_bit_cnt[0]),
	.b(n379),
	.c(n548));
   na03m02 U411 (.o(n457),
	.a(i_rx_phy_bit_cnt[1]),
	.b(rst),
	.c(n480));
   ao22f01 U412 (.o(n570),
	.a(n569),
	.b(rst_cnt[3]),
	.c(n568),
	.d(n567));
   no02m02 U413 (.o(n523),
	.a(n517),
	.b(n524));
   no02f02 U414 (.o(n558),
	.a(n551),
	.b(n550));
   no02m02 U415 (.o(n578),
	.a(n581),
	.b(i_tx_phy_one_cnt[0]));
   na02m01 U416 (.o(n508),
	.a(n510),
	.b(n529));
   na02m03 U417 (.o(n581),
	.a(n524),
	.b(i_tx_phy_sd_raw_o));
   ao12f02 U418 (.o(n573),
	.a(n435),
	.b(n370),
	.c(n369));
   in01m02 U419 (.o(n520),
	.a(i_tx_phy_bit_cnt[1]));
   na02f01 U420 (.o(n370),
	.a(n416),
	.b(i_rx_phy_rxd_r));
   no02m02 U421 (.o(n423),
	.a(FE_DBTN0_i_tx_phy_state_1_),
	.b(i_tx_phy_state[0]));
   no04f04 U422 (.o(n443),
	.a(FE_OFN1_fs_ce),
	.b(n592),
	.c(RxActive_o),
	.d(i_rx_phy_se0_s));
   na02f02 U423 (.o(n477),
	.a(n424),
	.b(n339));
   no02f04 U424 (.o(n592),
	.a(i_rx_phy_rxdp_s),
	.b(i_rx_phy_rxdn_s));
   no04f06 U425 (.o(n529),
	.a(n590),
	.b(LineState_o[0]),
	.c(LineState_o[1]),
	.d(usb_rst));
   no02m02 U426 (.o(n410),
	.a(FE_DBTN0_i_tx_phy_state_1_),
	.b(n426));
   na02m01 U427 (.o(n531),
	.a(rst_cnt[0]),
	.b(rst_cnt[1]));
   no03s02 U428 (.o(n366),
	.a(LineState_o[0]),
	.b(LineState_o[1]),
	.c(n583));
   na02m02 U429 (.o(n426),
	.a(n331),
	.b(i_tx_phy_sft_done));
   na02m02 U430 (.o(n378),
	.a(rst),
	.b(i_rx_phy_shift_en));
   na02m02 U431 (.o(n326),
	.a(i_tx_phy_state[2]),
	.b(n327));
   in01s06 U432 (.o(n583),
	.a(rst));
   in01s02 U433 (.o(n331),
	.a(i_tx_phy_sft_done_r));
   na02m02 U434 (.o(n513),
	.a(i_tx_phy_bit_cnt[2]),
	.b(i_tx_phy_bit_cnt[0]));
   no04f02 U435 (.o(n547),
	.a(n548),
	.b(n546),
	.c(n545),
	.d(n544));
   oa12f02 U436 (.o(n579),
	.a(i_tx_phy_one_cnt[1]),
	.b(n578),
	.c(n577));
   na02f08 U437 (.o(n590),
	.a(rst),
	.b(fs_ce));
   no02s02 U438 (.o(n500),
	.a(n485),
	.b(n484));
   in01m02 U439 (.o(n562),
	.a(n537));
   ao12f02 U440 (.o(n533),
	.a(n527),
	.b(n529),
	.c(n528));
   na02f02 U441 (.o(n527),
	.a(n509),
	.b(n508));
   no02f01 U442 (.o(n567),
	.a(n531),
	.b(n530));
   no02f04 U443 (.o(n456),
	.a(FE_OFN1_fs_ce),
	.b(n408));
   no02m02 U444 (.o(n386),
	.a(n367),
	.b(n529));
   in01f01 U445 (.o(n548),
	.a(n456));
   in01m01 U446 (.o(n569),
	.a(n564));
   oa12m02 U447 (.o(n496),
	.a(n441),
	.b(n583),
	.c(n443));
   ao12f02 U448 (.o(n564),
	.a(n386),
	.b(n529),
	.c(n387));
   in01m01 U449 (.o(n509),
	.a(n386));
   in01f02 U450 (.o(n550),
	.a(n477));
   na03m02 U451 (.o(n441),
	.a(n488),
	.b(n440),
	.c(n497));
   no03f03 U452 (.o(n471),
	.a(i_tx_phy_one_cnt[0]),
	.b(n576),
	.c(n476));
   oa22m01 U453 (.o(n100),
	.a(n470),
	.b(n464),
	.c(n466),
	.d(n467));
   oa22m01 U454 (.o(n99),
	.a(n470),
	.b(n469),
	.c(n468),
	.d(n467));
   no02s02 U455 (.o(n129),
	.a(n583),
	.b(n344));
   ao12f02 U456 (.o(n467),
	.a(n463),
	.b(n585),
	.c(i_rx_phy_shift_en));
   oa12f01 U457 (.o(n127),
	.a(n350),
	.b(n352),
	.c(FE_DBTN0_i_tx_phy_state_1_));
   no02f03 U458 (.o(n524),
	.a(n472),
	.b(n471));
   na02f02 U459 (.o(n472),
	.a(i_tx_phy_tx_ip_sync),
	.b(n505));
   oa22f01 U460 (.o(n103),
	.a(n503),
	.b(fs_ce),
	.c(FE_OFN1_fs_ce),
	.d(n501));
   ao12f01 U461 (.o(n501),
	.a(RxActive_o),
	.b(n500),
	.c(n499));
   na02f03 U462 (.o(n537),
	.a(i_rx_phy_shift_en),
	.b(n456));
   no02f01 U463 (.o(n488),
	.a(n583),
	.b(i_rx_phy_fs_state[0]));
   in01f01 U465 (.o(n333),
	.a(n326));
   in01f02 U466 (.o(n327),
	.a(i_tx_phy_append_eop_sync3));
   na03m02 U468 (.o(n481),
	.a(i_rx_phy_bit_cnt[2]),
	.b(rst),
	.c(n480));
   na02s02 U469 (.o(n572),
	.a(n571),
	.b(n573));
   oa22f01 U470 (.o(n141),
	.a(n566),
	.b(n533),
	.c(n532),
	.d(rst_cnt[2]));
   oa12m02 U471 (.o(n338),
	.a(i_tx_phy_state[2]),
	.b(FE_OFN1_fs_ce),
	.c(i_tx_phy_append_eop_sync3));
   ao22f02 U472 (.o(n344),
	.a(n352),
	.b(n345),
	.c(i_tx_phy_state[0]),
	.d(n343));
   oa12m01 U473 (.o(n98),
	.a(n538),
	.b(n539),
	.c(n562));
   oa12m01 U474 (.o(n96),
	.a(n542),
	.b(n543),
	.c(n562));
   na02f01 U475 (.o(n542),
	.a(n562),
	.b(DataIn_o[6]));
   oa12m01 U476 (.o(n94),
	.a(n561),
	.b(n563),
	.c(n562));
   na02f01 U477 (.o(n561),
	.a(n562),
	.b(DataIn_o[4]));
   oa12m01 U478 (.o(n92),
	.a(n540),
	.b(n541),
	.c(n562));
   na02f01 U479 (.o(n540),
	.a(n562),
	.b(DataIn_o[2]));
   no02m02 U480 (.o(n128),
	.a(n583),
	.b(n337));
   ao12f02 U481 (.o(n350),
	.a(n348),
	.b(n349),
	.c(n423));
   no04f02 U482 (.o(n348),
	.a(n347),
	.b(n346),
	.c(n345),
	.d(i_tx_phy_state[1]));
   no02f02 U483 (.o(n463),
	.a(n470),
	.b(i_rx_phy_one_cnt[0]));
   ao12f01 U484 (.o(n480),
	.a(n503),
	.b(i_rx_phy_bit_cnt[0]),
	.c(n456));
   in01f01 U485 (.o(n332),
	.a(n328));
   ao22f01 U486 (.o(n512),
	.a(n527),
	.b(rst_cnt[1]),
	.c(n511),
	.d(n529));
   in01f02 U487 (.o(n329),
	.a(i_tx_phy_state[2]));
   oa22f02 U489 (.o(n328),
	.a(i_tx_phy_append_eop_sync3),
	.b(FE_DBTN0_i_tx_phy_state_1_),
	.c(n329),
	.d(fs_ce));
   no02f02 U490 (.o(n424),
	.a(i_tx_phy_state[2]),
	.b(i_tx_phy_state[1]));
   oa12f02 U491 (.o(n334),
	.a(n332),
	.b(i_tx_phy_state[0]),
	.c(n333));
   ao12f02 U492 (.o(n342),
	.a(n334),
	.b(n424),
	.c(n426));
   na02s02 U493 (.o(n336),
	.a(n342),
	.b(i_tx_phy_state[0]));
   no03s02 U494 (.o(n335),
	.a(i_tx_phy_state[2]),
	.b(FE_DBTN0_i_tx_phy_state_1_),
	.c(n336));
   ao12f01 U495 (.o(n337),
	.a(n335),
	.b(i_tx_phy_state[2]),
	.c(n336));
   no02s01 U496 (.o(n411),
	.a(i_tx_phy_state[0]),
	.b(i_tx_phy_data_done));
   na03s02 U497 (.o(n340),
	.a(n410),
	.b(n411),
	.c(n338));
   in01f01 U498 (.o(n394),
	.a(TxValid_i));
   no02s02 U499 (.o(n339),
	.a(n394),
	.b(i_tx_phy_state[0]));
   na03f02 U500 (.o(n341),
	.a(rst),
	.b(n340),
	.c(n477));
   no02f02 U501 (.o(n346),
	.a(n341),
	.b(n342));
   in01s01 U502 (.o(n352),
	.a(n346));
   in01s01 U503 (.o(n345),
	.a(i_tx_phy_state[0]));
   in01s01 U504 (.o(n343),
	.a(n342));
   na02s01 U505 (.o(n347),
	.a(n329),
	.b(rst));
   in01s01 U506 (.o(n349),
	.a(n347));
   na02s01 U507 (.o(n517),
	.a(rst),
	.b(i_tx_phy_tx_ip_sync));
   in01s01 U508 (.o(n356),
	.a(n517));
   no02s01 U509 (.o(n354),
	.a(n590),
	.b(i_tx_phy_sd_bs_o));
   na02s01 U510 (.o(n353),
	.a(n354),
	.b(i_tx_phy_sd_nrzi_o));
   oa12s01 U511 (.o(n355),
	.a(n353),
	.b(i_tx_phy_sd_nrzi_o),
	.c(n354));
   na03m02 U512 (.o(n110),
	.a(n356),
	.b(i_tx_phy_txoe_r1),
	.c(n355));
   in01s01 U513 (.o(n358),
	.a(n592));
   in01s01 U514 (.o(n418),
	.a(RxActive_o));
   no02s01 U515 (.o(n357),
	.a(i_rx_phy_bit_cnt[1]),
	.b(i_rx_phy_bit_cnt[2]));
   no04s01 U516 (.o(i_rx_phy_N166),
	.a(n358),
	.b(i_rx_phy_se0_r),
	.c(n418),
	.d(n357));
   in01s01 U517 (.o(n574),
	.a(i_rx_phy_dpll_state[0]));
   no02s01 U518 (.o(i_rx_phy_fs_ce_d),
	.a(i_rx_phy_dpll_state[1]),
	.b(n574));
   in01s01 U519 (.o(n361),
	.a(i_rx_phy_rxd_s1));
   in01s01 U520 (.o(n360),
	.a(i_rx_phy_rxd_s0));
   oa12s01 U521 (.o(n359),
	.a(i_rx_phy_rxd_s),
	.b(i_rx_phy_rxd_s0),
	.c(i_rx_phy_rxd_s1));
   oa12s01 U522 (.o(n147),
	.a(n359),
	.b(n361),
	.c(n360));
   na02s01 U523 (.o(n362),
	.a(LineState_o[1]),
	.b(i_rx_phy_rxdn_s0));
   in01s01 U524 (.o(i_rx_phy_N28),
	.a(n362));
   na02s01 U525 (.o(n363),
	.a(LineState_o[0]),
	.b(i_rx_phy_rxdp_s0));
   in01s01 U526 (.o(i_rx_phy_N26),
	.a(n363));
   in01s01 U527 (.o(n416),
	.a(i_rx_phy_rxd_s));
   in01s01 U528 (.o(n417),
	.a(i_rx_phy_sd_r));
   oa22s01 U529 (.o(n146),
	.a(n416),
	.b(FE_OFN1_fs_ce),
	.c(n417),
	.d(fs_ce));
   in01s01 U530 (.o(n365),
	.a(i_tx_phy_txoe_r1));
   in01s01 U531 (.o(n364),
	.a(i_tx_phy_txoe_r2));
   no02f04 U532 (.o(n585),
	.a(n583),
	.b(fs_ce));
   in01f02 U533 (.o(n588),
	.a(n585));
   oa22s01 U534 (.o(n132),
	.a(n590),
	.b(n365),
	.c(n364),
	.d(n588));
   in01f02 U535 (.o(n505),
	.a(n590));
   oa12s01 U536 (.o(n133),
	.a(n472),
	.b(n588),
	.c(n365));
   in01s01 U537 (.o(n367),
	.a(n366));
   in01s01 U538 (.o(n510),
	.a(rst_cnt[0]));
   oa12s01 U539 (.o(n144),
	.a(n508),
	.b(n509),
	.c(n510));
   in01s01 U540 (.o(n571),
	.a(i_rx_phy_fs_ce_d));
   na02s01 U541 (.o(n371),
	.a(n574),
	.b(i_rx_phy_dpll_state[1]));
   in01s01 U542 (.o(n368),
	.a(i_rx_phy_rxd_r));
   na02s01 U543 (.o(n369),
	.a(n368),
	.b(i_rx_phy_rxd_s));
   in01s01 U544 (.o(n435),
	.a(i_rx_phy_rx_en));
   no02s01 U545 (.o(n372),
	.a(n371),
	.b(n573));
   in01s01 U546 (.o(n373),
	.a(n372));
   ao12s01 U547 (.o(i_rx_phy_N32),
	.a(n583),
	.b(n571),
	.c(n373));
   no02s02 U548 (.o(n374),
	.a(n378),
	.b(FE_OFN1_fs_ce));
   in01s01 U549 (.o(n377),
	.a(n374));
   in01s02 U550 (.o(n375),
	.a(i_rx_phy_one_cnt[0]));
   na03f02 U551 (.o(n376),
	.a(n375),
	.b(i_rx_phy_one_cnt[2]),
	.c(i_rx_phy_one_cnt[1]));
   in01f02 U552 (.o(n408),
	.a(n376));
   no02f02 U553 (.o(n455),
	.a(n377),
	.b(n408));
   in01s01 U554 (.o(n483),
	.a(n455));
   in01s01 U555 (.o(n379),
	.a(n378));
   oa12s01 U556 (.o(n90),
	.a(n380),
	.b(n483),
	.c(i_rx_phy_bit_cnt[0]));
   in01s01 U557 (.o(n541),
	.a(DataIn_o[1]));
   na02s01 U558 (.o(n381),
	.a(n537),
	.b(DataIn_o[0]));
   oa12s01 U559 (.o(n91),
	.a(n381),
	.b(n537),
	.c(n541));
   in01s01 U560 (.o(n563),
	.a(DataIn_o[3]));
   na02s01 U561 (.o(n382),
	.a(n537),
	.b(DataIn_o[2]));
   oa12s01 U562 (.o(n93),
	.a(n382),
	.b(n537),
	.c(n563));
   in01s01 U563 (.o(n539),
	.a(DataIn_o[7]));
   na02s01 U564 (.o(n383),
	.a(n537),
	.b(DataIn_o[6]));
   oa12s01 U565 (.o(n97),
	.a(n383),
	.b(n537),
	.c(n539));
   in01s01 U566 (.o(n543),
	.a(DataIn_o[5]));
   na02s01 U567 (.o(n384),
	.a(n537),
	.b(DataIn_o[4]));
   oa12s01 U568 (.o(n95),
	.a(n384),
	.b(n537),
	.c(n543));
   in01s01 U569 (.o(n389),
	.a(rst_cnt[4]));
   na02s01 U570 (.o(n385),
	.a(rst_cnt[2]),
	.b(rst_cnt[3]));
   no02f02 U571 (.o(n565),
	.a(n385),
	.b(n531));
   in01s01 U572 (.o(n387),
	.a(n565));
   na03s01 U573 (.o(n388),
	.a(n565),
	.b(n529),
	.c(n389));
   oa12s01 U574 (.o(n143),
	.a(n388),
	.b(n389),
	.c(n564));
   no03s01 U575 (.o(n390),
	.a(i_rx_phy_sync_err),
	.b(i_rx_phy_byte_err),
	.c(i_rx_phy_bit_stuff_err));
   in01s01 U576 (.o(RxError_o),
	.a(n390));
   no02s01 U577 (.o(n391),
	.a(i_rx_phy_N28),
	.b(i_rx_phy_rxdn_s_r));
   in01s01 U578 (.o(i_rx_phy_N29),
	.a(n391));
   no02s01 U579 (.o(n392),
	.a(i_rx_phy_N26),
	.b(i_rx_phy_rxdp_s_r));
   in01s01 U580 (.o(i_rx_phy_N27),
	.a(n392));
   in01s01 U581 (.o(n393),
	.a(i_tx_phy_data_done));
   na02s01 U582 (.o(n395),
	.a(n393),
	.b(i_tx_phy_tx_ip));
   no02s01 U583 (.o(n427),
	.a(n394),
	.b(n583));
   na02s01 U584 (.o(n396),
	.a(n395),
	.b(n427));
   in01s01 U585 (.o(n130),
	.a(n396));
   ao12s01 U586 (.o(n397),
	.a(RxValid_o),
	.b(i_rx_phy_rx_valid_r),
	.c(FE_OFN1_fs_ce));
   in01s01 U587 (.o(n86),
	.a(n397));
   oa12s01 U588 (.o(n398),
	.a(fs_ce),
	.b(i_tx_phy_txoe_r1),
	.c(i_tx_phy_txoe_r2));
   oa12s01 U589 (.o(n399),
	.a(n398),
	.b(fs_ce),
	.c(txoe));
   na02s01 U590 (.o(n131),
	.a(n399),
	.b(rst));
   na02s01 U591 (.o(n400),
	.a(n565),
	.b(rst_cnt[4]));
   in01s01 U592 (.o(N26),
	.a(n400));
   in01s01 U593 (.o(n551),
	.a(i_tx_phy_ld_data));
   oa22s01 U594 (.o(n401),
	.a(n551),
	.b(DataOut_i[7]),
	.c(i_tx_phy_ld_data),
	.d(i_tx_phy_hold_reg[7]));
   na02s01 U595 (.o(n126),
	.a(n401),
	.b(n477));
   in01s01 U596 (.o(n402),
	.a(i_tx_phy_sd_nrzi_o));
   ao12s01 U597 (.o(n403),
	.a(n402),
	.b(phy_tx_mode),
	.c(i_tx_phy_append_eop_sync3));
   oa22s01 U598 (.o(n404),
	.a(FE_OFN1_fs_ce),
	.b(n403),
	.c(fs_ce),
	.d(txdp));
   na02s01 U599 (.o(n108),
	.a(n404),
	.b(rst));
   ao22s01 U600 (.o(n405),
	.a(FE_OFN1_fs_ce),
	.b(i_rx_phy_se0_s),
	.c(fs_ce),
	.d(n592));
   in01s01 U601 (.o(n145),
	.a(n405));
   na03s01 U602 (.o(n406),
	.a(fs_ce),
	.b(i_rx_phy_sd_nrzi),
	.c(RxActive_o));
   no02s01 U603 (.o(n407),
	.a(n406),
	.b(n592));
   na02s01 U604 (.o(n409),
	.a(n408),
	.b(n407));
   in01s01 U605 (.o(i_rx_phy_N136),
	.a(n409));
   in01s01 U606 (.o(n587),
	.a(i_tx_phy_append_eop_sync2));
   ao22s01 U607 (.o(n412),
	.a(n587),
	.b(i_tx_phy_append_eop),
	.c(n411),
	.d(n410));
   no02s01 U608 (.o(n112),
	.a(n583),
	.b(n412));
   ao22s01 U609 (.o(n413),
	.a(n585),
	.b(i_tx_phy_append_eop_sync1),
	.c(i_tx_phy_append_eop),
	.d(n505));
   in01s01 U610 (.o(n139),
	.a(n413));
   no02s01 U611 (.o(n515),
	.a(n520),
	.b(n513));
   in01s01 U612 (.o(n414),
	.a(n515));
   in01f01 U613 (.o(n576),
	.a(i_tx_phy_one_cnt[1]));
   in01f01 U614 (.o(n476),
	.a(i_tx_phy_one_cnt[2]));
   no02s01 U615 (.o(i_tx_phy_N88),
	.a(n414),
	.b(n471));
   na02s01 U616 (.o(n415),
	.a(n456),
	.b(i_rx_phy_rx_valid1));
   in01s01 U617 (.o(i_rx_phy_N165),
	.a(n415));
   oa12s01 U618 (.o(n421),
	.a(n505),
	.b(n416),
	.c(i_rx_phy_sd_r));
   no02s01 U619 (.o(n420),
	.a(n417),
	.b(i_rx_phy_rxd_s));
   ao22s01 U620 (.o(n419),
	.a(n418),
	.b(rst),
	.c(n585),
	.d(i_rx_phy_sd_nrzi));
   oa12s01 U621 (.o(n102),
	.a(n419),
	.b(n421),
	.c(n420));
   in01s01 U622 (.o(n422),
	.a(i_tx_phy_append_eop_sync1));
   oa22s01 U623 (.o(n138),
	.a(n422),
	.b(n590),
	.c(n587),
	.d(n588));
   ao22s01 U624 (.o(n425),
	.a(n424),
	.b(i_tx_phy_state[0]),
	.c(i_tx_phy_data_done),
	.d(n423));
   no02f01 U625 (.o(n591),
	.a(n426),
	.b(n425));
   na02s01 U626 (.o(n428),
	.a(n427),
	.b(n591));
   in01s01 U627 (.o(i_tx_phy_N18),
	.a(n428));
   na02f02 U628 (.o(n470),
	.a(n455),
	.b(i_rx_phy_sd_nrzi));
   na03s01 U629 (.o(n429),
	.a(i_rx_phy_shift_en),
	.b(n585),
	.c(i_rx_phy_one_cnt[0]));
   in01s01 U630 (.o(n430),
	.a(n429));
   no02s01 U631 (.o(n431),
	.a(n463),
	.b(n430));
   in01s01 U632 (.o(n101),
	.a(n431));
   no02s01 U633 (.o(n440),
	.a(i_rx_phy_fs_state[1]),
	.b(i_rx_phy_fs_state[2]));
   in01s01 U634 (.o(n433),
	.a(n440));
   in01s01 U635 (.o(n432),
	.a(i_rx_phy_rxdp_s));
   na02s02 U636 (.o(n497),
	.a(n432),
	.b(i_rx_phy_rx_en));
   na02f01 U637 (.o(n442),
	.a(n433),
	.b(n497));
   in01s01 U638 (.o(n437),
	.a(n442));
   in01s01 U639 (.o(n489),
	.a(n497));
   in01s01 U640 (.o(n434),
	.a(i_rx_phy_fs_state[0]));
   no03s02 U641 (.o(n492),
	.a(i_rx_phy_rxdn_s),
	.b(n435),
	.c(n434));
   ao12s01 U642 (.o(n436),
	.a(n492),
	.b(n489),
	.c(i_rx_phy_fs_state[2]));
   oa12f01 U643 (.o(n439),
	.a(n436),
	.b(i_rx_phy_fs_state[0]),
	.c(n437));
   na02s01 U644 (.o(n485),
	.a(i_rx_phy_fs_state[2]),
	.b(i_rx_phy_fs_state[0]));
   in01s01 U645 (.o(n498),
	.a(i_rx_phy_fs_state[1]));
   oa12s01 U646 (.o(n438),
	.a(n443),
	.b(n485),
	.c(n498));
   na02s01 U647 (.o(n445),
	.a(n442),
	.b(n488));
   in01f01 U648 (.o(n484),
	.a(n443));
   na03s01 U649 (.o(n444),
	.a(rst),
	.b(i_rx_phy_fs_state[0]),
	.c(n484));
   oa12s01 U650 (.o(n107),
	.a(n444),
	.b(n496),
	.c(n445));
   in01s01 U651 (.o(n446),
	.a(i_tx_phy_hold_reg_d[5]));
   no03s01 U652 (.o(n447),
	.a(i_tx_phy_bit_cnt[1]),
	.b(n513),
	.c(n446));
   ao12s01 U653 (.o(n454),
	.a(n447),
	.b(i_tx_phy_hold_reg_d[7]),
	.c(n515));
   oa22s01 U654 (.o(n449),
	.a(n520),
	.b(i_tx_phy_hold_reg_d[2]),
	.c(i_tx_phy_bit_cnt[1]),
	.d(i_tx_phy_hold_reg_d[0]));
   in01s01 U655 (.o(n516),
	.a(i_tx_phy_bit_cnt[2]));
   oa22s01 U656 (.o(n448),
	.a(n520),
	.b(i_tx_phy_hold_reg_d[6]),
	.c(i_tx_phy_bit_cnt[1]),
	.d(i_tx_phy_hold_reg_d[4]));
   ao22f01 U657 (.o(n452),
	.a(n449),
	.b(n516),
	.c(i_tx_phy_bit_cnt[2]),
	.d(n448));
   ao22s01 U658 (.o(n450),
	.a(n520),
	.b(i_tx_phy_hold_reg_d[1]),
	.c(i_tx_phy_bit_cnt[1]),
	.d(i_tx_phy_hold_reg_d[3]));
   oa12s01 U659 (.o(n451),
	.a(i_tx_phy_bit_cnt[0]),
	.b(i_tx_phy_bit_cnt[2]),
	.c(n450));
   oa12f01 U660 (.o(n453),
	.a(n451),
	.b(i_tx_phy_bit_cnt[0]),
	.c(n452));
   in01s01 U661 (.o(n459),
	.a(i_tx_phy_tx_ip_sync));
   ao12f01 U662 (.o(i_tx_phy_N87),
	.a(n459),
	.b(n454),
	.c(n453));
   in01s01 U663 (.o(n545),
	.a(i_rx_phy_bit_cnt[1]));
   na03s01 U664 (.o(n458),
	.a(n455),
	.b(i_rx_phy_bit_cnt[0]),
	.c(n545));
   in01s01 U665 (.o(n503),
	.a(i_rx_phy_shift_en));
   na02s01 U666 (.o(n89),
	.a(n458),
	.b(n457));
   no02f02 U667 (.o(n577),
	.a(n459),
	.b(n588));
   in01s01 U668 (.o(n460),
	.a(i_tx_phy_tx_ip));
   no02s01 U669 (.o(n461),
	.a(n460),
	.b(n590));
   no02s01 U670 (.o(n462),
	.a(n577),
	.b(n461));
   in01s01 U671 (.o(n134),
	.a(n462));
   in01s01 U672 (.o(n466),
	.a(i_rx_phy_one_cnt[1]));
   na02s01 U673 (.o(n464),
	.a(n466),
	.b(i_rx_phy_one_cnt[0]));
   no02s01 U674 (.o(n465),
	.a(n466),
	.b(i_rx_phy_one_cnt[2]));
   ao22s01 U675 (.o(n469),
	.a(n466),
	.b(i_rx_phy_one_cnt[2]),
	.c(n465),
	.d(i_rx_phy_one_cnt[0]));
   in01s01 U676 (.o(n468),
	.a(i_rx_phy_one_cnt[2]));
   in01s01 U677 (.o(n475),
	.a(n577));
   no02s01 U678 (.o(n473),
	.a(n576),
	.b(i_tx_phy_one_cnt[2]));
   ao22s01 U679 (.o(n474),
	.a(n576),
	.b(i_tx_phy_one_cnt[2]),
	.c(i_tx_phy_one_cnt[0]),
	.d(n473));
   oa22s01 U680 (.o(n116),
	.a(n476),
	.b(n475),
	.c(n581),
	.d(n474));
   ao12s01 U681 (.o(n478),
	.a(n550),
	.b(i_tx_phy_tx_ip),
	.c(n327));
   no02s01 U682 (.o(n135),
	.a(n583),
	.b(n478));
   no02s01 U683 (.o(n479),
	.a(n545),
	.b(i_rx_phy_bit_cnt[2]));
   ao22s01 U684 (.o(n482),
	.a(n545),
	.b(i_rx_phy_bit_cnt[2]),
	.c(i_rx_phy_bit_cnt[0]),
	.d(n479));
   oa12s01 U685 (.o(n88),
	.a(n481),
	.b(n483),
	.c(n482));
   na02s01 U686 (.o(n486),
	.a(n592),
	.b(i_rx_phy_rx_valid_r));
   ao22f01 U687 (.o(n487),
	.a(n486),
	.b(RxActive_o),
	.c(n500),
	.d(n489));
   no02f01 U688 (.o(n104),
	.a(n583),
	.b(n487));
   na03s01 U689 (.o(n490),
	.a(rst),
	.b(n492),
	.c(n498));
   oa22f01 U690 (.o(n105),
	.a(n496),
	.b(n490),
	.c(n498),
	.d(n493));
   in01s01 U691 (.o(n494),
	.a(i_rx_phy_fs_state[2]));
   oa22s01 U692 (.o(n491),
	.a(n498),
	.b(i_rx_phy_fs_state[2]),
	.c(i_rx_phy_fs_state[1]),
	.d(n494));
   na03f01 U693 (.o(n495),
	.a(rst),
	.b(n492),
	.c(n491));
   oa22f01 U694 (.o(n106),
	.a(n496),
	.b(n495),
	.c(n494),
	.d(n493));
   oa12s01 U695 (.o(n499),
	.a(n497),
	.b(n498),
	.c(i_rx_phy_rxdp_s));
   na02s01 U696 (.o(n504),
	.a(n327),
	.b(phy_tx_mode));
   oa22s01 U697 (.o(n506),
	.a(n504),
	.b(i_tx_phy_sd_nrzi_o),
	.c(n327),
	.d(phy_tx_mode));
   ao22s01 U698 (.o(n507),
	.a(n506),
	.b(n505),
	.c(txdn),
	.d(n585));
   in01s01 U699 (.o(n109),
	.a(n507));
   no02s01 U700 (.o(n511),
	.a(n510),
	.b(rst_cnt[1]));
   in01s01 U701 (.o(n140),
	.a(n512));
   na03s01 U702 (.o(n514),
	.a(i_tx_phy_bit_cnt[0]),
	.b(i_tx_phy_bit_cnt[1]),
	.c(n513));
   oa12s01 U703 (.o(n518),
	.a(n514),
	.b(n516),
	.c(n515));
   ao22f01 U704 (.o(n519),
	.a(n518),
	.b(n524),
	.c(i_tx_phy_bit_cnt[2]),
	.d(n523));
   in01s01 U705 (.o(n113),
	.a(n519));
   in01s01 U706 (.o(n525),
	.a(i_tx_phy_bit_cnt[0]));
   oa22s01 U707 (.o(n521),
	.a(n520),
	.b(i_tx_phy_bit_cnt[0]),
	.c(n525),
	.d(i_tx_phy_bit_cnt[1]));
   ao22f01 U708 (.o(n522),
	.a(n521),
	.b(n524),
	.c(i_tx_phy_bit_cnt[1]),
	.d(n523));
   in01s01 U709 (.o(n114),
	.a(n522));
   ao22f01 U710 (.o(n526),
	.a(n525),
	.b(n524),
	.c(i_tx_phy_bit_cnt[0]),
	.d(n523));
   in01s01 U711 (.o(n115),
	.a(n526));
   in01s01 U712 (.o(n566),
	.a(rst_cnt[2]));
   in01s01 U713 (.o(n528),
	.a(rst_cnt[1]));
   in01s01 U714 (.o(n530),
	.a(n529));
   in01s01 U715 (.o(n532),
	.a(n567));
   na02f01 U716 (.o(n534),
	.a(n577),
	.b(i_tx_phy_one_cnt[0]));
   in01s01 U717 (.o(n535),
	.a(n534));
   no02f01 U718 (.o(n536),
	.a(n578),
	.b(n535));
   in01s01 U719 (.o(n118),
	.a(n536));
   in01s01 U720 (.o(n546),
	.a(i_rx_phy_bit_cnt[2]));
   in01s01 U721 (.o(n544),
	.a(i_rx_phy_bit_cnt[0]));
   ao12f01 U722 (.o(n549),
	.a(n547),
	.b(i_rx_phy_rx_valid1),
	.c(n548));
   no02s01 U723 (.o(n87),
	.a(n583),
	.b(n549));
   no02f02 U724 (.o(n559),
	.a(n550),
	.b(i_tx_phy_ld_data));
   ao22s01 U725 (.o(n552),
	.a(n559),
	.b(i_tx_phy_hold_reg[4]),
	.c(n558),
	.d(DataOut_i[4]));
   in01s01 U726 (.o(n123),
	.a(n552));
   ao22s01 U727 (.o(n553),
	.a(n559),
	.b(i_tx_phy_hold_reg[6]),
	.c(n558),
	.d(DataOut_i[6]));
   in01s01 U728 (.o(n125),
	.a(n553));
   ao22s01 U729 (.o(n554),
	.a(n559),
	.b(i_tx_phy_hold_reg[0]),
	.c(n558),
	.d(DataOut_i[0]));
   in01s01 U730 (.o(n119),
	.a(n554));
   ao22s01 U731 (.o(n555),
	.a(n559),
	.b(i_tx_phy_hold_reg[1]),
	.c(n558),
	.d(DataOut_i[1]));
   in01s01 U732 (.o(n120),
	.a(n555));
   ao22s01 U733 (.o(n556),
	.a(n559),
	.b(i_tx_phy_hold_reg[2]),
	.c(n558),
	.d(DataOut_i[2]));
   in01s01 U734 (.o(n121),
	.a(n556));
   ao22s01 U735 (.o(n557),
	.a(n559),
	.b(i_tx_phy_hold_reg[3]),
	.c(n558),
	.d(DataOut_i[3]));
   in01s01 U736 (.o(n122),
	.a(n557));
   ao22s01 U737 (.o(n560),
	.a(n559),
	.b(i_tx_phy_hold_reg[5]),
	.c(n558),
	.d(DataOut_i[5]));
   in01s01 U738 (.o(n124),
	.a(n560));
   no02s01 U739 (.o(n568),
	.a(n566),
	.b(n565));
   in01s01 U740 (.o(n142),
	.a(n570));
   oa12s01 U741 (.o(n575),
	.a(n572),
	.b(n574),
	.c(n573));
   na02s01 U742 (.o(i_rx_phy_N31),
	.a(n575),
	.b(rst));
   na02s01 U743 (.o(n580),
	.a(n576),
	.b(i_tx_phy_one_cnt[0]));
   oa12f01 U744 (.o(n117),
	.a(n579),
	.b(n581),
	.c(n580));
   in01s01 U745 (.o(n582),
	.a(i_tx_phy_sd_bs_o));
   oa12s01 U746 (.o(n111),
	.a(n581),
	.b(n588),
	.c(n582));
   no02s01 U747 (.o(n584),
	.a(n583),
	.b(i_tx_phy_append_eop_sync4));
   no02s01 U748 (.o(n586),
	.a(n585),
	.b(n584));
   oa22s01 U749 (.o(n137),
	.a(n590),
	.b(n587),
	.c(n327),
	.d(n586));
   in01s01 U750 (.o(n589),
	.a(i_tx_phy_append_eop_sync4));
   oa22s01 U751 (.o(n136),
	.a(n590),
	.b(n327),
	.c(n589),
	.d(n588));
endmodule


/*
###############################################################
#  Design:            mpeg2_top
###############################################################
*/
module mpeg2_top (
	clk, 
	wbb_stb_i, 
	wbb_we_i, 
	wbb_adr_i, 
	wbb_dat_i, 
	wbb_dat_o, 
	wbb_ack_o, 
	v1_int18_n, 
	v1_int23_n, 
	v1_dmareq8_n, 
	mr_dmaack8_n, 
	sc_dmaack8_n, 
	y1_bs_wait_n, 
	v1_bs_req_n, 
	v1_sd_pichead_s, 
	y1_bs_data, 
	v1_dspfld_num1, 
	v1_dspfld_sc1, 
	v1_dspfld_num2, 
	v1_dspfld_sc2, 
	v1_dsp_ps, 
	vmem_wen, 
	vmem_we, 
	vmem_we_n, 
	vmem_ren, 
	vmem_add, 
	vmem_data_out, 
	vmem_data_in, 
	v_mode_mpeg1, 
	vmem_ch);
   input clk;
   input wbb_stb_i;
   input wbb_we_i;
   input [8:2] wbb_adr_i;
   input [31:0] wbb_dat_i;
   output [31:0] wbb_dat_o;
   output wbb_ack_o;
   output v1_int18_n;
   output v1_int23_n;
   output v1_dmareq8_n;
   input mr_dmaack8_n;
   input sc_dmaack8_n;
   input y1_bs_wait_n;
   output v1_bs_req_n;
   output v1_sd_pichead_s;
   input [31:0] y1_bs_data;
   output [3:0] v1_dspfld_num1;
   output v1_dspfld_sc1;
   output [3:0] v1_dspfld_num2;
   output v1_dspfld_sc2;
   output v1_dsp_ps;
   output vmem_wen;
   output [3:0] vmem_we;
   output [3:0] vmem_we_n;
   output vmem_ren;
   output [25:0] vmem_add;
   output [31:0] vmem_data_out;
   input [31:0] vmem_data_in;
   input v_mode_mpeg1;
   input vmem_ch;

   // Internal wires
   wire FE_OCPN583_n247126;
   wire FE_OCPN582_n247126;
   wire FE_OFN581_n248442;
   wire FE_OFN580_n248442;
   wire FE_OFN579_n248820;
   wire FE_OFN578_n248820;
   wire FE_OFN577_n247126;
   wire FE_OFN576_n247126;
   wire FE_OFN575_n245444;
   wire FE_OFN574_n245444;
   wire FE_OFN573_n249242;
   wire FE_OFN572_n249242;
   wire FE_OFN571_n248074;
   wire FE_OFN570_n248074;
   wire FE_OFN569_n247780;
   wire FE_OFN568_n247780;
   wire FE_OFN567_n247541;
   wire FE_OFN566_n247541;
   wire FE_OFN565_n247738;
   wire FE_OFN564_n247738;
   wire FE_OFN563_n250717;
   wire FE_OFN562_n250717;
   wire FE_OFN561_n251852;
   wire FE_OFN560_n251852;
   wire FE_OFN559_n251852;
   wire FE_OFN558_n252630;
   wire FE_OFN557_n252630;
   wire FE_OFN556_n250770;
   wire FE_OFN555_n250770;
   wire FE_OFN554_n247778;
   wire FE_OFN553_n247778;
   wire FE_RN_9_0;
   wire FE_RN_8_0;
   wire FE_RN_7_0;
   wire FE_RN_6_0;
   wire FE_RN_5_0;
   wire FE_RN_4_0;
   wire FE_RN_3_0;
   wire FE_RN_2_0;
   wire FE_RN_1_0;
   wire FE_RN_0_0;
   wire FE_OFN552_n245462;
   wire FE_OFN551_n249140;
   wire FE_OFN550_n249113;
   wire FE_OFN549_regtop_g_a_r_2_;
   wire FE_OFN548_regtop_g_a_r_2_;
   wire FE_OFN547_n245460;
   wire FE_OFN546_n245460;
   wire FE_OFN545_n245460;
   wire FE_OFN544_n252912;
   wire FE_OFN543_vldtop_vld_syndec_vld_vlfeed_lower_26_;
   wire FE_OFN542_n248424;
   wire FE_OFN541_n248424;
   wire FE_OFN540_vldtop_vld_syndec_vld_vlfeed_lower_12_;
   wire FE_OFN537_vldtop_vld_syndec_vld_vlfeed_lower_18_;
   wire FE_OFN534_regtop_g_a_r_5_;
   wire FE_OFN532_regtop_g_a_r_5_;
   wire FE_OFN530_vldtop_vld_syndec_vld_vlfeed_lower_14_;
   wire FE_OFN527_n249828;
   wire FE_OFN526_n249548;
   wire FE_OFN525_vldtop_vld_syndec_vld_vlfeed_lower_16_;
   wire FE_OFN524_n247696;
   wire FE_OFN523_n247696;
   wire FE_OFN522_n248508;
   wire FE_OFN521_n248508;
   wire FE_OFN520_regtop_g_a_r_6_;
   wire FE_OFN519_regtop_g_a_r_6_;
   wire FE_OFN517_regtop_g_a_r_6_;
   wire FE_OFN516_regtop_v1_hdi00_a_0_;
   wire FE_OFN514_n247538;
   wire FE_OFN513_n247538;
   wire FE_OFN512_n248634;
   wire FE_OFN511_n248634;
   wire FE_OFN510_regtop_g_a_r_7_;
   wire FE_OFN509_regtop_g_a_r_7_;
   wire FE_OFN508_n252540;
   wire FE_OFN507_regtop_g_a_r_4_;
   wire FE_OFN506_regtop_g_a_r_4_;
   wire FE_OFN505_regtop_g_a_r_4_;
   wire FE_OFN504_regtop_g_a_r_4_;
   wire FE_OFN503_n246205;
   wire FE_OFN502_n246205;
   wire FE_OFN501_n246205;
   wire FE_OFN500_n246205;
   wire FE_OFN499_n253015;
   wire FE_OFN498_n253015;
   wire FE_OFN497_n249947;
   wire FE_OFN496_n249242;
   wire FE_OFN494_n252377;
   wire FE_OFN493_n252377;
   wire FE_OFN492_n252377;
   wire FE_OFN491_regtop_g_a_r_3_;
   wire FE_OFN490_regtop_g_a_r_3_;
   wire FE_OFN489_n249763;
   wire FE_OFN488_n245940;
   wire FE_OFN486_n245940;
   wire FE_OFN485_n245940;
   wire FE_OFN484_n245940;
   wire FE_OFN483_n249211;
   wire FE_OFN478_n249800;
   wire FE_OFN477_n249800;
   wire FE_OFN472_n244982;
   wire FE_OFN471_n244982;
   wire FE_OFN470_n244978;
   wire FE_OFN469_n244978;
   wire FE_OFN468_n244218;
   wire FE_OFN467_n244218;
   wire FE_OFN466_n249845;
   wire FE_OFN465_n249845;
   wire FE_OFN464_n249821;
   wire FE_OFN463_n249821;
   wire FE_OFN462_n249378;
   wire FE_OFN461_n249378;
   wire FE_OFN458_n252996;
   wire FE_OFN457_n252996;
   wire FE_OFN456_n252942;
   wire FE_OFN455_n252942;
   wire FE_OFN454_n252863;
   wire FE_OFN453_n252863;
   wire FE_OFN449_n249831;
   wire FE_OFN448_n249831;
   wire FE_OFN445_n249391;
   wire FE_OFN444_n249391;
   wire FE_OFN441_n252905;
   wire FE_OFN440_n252905;
   wire FE_OFN439_n252264;
   wire FE_OFN437_n252069;
   wire FE_OFN436_n252069;
   wire FE_OFN435_n252069;
   wire FE_OFN434_n251996;
   wire FE_OFN433_n251996;
   wire FE_OFN432_n251781;
   wire FE_OFN431_n251781;
   wire FE_OFN430_n251710;
   wire FE_OFN429_n251710;
   wire FE_OFN428_n251494;
   wire FE_OFN427_n251494;
   wire FE_OFN426_n251424;
   wire FE_OFN425_n251424;
   wire FE_OFN424_n251300;
   wire FE_OFN423_n251300;
   wire FE_OFN422_n251211;
   wire FE_OFN421_n251211;
   wire FE_OFN420_n251140;
   wire FE_OFN419_n251140;
   wire FE_OFN418_n250930;
   wire FE_OFN417_n250930;
   wire FE_OFN416_n250859;
   wire FE_OFN415_n250859;
   wire FE_OFN414_n250646;
   wire FE_OFN413_n250646;
   wire FE_OFN412_n250576;
   wire FE_OFN411_n250576;
   wire FE_OFN410_n250360;
   wire FE_OFN409_n250360;
   wire FE_OFN408_n250289;
   wire FE_OFN407_n250289;
   wire FE_OFN406_n250162;
   wire FE_OFN405_n250162;
   wire FE_OFN404_n250071;
   wire FE_OFN403_n250071;
   wire FE_OFN402_n249999;
   wire FE_OFN401_n249999;
   wire FE_OFN400_n249836;
   wire FE_OFN399_n249836;
   wire FE_OFN398_n249646;
   wire FE_OFN397_n249646;
   wire FE_OFN396_n249640;
   wire FE_OFN395_n249640;
   wire FE_OFN392_n249635;
   wire FE_OFN391_n249635;
   wire FE_OFN390_n249480;
   wire FE_OFN389_n249480;
   wire FE_OFN388_n249468;
   wire FE_OFN387_n249468;
   wire FE_OFN386_n248760;
   wire FE_OFN385_n248760;
   wire FE_OFN384_n248677;
   wire FE_OFN383_n248677;
   wire FE_OFN382_n248549;
   wire FE_OFN381_n248549;
   wire FE_OFN376_n248352;
   wire FE_OFN375_n248352;
   wire FE_OFN374_n248311;
   wire FE_OFN373_n248311;
   wire FE_OFN372_n247737;
   wire FE_OFN371_n247737;
   wire FE_OFN368_n247123;
   wire FE_OFN367_n247123;
   wire FE_OFN366_n246266;
   wire FE_OFN365_n246266;
   wire FE_OFN362_n252748;
   wire FE_OFN361_n252748;
   wire FE_OFN360_n252728;
   wire FE_OFN359_n252728;
   wire FE_OFN356_n252508;
   wire FE_OFN355_n252508;
   wire FE_OFN354_n252338;
   wire FE_OFN353_n252338;
   wire FE_OFN352_n252242;
   wire FE_OFN351_n252242;
   wire FE_OFN350_n252215;
   wire FE_OFN349_n252215;
   wire FE_OFN348_n252178;
   wire FE_OFN347_n252178;
   wire FE_OFN346_n252141;
   wire FE_OFN345_n252141;
   wire FE_OFN344_n252141;
   wire FE_OFN343_n252032;
   wire FE_OFN342_n252032;
   wire FE_OFN341_n251960;
   wire FE_OFN340_n251960;
   wire FE_OFN339_n251923;
   wire FE_OFN338_n251923;
   wire FE_OFN337_n251887;
   wire FE_OFN336_n251887;
   wire FE_OFN335_n251852;
   wire FE_OFN334_n251852;
   wire FE_OFN333_n251746;
   wire FE_OFN332_n251746;
   wire FE_OFN331_n251675;
   wire FE_OFN330_n251675;
   wire FE_OFN329_n251637;
   wire FE_OFN328_n251637;
   wire FE_OFN327_n251600;
   wire FE_OFN326_n251600;
   wire FE_OFN325_n251565;
   wire FE_OFN324_n251565;
   wire FE_OFN323_n251565;
   wire FE_OFN322_n251459;
   wire FE_OFN321_n251459;
   wire FE_OFN320_n251388;
   wire FE_OFN319_n251388;
   wire FE_OFN318_n251353;
   wire FE_OFN317_n251353;
   wire FE_OFN316_n251317;
   wire FE_OFN315_n251317;
   wire FE_OFN314_n251281;
   wire FE_OFN313_n251281;
   wire FE_OFN312_n251281;
   wire FE_OFN311_n251175;
   wire FE_OFN310_n251175;
   wire FE_OFN309_n251105;
   wire FE_OFN308_n251105;
   wire FE_OFN307_n251072;
   wire FE_OFN306_n251072;
   wire FE_OFN305_n251072;
   wire FE_OFN304_n251036;
   wire FE_OFN303_n251036;
   wire FE_OFN302_n251001;
   wire FE_OFN301_n251001;
   wire FE_OFN300_n250895;
   wire FE_OFN299_n250895;
   wire FE_OFN298_n250824;
   wire FE_OFN297_n250824;
   wire FE_OFN296_n250789;
   wire FE_OFN295_n250789;
   wire FE_OFN294_n250752;
   wire FE_OFN293_n250752;
   wire FE_OFN292_n250717;
   wire FE_OFN291_n250717;
   wire FE_OFN290_n250611;
   wire FE_OFN289_n250611;
   wire FE_OFN288_n250540;
   wire FE_OFN287_n250540;
   wire FE_OFN286_n250502;
   wire FE_OFN285_n250502;
   wire FE_OFN284_n250466;
   wire FE_OFN283_n250466;
   wire FE_OFN282_n250430;
   wire FE_OFN281_n250430;
   wire FE_OFN280_n250324;
   wire FE_OFN279_n250324;
   wire FE_OFN278_n250254;
   wire FE_OFN277_n250254;
   wire FE_OFN276_n250218;
   wire FE_OFN275_n250218;
   wire FE_OFN274_n250180;
   wire FE_OFN273_n250180;
   wire FE_OFN272_n250144;
   wire FE_OFN271_n250144;
   wire FE_OFN270_n250035;
   wire FE_OFN269_n250035;
   wire FE_OFN268_n249964;
   wire FE_OFN267_n249964;
   wire FE_OFN266_n249787;
   wire FE_OFN265_n249787;
   wire FE_OFN264_n249636;
   wire FE_OFN263_n249636;
   wire FE_OFN256_n248843;
   wire FE_OFN255_n248843;
   wire FE_OFN252_n248799;
   wire FE_OFN251_n248799;
   wire FE_OFN248_n248527;
   wire FE_OFN247_n248527;
   wire FE_OFN246_n248465;
   wire FE_OFN245_n248465;
   wire FE_OFN244_n248463;
   wire FE_OFN243_n248463;
   wire FE_OFN240_n248389;
   wire FE_OFN239_n248389;
   wire FE_OFN236_n248245;
   wire FE_OFN235_n248245;
   wire FE_OFN234_n248115;
   wire FE_OFN233_n248115;
   wire FE_OFN230_n247987;
   wire FE_OFN229_n247987;
   wire FE_OFN228_n247903;
   wire FE_OFN227_n247903;
   wire FE_OFN220_n246261;
   wire FE_OFN219_n246261;
   wire FE_OFN218_n246238;
   wire FE_OFN217_n246238;
   wire FE_OFN214_n252483;
   wire FE_OFN213_n252483;
   wire FE_OFN212_n252422;
   wire FE_OFN211_n252422;
   wire FE_OFN210_n252159;
   wire FE_OFN209_n252159;
   wire FE_OFN208_n252105;
   wire FE_OFN207_n252105;
   wire FE_OFN206_n251816;
   wire FE_OFN205_n251816;
   wire FE_OFN204_n251530;
   wire FE_OFN203_n251530;
   wire FE_OFN202_n251246;
   wire FE_OFN201_n251246;
   wire FE_OFN200_n250965;
   wire FE_OFN199_n250965;
   wire FE_OFN198_n250682;
   wire FE_OFN197_n250682;
   wire FE_OFN196_n250682;
   wire FE_OFN195_n250395;
   wire FE_OFN194_n250395;
   wire FE_OFN193_n250107;
   wire FE_OFN192_n250107;
   wire FE_OFN191_n250107;
   wire FE_OFN185_n248415;
   wire FE_OFN184_n248415;
   wire FE_OFN183_n248414;
   wire FE_OFN182_n248414;
   wire FE_OFN181_n248413;
   wire FE_OFN180_n248413;
   wire FE_OFN179_n248408;
   wire FE_OFN178_n248408;
   wire FE_OFN177_n248407;
   wire FE_OFN176_n248407;
   wire FE_OFN175_n248406;
   wire FE_OFN174_n248406;
   wire FE_OFN173_n248405;
   wire FE_OFN172_n248405;
   wire FE_OFN171_n248404;
   wire FE_OFN170_n248404;
   wire FE_OFN169_n248399;
   wire FE_OFN168_n248399;
   wire FE_OFN167_n248398;
   wire FE_OFN166_n248398;
   wire FE_OFN165_n248393;
   wire FE_OFN164_n248393;
   wire FE_OFN163_n248392;
   wire FE_OFN162_n248392;
   wire FE_OFN161_n248391;
   wire FE_OFN160_n248391;
   wire FE_OFN159_n248382;
   wire FE_OFN158_n248382;
   wire FE_OFN157_n248381;
   wire FE_OFN156_n248381;
   wire FE_OFN155_n248380;
   wire FE_OFN154_n248380;
   wire FE_OFN153_n248375;
   wire FE_OFN152_n248375;
   wire FE_OFN151_n248374;
   wire FE_OFN150_n248374;
   wire FE_OFN149_n248373;
   wire FE_OFN148_n248373;
   wire FE_OFN147_n248372;
   wire FE_OFN146_n248372;
   wire FE_OFN145_n248372;
   wire FE_OFN144_n248371;
   wire FE_OFN143_n248371;
   wire FE_OFN142_n248370;
   wire FE_OFN141_n248370;
   wire FE_OFN140_n248369;
   wire FE_OFN139_n248369;
   wire FE_OFN138_n248364;
   wire FE_OFN137_n248364;
   wire FE_OFN136_n248363;
   wire FE_OFN135_n248363;
   wire FE_OFN134_n248362;
   wire FE_OFN133_n248362;
   wire FE_OFN132_n248357;
   wire FE_OFN131_n248357;
   wire FE_OFN130_n248356;
   wire FE_OFN129_n248356;
   wire FE_OFN128_n248355;
   wire FE_OFN127_n248355;
   wire FE_OFN126_n248176;
   wire FE_OFN125_n248176;
   wire FE_OFN124_n248175;
   wire FE_OFN123_n248175;
   wire FE_OFN122_n248174;
   wire FE_OFN121_n248174;
   wire FE_OFN120_n248173;
   wire FE_OFN119_n248173;
   wire FE_OFN116_n248167;
   wire FE_OFN115_n248167;
   wire FE_OFN114_n248162;
   wire FE_OFN113_n248162;
   wire FE_OFN112_n248162;
   wire FE_OFN109_n248160;
   wire FE_OFN108_n248160;
   wire FE_OFN107_n248160;
   wire FE_OFN106_n248159;
   wire FE_OFN105_n248159;
   wire FE_OFN104_n248158;
   wire FE_OFN103_n248158;
   wire FE_OFN102_n248153;
   wire FE_OFN101_n248153;
   wire FE_OFN100_n248152;
   wire FE_OFN99_n248152;
   wire FE_OFN98_n248151;
   wire FE_OFN97_n248151;
   wire FE_OFN96_n248150;
   wire FE_OFN95_n248150;
   wire FE_OFN94_n248141;
   wire FE_OFN93_n248141;
   wire FE_OFN90_n248139;
   wire FE_OFN89_n248139;
   wire FE_OFN88_n248138;
   wire FE_OFN87_n248138;
   wire FE_OFN86_n248129;
   wire FE_OFN85_n248129;
   wire FE_OFN84_n248128;
   wire FE_OFN83_n248128;
   wire FE_OFN82_n248127;
   wire FE_OFN81_n248127;
   wire FE_OFN80_n248127;
   wire FE_OFN79_n248126;
   wire FE_OFN78_n248126;
   wire FE_OFN77_n248121;
   wire FE_OFN76_n248121;
   wire FE_OFN75_n248120;
   wire FE_OFN74_n248120;
   wire FE_OFN73_n248119;
   wire FE_OFN72_n248119;
   wire FE_OFN71_n248119;
   wire FE_OFN70_n248118;
   wire FE_OFN69_n248118;
   wire FE_OFN68_n247591;
   wire FE_OFN67_n247591;
   wire FE_OFN66_n247531;
   wire FE_OFN65_n247531;
   wire FE_OFN64_n247509;
   wire FE_OFN63_n247509;
   wire FE_OFN62_n247107;
   wire FE_OFN61_n247107;
   wire FE_OFN60_n247099;
   wire FE_OFN59_n247099;
   wire FE_OFN58_n247092;
   wire FE_OFN57_n247092;
   wire FE_OFN56_n247074;
   wire FE_OFN55_n247074;
   wire FE_OFN54_n247067;
   wire FE_OFN53_n247067;
   wire FE_OFN52_n247067;
   wire FE_OFN51_n247057;
   wire FE_OFN50_n247057;
   wire FE_OFN45_n252700;
   wire FE_OFN44_n252700;
   wire FE_OFN43_n252668;
   wire FE_OFN42_n252668;
   wire FE_OFN41_n252640;
   wire FE_OFN40_n252640;
   wire FE_OFN39_n252462;
   wire FE_OFN38_n252462;
   wire FE_OFN37_n252446;
   wire FE_OFN36_n252446;
   wire FE_OFN33_n251904;
   wire FE_OFN32_n251904;
   wire FE_OFN31_n251904;
   wire FE_OFN28_n251337;
   wire FE_OFN27_n251337;
   wire FE_OFN24_n250486;
   wire FE_OFN23_n250486;
   wire FE_OFN22_n250202;
   wire FE_OFN21_n250202;
   wire FE_OFN20_n249394;
   wire FE_OFN19_n249394;
   wire FE_OFN18_n247494;
   wire FE_OFN17_n247494;
   wire FE_OFN16_n247350;
   wire FE_OFN15_n247350;
   wire FE_OFN14_n247150;
   wire FE_OFN13_n247150;
   wire FE_OFN8_n247076;
   wire FE_OFN7_n247076;
   wire FE_OFN6_n246618;
   wire FE_OFN5_n246618;
   wire FE_OFN4_n245443;
   wire FE_OFN3_n245443;
   wire FE_OFN2_g_swrst_r_n;
   wire FE_OFN1_g_swrst_r_n;
   wire g_mbc_en_r;
   wire g_pmod_r;
   wire g_swrst_r_n;
   wire g_vden_r;
   wire g_fcyc_en_r;
   wire v_ferror_r;
   wire v_seqstrt_r;
   wire c_tmg_ferr_hit_r;
   wire v_nferror_r;
   wire g_init_vld_r_s;
   wire g_line_offset_r;
   wire g_bmod_r;
   wire cntrltop_ctmg_ctpedet_N22;
   wire cntrltop_ctmg_ctpedet_c_tmg_ferr_pre_d1_r;
   wire cntrltop_ctmg_ctpedet_c_tmg_ferr_pre;
   wire cntrltop_ctmg_ctpedet_c_bigpictdet_r;
   wire vldtop_vld_syndec_vld_seqhed_state_0_;
   wire vldtop_vld_syndec_vld_outbuf_N487;
   wire vldtop_vld_syndec_vld_outbuf_N486;
   wire vldtop_vld_syndec_vld_outbuf_N485;
   wire vldtop_vld_syndec_vld_outbuf_N484;
   wire vldtop_vld_syndec_vld_outbuf_N483;
   wire vldtop_vld_syndec_vld_outbuf_N482;
   wire vldtop_vld_syndec_vld_outbuf_N481;
   wire vldtop_vld_syndec_vld_outbuf_N480;
   wire vldtop_vld_syndec_vld_outbuf_N479;
   wire vldtop_vld_syndec_vld_outbuf_N478;
   wire vldtop_vld_syndec_vld_outbuf_N477;
   wire vldtop_vld_syndec_vld_outbuf_N476;
   wire vldtop_vld_syndec_vld_outbuf_N475;
   wire vldtop_vld_syndec_vld_outbuf_N474;
   wire vldtop_vld_syndec_vld_outbuf_N473;
   wire vldtop_vld_syndec_vld_outbuf_N472;
   wire vldtop_vld_syndec_vld_outbuf_N471;
   wire vldtop_vld_syndec_vld_outbuf_N470;
   wire vldtop_vld_syndec_vld_outbuf_N469;
   wire vldtop_vld_syndec_vld_outbuf_N468;
   wire vldtop_vld_syndec_vld_outbuf_N467;
   wire vldtop_vld_syndec_vld_outbuf_N466;
   wire vldtop_vld_syndec_vld_outbuf_N465;
   wire vldtop_vld_syndec_vld_outbuf_N464;
   wire vldtop_vld_syndec_vld_outbuf_N463;
   wire vldtop_vld_syndec_vld_outbuf_N52;
   wire vldtop_vld_syndec_vld_outbuf_N46;
   wire vldtop_vld_syndec_vld_outbuf_N44;
   wire vldtop_vld_syndec_vld_vscdet_v_search_1st_r;
   wire vldtop_vld_syndec_vld_vscdet_v_seqerr_r;
   wire vldtop_vld_syndec_vld_vlfeed_dselect_r;
   wire vldtop_vld_syndec_vld_vlfeed_feed_on;
   wire busrtop_b_rreq_N431;
   wire busrtop_b_rreq_N430;
   wire busrtop_b_rreq_N429;
   wire busrtop_b_rreq_N428;
   wire busrtop_b_rreq_N427;
   wire busrtop_b_rreq_N426;
   wire busrtop_b_rreq_N425;
   wire busrtop_b_rreq_N424;
   wire busrtop_b_rreq_N423;
   wire busrtop_b_rreq_N296;
   wire busrtop_b_rreq_N295;
   wire busrtop_b_rreq_N229;
   wire busrtop_b_rreq_N106;
   wire busrtop_b_rreq_N105;
   wire busrtop_b_rreq_N104;
   wire busrtop_b_rreq_N103;
   wire busrtop_b_rreq_N102;
   wire busrtop_b_rreq_N101;
   wire busrtop_b_rreq_N100;
   wire busrtop_b_rreq_N99;
   wire busrtop_b_rreq_N98;
   wire busrtop_b_rreq_N97;
   wire busrtop_b_rreq_N96;
   wire busrtop_b_rreq_N95;
   wire busrtop_b_rreq_N94;
   wire busrtop_b_rreq_N93;
   wire busrtop_b_rreq_N92;
   wire busrtop_b_rreq_N91;
   wire busrtop_b_rreq_N90;
   wire busrtop_b_rreq_N89;
   wire busrtop_b_rreq_N88;
   wire busrtop_b_rreq_N87;
   wire busrtop_b_rreq_N86;
   wire busrtop_b_rreq_N85;
   wire regtop_N2024;
   wire regtop_N2023;
   wire regtop_N2022;
   wire regtop_N2021;
   wire regtop_N2020;
   wire regtop_N2019;
   wire regtop_N2018;
   wire regtop_N2017;
   wire regtop_N2016;
   wire regtop_N2015;
   wire regtop_N2014;
   wire regtop_N2013;
   wire regtop_N2012;
   wire regtop_N2011;
   wire regtop_N2010;
   wire regtop_N2009;
   wire regtop_N2008;
   wire regtop_N2007;
   wire regtop_N2006;
   wire regtop_N2005;
   wire regtop_N2004;
   wire regtop_N2003;
   wire regtop_N2002;
   wire regtop_N2001;
   wire regtop_N2000;
   wire regtop_N1999;
   wire regtop_N1998;
   wire regtop_N1997;
   wire regtop_N1996;
   wire regtop_N1995;
   wire regtop_N1994;
   wire regtop_N1993;
   wire regtop_g_rd_en_r;
   wire regtop_g_rd_en2_r;
   wire regtop_N1991;
   wire regtop_N1990;
   wire regtop_v1_hdi00_we;
   wire regtop_v1_hdi00_bs;
   wire regtop_g_sc_r;
   wire regtop_g_va_r;
   wire regtop_g_cdf_r;
   wire regtop_g_pf_r;
   wire regtop_g_rff_r;
   wire regtop_g_tff_r;
   wire regtop_g_bl_r;
   wire regtop_g_cg_r;
   wire regtop_g_cd_r;
   wire regtop_g_ld_r;
   wire regtop_g_ps_r;
   wire regtop_g_cpf_r;
   wire regtop_g_hclr_r_s;
   wire regtop_g_dcnt_r;
   wire regtop_N1279;
   wire regtop_g_prev_enfst_r;
   wire regtop_N1267;
   wire regtop_g_prev_efbst_r;
   wire regtop_g_issh_r;
   wire regtop_g_ispi_r;
   wire regtop_g_issr_r;
   wire regtop_g_issw_r;
   wire regtop_g_isuc_r;
   wire regtop_g_isdc_r;
   wire regtop_g_isnf_r;
   wire regtop_g_isfb_r;
   wire regtop_g_dsts_r;
   wire regtop_g_isph_r;
   wire regtop_g_isfp_r;
   wire regtop_g_icsh_r;
   wire regtop_g_icph_r;
   wire regtop_g_icpi_r;
   wire regtop_g_icnf_r;
   wire regtop_g_icfb_r;
   wire regtop_g_icfp_r;
   wire regtop_g_icsr_r;
   wire regtop_g_icsw_r;
   wire regtop_g_icuc_r;
   wire regtop_g_icdc_r;
   wire regtop_g_mpeg_r;
   wire regtop_g_imod_r;
   wire regtop_g_dmod_r;
   wire regtop_g_memr_ok_r;
   wire regtop_g_tmg_ferr_hit_r;
   wire regtop_g_nferror_r;
   wire regtop_g_ferror_r;
   wire regtop_g_seqstrt_r;
   wire regtop_g_dacksh_r_n;
   wire regtop_g_dack32_r_n;
   wire regtop_g_write_r_n;
   wire regtop_g_read_r_n;
   wire regtop_g_ms_r_n;
   wire busiftop_status_b_current_0_;
   wire busiftop_N61;
   wire busiftop_N60;
   wire busiftop_N59;
   wire busiftop_N58;
   wire busiftop_N57;
   wire busiftop_N56;
   wire busiftop_N55;
   wire busiftop_N54;
   wire busiftop_N53;
   wire busiftop_N52;
   wire busiftop_N51;
   wire busiftop_N50;
   wire busiftop_N49;
   wire busiftop_N48;
   wire busiftop_N47;
   wire busiftop_N46;
   wire busiftop_N45;
   wire busiftop_N44;
   wire busiftop_N43;
   wire busiftop_N42;
   wire busiftop_N41;
   wire busiftop_N40;
   wire busiftop_N39;
   wire busiftop_N38;
   wire busiftop_N37;
   wire busiftop_N36;
   wire busiftop_N35;
   wire busiftop_vmem_ren_g;
   wire busiftop_vmem_ch_r;
   wire busiftop_N32;
   wire busiftop_N28;
   wire n157815;
   wire n157831;
   wire n157832;
   wire n157833;
   wire n157834;
   wire n157835;
   wire n157836;
   wire n157837;
   wire n157838;
   wire n157839;
   wire n157840;
   wire n162088;
   wire n170932;
   wire n170937;
   wire n170938;
   wire n170939;
   wire n170951;
   wire n170952;
   wire n170953;
   wire n170954;
   wire n170955;
   wire n170956;
   wire n170957;
   wire n170958;
   wire n170959;
   wire n170960;
   wire n170961;
   wire n170962;
   wire n170963;
   wire n170964;
   wire n170965;
   wire n184629;
   wire n184630;
   wire n184631;
   wire n184632;
   wire n184633;
   wire n184634;
   wire n184635;
   wire n184636;
   wire n184637;
   wire n184638;
   wire n184639;
   wire n184640;
   wire n184641;
   wire n184642;
   wire n184643;
   wire n184644;
   wire n184645;
   wire n184646;
   wire n184647;
   wire n184648;
   wire n184649;
   wire n184650;
   wire n184651;
   wire n184652;
   wire n184653;
   wire n184654;
   wire n184655;
   wire n184656;
   wire n184657;
   wire n184658;
   wire n184659;
   wire n184660;
   wire n184661;
   wire n184662;
   wire n184663;
   wire n184664;
   wire n184665;
   wire n184666;
   wire n184667;
   wire n184668;
   wire n184669;
   wire n184670;
   wire n184671;
   wire n184672;
   wire n184673;
   wire n184674;
   wire n184675;
   wire n184676;
   wire n184677;
   wire n184678;
   wire n184679;
   wire n184680;
   wire n184681;
   wire n184682;
   wire n184683;
   wire n184684;
   wire n184685;
   wire n184686;
   wire n184687;
   wire n184688;
   wire n184689;
   wire n184690;
   wire n184691;
   wire n184692;
   wire n184693;
   wire n184694;
   wire n184695;
   wire n184696;
   wire n184697;
   wire n184698;
   wire n184699;
   wire n184700;
   wire n184701;
   wire n184702;
   wire n184703;
   wire n184704;
   wire n184705;
   wire n184706;
   wire n184707;
   wire n184708;
   wire n184709;
   wire n184710;
   wire n184711;
   wire n184712;
   wire n184713;
   wire n184714;
   wire n184715;
   wire n184716;
   wire n184717;
   wire n184718;
   wire n184719;
   wire n184720;
   wire n184721;
   wire n184722;
   wire n184723;
   wire n184724;
   wire n184725;
   wire n184726;
   wire n184727;
   wire n184728;
   wire n184729;
   wire n184730;
   wire n184731;
   wire n184732;
   wire n184733;
   wire n184734;
   wire n184735;
   wire n184736;
   wire n184737;
   wire n184738;
   wire n184739;
   wire n184740;
   wire n184741;
   wire n184742;
   wire n184743;
   wire n184744;
   wire n184745;
   wire n184746;
   wire n184747;
   wire n184748;
   wire n184749;
   wire n184750;
   wire n184751;
   wire n184752;
   wire n184753;
   wire n184754;
   wire n184755;
   wire n184756;
   wire n184757;
   wire n184758;
   wire n184759;
   wire n184760;
   wire n184761;
   wire n184762;
   wire n184763;
   wire n184764;
   wire n184765;
   wire n184766;
   wire n184767;
   wire n184768;
   wire n184769;
   wire n184770;
   wire n184771;
   wire n184772;
   wire n184773;
   wire n184774;
   wire n184775;
   wire n184776;
   wire n184777;
   wire n184778;
   wire n184779;
   wire n184780;
   wire n184781;
   wire n184782;
   wire n184783;
   wire n184784;
   wire n184785;
   wire n184786;
   wire n184787;
   wire n184788;
   wire n184789;
   wire n184790;
   wire n184791;
   wire n184792;
   wire n184793;
   wire n184794;
   wire n184795;
   wire n184796;
   wire n184797;
   wire n184798;
   wire n184799;
   wire n184800;
   wire n184801;
   wire n184802;
   wire n184803;
   wire n184804;
   wire n184805;
   wire n184806;
   wire n184807;
   wire n184808;
   wire n184809;
   wire n184810;
   wire n184811;
   wire n184812;
   wire n184813;
   wire n184814;
   wire n184815;
   wire n184816;
   wire n184817;
   wire n184818;
   wire n184819;
   wire n184820;
   wire n184821;
   wire n184822;
   wire n184823;
   wire n184824;
   wire n184825;
   wire n184826;
   wire n184827;
   wire n184828;
   wire n184829;
   wire n184830;
   wire n184831;
   wire n184832;
   wire n184833;
   wire n184834;
   wire n184835;
   wire n184836;
   wire n184837;
   wire n184838;
   wire n184839;
   wire n184840;
   wire n184841;
   wire n184842;
   wire n184843;
   wire n184844;
   wire n184845;
   wire n184846;
   wire n184847;
   wire n184848;
   wire n184849;
   wire n184850;
   wire n184851;
   wire n184852;
   wire n184853;
   wire n184854;
   wire n184855;
   wire n184856;
   wire n184857;
   wire n184858;
   wire n184859;
   wire n184860;
   wire n184861;
   wire n184862;
   wire n184863;
   wire n184864;
   wire n184865;
   wire n184866;
   wire n184867;
   wire n184868;
   wire n184869;
   wire n184870;
   wire n184871;
   wire n184872;
   wire n184873;
   wire n184874;
   wire n184875;
   wire n184876;
   wire n184877;
   wire n184878;
   wire n184879;
   wire n184880;
   wire n184881;
   wire n184882;
   wire n184883;
   wire n184884;
   wire n184885;
   wire n184886;
   wire n184887;
   wire n184888;
   wire n184889;
   wire n184890;
   wire n184891;
   wire n184892;
   wire n184893;
   wire n184894;
   wire n184895;
   wire n184896;
   wire n184897;
   wire n184898;
   wire n184899;
   wire n184900;
   wire n184901;
   wire n184902;
   wire n184903;
   wire n184904;
   wire n184905;
   wire n184906;
   wire n184907;
   wire n184908;
   wire n184909;
   wire n184910;
   wire n184911;
   wire n184912;
   wire n184913;
   wire n184914;
   wire n184915;
   wire n184916;
   wire n184917;
   wire n184918;
   wire n184919;
   wire n184920;
   wire n184921;
   wire n184922;
   wire n184923;
   wire n184924;
   wire n184925;
   wire n184926;
   wire n184927;
   wire n184928;
   wire n184929;
   wire n184930;
   wire n184931;
   wire n184932;
   wire n184933;
   wire n184934;
   wire n184935;
   wire n184936;
   wire n184937;
   wire n184938;
   wire n184939;
   wire n184940;
   wire n184941;
   wire n184942;
   wire n184943;
   wire n184944;
   wire n184945;
   wire n184946;
   wire n184947;
   wire n184948;
   wire n184949;
   wire n184950;
   wire n184951;
   wire n184952;
   wire n184953;
   wire n184954;
   wire n184955;
   wire n184956;
   wire n184957;
   wire n184958;
   wire n184959;
   wire n184960;
   wire n184961;
   wire n184962;
   wire n184963;
   wire n184964;
   wire n184965;
   wire n184966;
   wire n184967;
   wire n184968;
   wire n184969;
   wire n184970;
   wire n184971;
   wire n184972;
   wire n184973;
   wire n184974;
   wire n184975;
   wire n184976;
   wire n184977;
   wire n184978;
   wire n184979;
   wire n184980;
   wire n184981;
   wire n184982;
   wire n184983;
   wire n184984;
   wire n184985;
   wire n184986;
   wire n184987;
   wire n184988;
   wire n184989;
   wire n184990;
   wire n184991;
   wire n184992;
   wire n184993;
   wire n184994;
   wire n184995;
   wire n184996;
   wire n184997;
   wire n184998;
   wire n184999;
   wire n185000;
   wire n185001;
   wire n185002;
   wire n185003;
   wire n185004;
   wire n185005;
   wire n185006;
   wire n185007;
   wire n185008;
   wire n185009;
   wire n185010;
   wire n185011;
   wire n185012;
   wire n185013;
   wire n185014;
   wire n185015;
   wire n185016;
   wire n185017;
   wire n185018;
   wire n185019;
   wire n185020;
   wire n185021;
   wire n185022;
   wire n185023;
   wire n185024;
   wire n185025;
   wire n185026;
   wire n185027;
   wire n185028;
   wire n185029;
   wire n185030;
   wire n185031;
   wire n185032;
   wire n185033;
   wire n185034;
   wire n185035;
   wire n185036;
   wire n185037;
   wire n185038;
   wire n185039;
   wire n185040;
   wire n185041;
   wire n185042;
   wire n185043;
   wire n185044;
   wire n185045;
   wire n185046;
   wire n185047;
   wire n185048;
   wire n185049;
   wire n185050;
   wire n185051;
   wire n185052;
   wire n185053;
   wire n185054;
   wire n185055;
   wire n185056;
   wire n185057;
   wire n185058;
   wire n185059;
   wire n185060;
   wire n185061;
   wire n185062;
   wire n185063;
   wire n185064;
   wire n185065;
   wire n185066;
   wire n185067;
   wire n185068;
   wire n185069;
   wire n185070;
   wire n185071;
   wire n185072;
   wire n185073;
   wire n185074;
   wire n185075;
   wire n185076;
   wire n185077;
   wire n185078;
   wire n185079;
   wire n185080;
   wire n185081;
   wire n185082;
   wire n185083;
   wire n185084;
   wire n185085;
   wire n185086;
   wire n185087;
   wire n185088;
   wire n185089;
   wire n185090;
   wire n185091;
   wire n185092;
   wire n185093;
   wire n185094;
   wire n185095;
   wire n185096;
   wire n185097;
   wire n185098;
   wire n185099;
   wire n185100;
   wire n185101;
   wire n185102;
   wire n185103;
   wire n185104;
   wire n185105;
   wire n185106;
   wire n185107;
   wire n185108;
   wire n185109;
   wire n185110;
   wire n185111;
   wire n185112;
   wire n185113;
   wire n185114;
   wire n185115;
   wire n185116;
   wire n185117;
   wire n185118;
   wire n185119;
   wire n185120;
   wire n185121;
   wire n185122;
   wire n185123;
   wire n185124;
   wire n185125;
   wire n185126;
   wire n185127;
   wire n185128;
   wire n185129;
   wire n185130;
   wire n185131;
   wire n185132;
   wire n185133;
   wire n185134;
   wire n185135;
   wire n185136;
   wire n185137;
   wire n185138;
   wire n185139;
   wire n185140;
   wire n185141;
   wire n185142;
   wire n185143;
   wire n185144;
   wire n185145;
   wire n185146;
   wire n185147;
   wire n185148;
   wire n185149;
   wire n185150;
   wire n185151;
   wire n185152;
   wire n185153;
   wire n185154;
   wire n185155;
   wire n185156;
   wire n185157;
   wire n185158;
   wire n185159;
   wire n185160;
   wire n185161;
   wire n185162;
   wire n185163;
   wire n185164;
   wire n185165;
   wire n185166;
   wire n185167;
   wire n185168;
   wire n185169;
   wire n185170;
   wire n185171;
   wire n185172;
   wire n185173;
   wire n185174;
   wire n185175;
   wire n185176;
   wire n185177;
   wire n185178;
   wire n185179;
   wire n185180;
   wire n185181;
   wire n185182;
   wire n185183;
   wire n185184;
   wire n185185;
   wire n185186;
   wire n185187;
   wire n185188;
   wire n185189;
   wire n185190;
   wire n185191;
   wire n185192;
   wire n185193;
   wire n185194;
   wire n185195;
   wire n185196;
   wire n185197;
   wire n185198;
   wire n185199;
   wire n185200;
   wire n185201;
   wire n185202;
   wire n185203;
   wire n185204;
   wire n185205;
   wire n185206;
   wire n185207;
   wire n185208;
   wire n185209;
   wire n185210;
   wire n185211;
   wire n185212;
   wire n185213;
   wire n185214;
   wire n185215;
   wire n185216;
   wire n185217;
   wire n185218;
   wire n185219;
   wire n185220;
   wire n185221;
   wire n185222;
   wire n185223;
   wire n185224;
   wire n185225;
   wire n185226;
   wire n185227;
   wire n185228;
   wire n185229;
   wire n185230;
   wire n185231;
   wire n185232;
   wire n185233;
   wire n185234;
   wire n185235;
   wire n185236;
   wire n185237;
   wire n185238;
   wire n185239;
   wire n185240;
   wire n185241;
   wire n185242;
   wire n185243;
   wire n185244;
   wire n185245;
   wire n185246;
   wire n185247;
   wire n185248;
   wire n185249;
   wire n185250;
   wire n185251;
   wire n185252;
   wire n185253;
   wire n185254;
   wire n185255;
   wire n185256;
   wire n185257;
   wire n185258;
   wire n185259;
   wire n185260;
   wire n185261;
   wire n185262;
   wire n185263;
   wire n185264;
   wire n185265;
   wire n185266;
   wire n185267;
   wire n185268;
   wire n185269;
   wire n185270;
   wire n185271;
   wire n185272;
   wire n185273;
   wire n185274;
   wire n185275;
   wire n185276;
   wire n185277;
   wire n185278;
   wire n185279;
   wire n185280;
   wire n185281;
   wire n185282;
   wire n185283;
   wire n185284;
   wire n185285;
   wire n185286;
   wire n185287;
   wire n185288;
   wire n185289;
   wire n185290;
   wire n185291;
   wire n185292;
   wire n185293;
   wire n185294;
   wire n185295;
   wire n185296;
   wire n185297;
   wire n185298;
   wire n185299;
   wire n185300;
   wire n185301;
   wire n185302;
   wire n185303;
   wire n185304;
   wire n185305;
   wire n185306;
   wire n185307;
   wire n185308;
   wire n185309;
   wire n185310;
   wire n185311;
   wire n185312;
   wire n185313;
   wire n185314;
   wire n185315;
   wire n185316;
   wire n185317;
   wire n185318;
   wire n185319;
   wire n185320;
   wire n185321;
   wire n185322;
   wire n185323;
   wire n185324;
   wire n185325;
   wire n185326;
   wire n185327;
   wire n185328;
   wire n185329;
   wire n185330;
   wire n185331;
   wire n185332;
   wire n185333;
   wire n185334;
   wire n185335;
   wire n185336;
   wire n185337;
   wire n185338;
   wire n185339;
   wire n185340;
   wire n185341;
   wire n185342;
   wire n185343;
   wire n185344;
   wire n185345;
   wire n185346;
   wire n185347;
   wire n185348;
   wire n185349;
   wire n185350;
   wire n185351;
   wire n185352;
   wire n185353;
   wire n185354;
   wire n185355;
   wire n185356;
   wire n185357;
   wire n185358;
   wire n185359;
   wire n185360;
   wire n185361;
   wire n185362;
   wire n185363;
   wire n185364;
   wire n185365;
   wire n185366;
   wire n185367;
   wire n185368;
   wire n185369;
   wire n185370;
   wire n185371;
   wire n185372;
   wire n185373;
   wire n185374;
   wire n185375;
   wire n185376;
   wire n185377;
   wire n185378;
   wire n185379;
   wire n185380;
   wire n185381;
   wire n185382;
   wire n185383;
   wire n185384;
   wire n185385;
   wire n185386;
   wire n185387;
   wire n185388;
   wire n185389;
   wire n185390;
   wire n185391;
   wire n185392;
   wire n185393;
   wire n185394;
   wire n185395;
   wire n185396;
   wire n185397;
   wire n185398;
   wire n185399;
   wire n185400;
   wire n185401;
   wire n185402;
   wire n185403;
   wire n185404;
   wire n185405;
   wire n185406;
   wire n185407;
   wire n185408;
   wire n185409;
   wire n185410;
   wire n185411;
   wire n185412;
   wire n185413;
   wire n185414;
   wire n185415;
   wire n185416;
   wire n185417;
   wire n185418;
   wire n185419;
   wire n185420;
   wire n185421;
   wire n185422;
   wire n185423;
   wire n185424;
   wire n185425;
   wire n185426;
   wire n185427;
   wire n185428;
   wire n185429;
   wire n185430;
   wire n185431;
   wire n185432;
   wire n185433;
   wire n185434;
   wire n185435;
   wire n185436;
   wire n185437;
   wire n185438;
   wire n185439;
   wire n185440;
   wire n185441;
   wire n185442;
   wire n185443;
   wire n185444;
   wire n185445;
   wire n185446;
   wire n185447;
   wire n185448;
   wire n185449;
   wire n185450;
   wire n185451;
   wire n185452;
   wire n185453;
   wire n185454;
   wire n185455;
   wire n185456;
   wire n185457;
   wire n185458;
   wire n185459;
   wire n185460;
   wire n185461;
   wire n185462;
   wire n185463;
   wire n185464;
   wire n185465;
   wire n185466;
   wire n185467;
   wire n185468;
   wire n185469;
   wire n185470;
   wire n185471;
   wire n185472;
   wire n185473;
   wire n185474;
   wire n185475;
   wire n185476;
   wire n185477;
   wire n185478;
   wire n185479;
   wire n185480;
   wire n185481;
   wire n185482;
   wire n185483;
   wire n185484;
   wire n185485;
   wire n185486;
   wire n185487;
   wire n185488;
   wire n185489;
   wire n185490;
   wire n185491;
   wire n185492;
   wire n185493;
   wire n185494;
   wire n185495;
   wire n185496;
   wire n185497;
   wire n185498;
   wire n185499;
   wire n185500;
   wire n185501;
   wire n185502;
   wire n185503;
   wire n185504;
   wire n185505;
   wire n185506;
   wire n185507;
   wire n185508;
   wire n185509;
   wire n185510;
   wire n185511;
   wire n185512;
   wire n185513;
   wire n185514;
   wire n185515;
   wire n185516;
   wire n185517;
   wire n185518;
   wire n185519;
   wire n185520;
   wire n185521;
   wire n185522;
   wire n185523;
   wire n185524;
   wire n185525;
   wire n185526;
   wire n185527;
   wire n185528;
   wire n185529;
   wire n185530;
   wire n185531;
   wire n185532;
   wire n185533;
   wire n185534;
   wire n185535;
   wire n185536;
   wire n185537;
   wire n185538;
   wire n185539;
   wire n185540;
   wire n185541;
   wire n185542;
   wire n185543;
   wire n185544;
   wire n185545;
   wire n185546;
   wire n185547;
   wire n185548;
   wire n185549;
   wire n185550;
   wire n185551;
   wire n185552;
   wire n185553;
   wire n185554;
   wire n185555;
   wire n185556;
   wire n185557;
   wire n185558;
   wire n185559;
   wire n185560;
   wire n185561;
   wire n185562;
   wire n185563;
   wire n185564;
   wire n185565;
   wire n185566;
   wire n185567;
   wire n185568;
   wire n185569;
   wire n185570;
   wire n185571;
   wire n185572;
   wire n185573;
   wire n185574;
   wire n185575;
   wire n185576;
   wire n185577;
   wire n185578;
   wire n185579;
   wire n185580;
   wire n185581;
   wire n185582;
   wire n185583;
   wire n185584;
   wire n185585;
   wire n185586;
   wire n185587;
   wire n185588;
   wire n185589;
   wire n185590;
   wire n185591;
   wire n185592;
   wire n185593;
   wire n185594;
   wire n185595;
   wire n185596;
   wire n185597;
   wire n185598;
   wire n185599;
   wire n185600;
   wire n185601;
   wire n185602;
   wire n185603;
   wire n185604;
   wire n185605;
   wire n185606;
   wire n185607;
   wire n185608;
   wire n185609;
   wire n185610;
   wire n185611;
   wire n185612;
   wire n185613;
   wire n185614;
   wire n185615;
   wire n185616;
   wire n185617;
   wire n185618;
   wire n185619;
   wire n185620;
   wire n185621;
   wire n185622;
   wire n185623;
   wire n185624;
   wire n185625;
   wire n185626;
   wire n185627;
   wire n185628;
   wire n185629;
   wire n185630;
   wire n185631;
   wire n185632;
   wire n185633;
   wire n185634;
   wire n185635;
   wire n185636;
   wire n185637;
   wire n185638;
   wire n185639;
   wire n185640;
   wire n185641;
   wire n185642;
   wire n185643;
   wire n185644;
   wire n185645;
   wire n185646;
   wire n185647;
   wire n185648;
   wire n185649;
   wire n185650;
   wire n185651;
   wire n185652;
   wire n185653;
   wire n185654;
   wire n185655;
   wire n185656;
   wire n185657;
   wire n185658;
   wire n185659;
   wire n185660;
   wire n185661;
   wire n185662;
   wire n185663;
   wire n185664;
   wire n185665;
   wire n185666;
   wire n185667;
   wire n185668;
   wire n185669;
   wire n185670;
   wire n185671;
   wire n185672;
   wire n185673;
   wire n185674;
   wire n185675;
   wire n185676;
   wire n185677;
   wire n185678;
   wire n185679;
   wire n185680;
   wire n185681;
   wire n185682;
   wire n185683;
   wire n185684;
   wire n185685;
   wire n185686;
   wire n185687;
   wire n185688;
   wire n185689;
   wire n185690;
   wire n185691;
   wire n185692;
   wire n185693;
   wire n185694;
   wire n185695;
   wire n185696;
   wire n185697;
   wire n185698;
   wire n185699;
   wire n185700;
   wire n185701;
   wire n185702;
   wire n185703;
   wire n185704;
   wire n185705;
   wire n185706;
   wire n185707;
   wire n185708;
   wire n185709;
   wire n185710;
   wire n185711;
   wire n185712;
   wire n185713;
   wire n185714;
   wire n185715;
   wire n185716;
   wire n185717;
   wire n185718;
   wire n185719;
   wire n185720;
   wire n185721;
   wire n185722;
   wire n185723;
   wire n185724;
   wire n185725;
   wire n185726;
   wire n185727;
   wire n185728;
   wire n185729;
   wire n185730;
   wire n185731;
   wire n185732;
   wire n185733;
   wire n185734;
   wire n185735;
   wire n185736;
   wire n185737;
   wire n185738;
   wire n185739;
   wire n185740;
   wire n185741;
   wire n185742;
   wire n185743;
   wire n185744;
   wire n185745;
   wire n185746;
   wire n185747;
   wire n185748;
   wire n185749;
   wire n185750;
   wire n185751;
   wire n185752;
   wire n185753;
   wire n185754;
   wire n185755;
   wire n185756;
   wire n185757;
   wire n185758;
   wire n185759;
   wire n185760;
   wire n185761;
   wire n185762;
   wire n185763;
   wire n185764;
   wire n185765;
   wire n185766;
   wire n185767;
   wire n185768;
   wire n185769;
   wire n185770;
   wire n185771;
   wire n185772;
   wire n185773;
   wire n185774;
   wire n185775;
   wire n185776;
   wire n185777;
   wire n185778;
   wire n185779;
   wire n185780;
   wire n185781;
   wire n185782;
   wire n185783;
   wire n185784;
   wire n185785;
   wire n185786;
   wire n185787;
   wire n185788;
   wire n185789;
   wire n185790;
   wire n185791;
   wire n185792;
   wire n185793;
   wire n185794;
   wire n185795;
   wire n185796;
   wire n185797;
   wire n185798;
   wire n185799;
   wire n185800;
   wire n185801;
   wire n185802;
   wire n185803;
   wire n185804;
   wire n185805;
   wire n185806;
   wire n185807;
   wire n185808;
   wire n185809;
   wire n185810;
   wire n185811;
   wire n185812;
   wire n185813;
   wire n185814;
   wire n185815;
   wire n185816;
   wire n185817;
   wire n185818;
   wire n185819;
   wire n185820;
   wire n185821;
   wire n185822;
   wire n185823;
   wire n185824;
   wire n185825;
   wire n185826;
   wire n185827;
   wire n185828;
   wire n185829;
   wire n185830;
   wire n185831;
   wire n185832;
   wire n185833;
   wire n185834;
   wire n185835;
   wire n185836;
   wire n185837;
   wire n185838;
   wire n185839;
   wire n185840;
   wire n185841;
   wire n185842;
   wire n185843;
   wire n185844;
   wire n185845;
   wire n185846;
   wire n185847;
   wire n185848;
   wire n185849;
   wire n185850;
   wire n185851;
   wire n185852;
   wire n185853;
   wire n185854;
   wire n185855;
   wire n185856;
   wire n185857;
   wire n185858;
   wire n185859;
   wire n185860;
   wire n185861;
   wire n185862;
   wire n185863;
   wire n185864;
   wire n185865;
   wire n185866;
   wire n185867;
   wire n185868;
   wire n185869;
   wire n185870;
   wire n185871;
   wire n185872;
   wire n185873;
   wire n185874;
   wire n185875;
   wire n185876;
   wire n185877;
   wire n185878;
   wire n185879;
   wire n185880;
   wire n185881;
   wire n185882;
   wire n185883;
   wire n185884;
   wire n185885;
   wire n185886;
   wire n185887;
   wire n185888;
   wire n185889;
   wire n185890;
   wire n185891;
   wire n185892;
   wire n185893;
   wire n185894;
   wire n185895;
   wire n185896;
   wire n185897;
   wire n185898;
   wire n185899;
   wire n185900;
   wire n185901;
   wire n185902;
   wire n185903;
   wire n185904;
   wire n185905;
   wire n185906;
   wire n185907;
   wire n185908;
   wire n185909;
   wire n185910;
   wire n185911;
   wire n185912;
   wire n185913;
   wire n185914;
   wire n185915;
   wire n185916;
   wire n185917;
   wire n185918;
   wire n185919;
   wire n185920;
   wire n185921;
   wire n185922;
   wire n185923;
   wire n185924;
   wire n185925;
   wire n185926;
   wire n185927;
   wire n185928;
   wire n185929;
   wire n185930;
   wire n185931;
   wire n185932;
   wire n185933;
   wire n185934;
   wire n185935;
   wire n185936;
   wire n185937;
   wire n185938;
   wire n185939;
   wire n185940;
   wire n185941;
   wire n185942;
   wire n185943;
   wire n185944;
   wire n185945;
   wire n185946;
   wire n185947;
   wire n185948;
   wire n185949;
   wire n185950;
   wire n185951;
   wire n185952;
   wire n185953;
   wire n185954;
   wire n185955;
   wire n185956;
   wire n185957;
   wire n185958;
   wire n185959;
   wire n185960;
   wire n185961;
   wire n185962;
   wire n185963;
   wire n185964;
   wire n185965;
   wire n185966;
   wire n185967;
   wire n185968;
   wire n185969;
   wire n185970;
   wire n185971;
   wire n185972;
   wire n185973;
   wire n185974;
   wire n185975;
   wire n185976;
   wire n185977;
   wire n185978;
   wire n185979;
   wire n185980;
   wire n185981;
   wire n185982;
   wire n185983;
   wire n185984;
   wire n185985;
   wire n185986;
   wire n185987;
   wire n185988;
   wire n185989;
   wire n185990;
   wire n185991;
   wire n185992;
   wire n185993;
   wire n185994;
   wire n185995;
   wire n185996;
   wire n185997;
   wire n185998;
   wire n185999;
   wire n186000;
   wire n186001;
   wire n186002;
   wire n186003;
   wire n186004;
   wire n186005;
   wire n186006;
   wire n186007;
   wire n186008;
   wire n186009;
   wire n186010;
   wire n186011;
   wire n186012;
   wire n186013;
   wire n186014;
   wire n186015;
   wire n186016;
   wire n186017;
   wire n186018;
   wire n186019;
   wire n186020;
   wire n186021;
   wire n186022;
   wire n186023;
   wire n186024;
   wire n186025;
   wire n186026;
   wire n186027;
   wire n186028;
   wire n186029;
   wire n186030;
   wire n186031;
   wire n186032;
   wire n186033;
   wire n186034;
   wire n186035;
   wire n186036;
   wire n186037;
   wire n186038;
   wire n186039;
   wire n186040;
   wire n186041;
   wire n186042;
   wire n186043;
   wire n186044;
   wire n186045;
   wire n186046;
   wire n186047;
   wire n186048;
   wire n186049;
   wire n186050;
   wire n186051;
   wire n186052;
   wire n186053;
   wire n186054;
   wire n186055;
   wire n186056;
   wire n186057;
   wire n186058;
   wire n186059;
   wire n186060;
   wire n186061;
   wire n186062;
   wire n186063;
   wire n186064;
   wire n186065;
   wire n186066;
   wire n186067;
   wire n186068;
   wire n186069;
   wire n186070;
   wire n186071;
   wire n186072;
   wire n186073;
   wire n186074;
   wire n186075;
   wire n186076;
   wire n186077;
   wire n186078;
   wire n186079;
   wire n186080;
   wire n186081;
   wire n186082;
   wire n186083;
   wire n186084;
   wire n186085;
   wire n186086;
   wire n186087;
   wire n186088;
   wire n186089;
   wire n186090;
   wire n186091;
   wire n186092;
   wire n186093;
   wire n186094;
   wire n186095;
   wire n186096;
   wire n186097;
   wire n186098;
   wire n186099;
   wire n186100;
   wire n186101;
   wire n186102;
   wire n186103;
   wire n186104;
   wire n186105;
   wire n186106;
   wire n186107;
   wire n186108;
   wire n186109;
   wire n186110;
   wire n186111;
   wire n186112;
   wire n186113;
   wire n186114;
   wire n186115;
   wire n186116;
   wire n186117;
   wire n186118;
   wire n186119;
   wire n186120;
   wire n186121;
   wire n186122;
   wire n186123;
   wire n186124;
   wire n186125;
   wire n186126;
   wire n186127;
   wire n186128;
   wire n186129;
   wire n186130;
   wire n186131;
   wire n186132;
   wire n186133;
   wire n186134;
   wire n186135;
   wire n186136;
   wire n186137;
   wire n186138;
   wire n186139;
   wire n186140;
   wire n186141;
   wire n186142;
   wire n186143;
   wire n186144;
   wire n186145;
   wire n186146;
   wire n186147;
   wire n186148;
   wire n186149;
   wire n186150;
   wire n186151;
   wire n186152;
   wire n186153;
   wire n186154;
   wire n186155;
   wire n186156;
   wire n186157;
   wire n186158;
   wire n186159;
   wire n186160;
   wire n186161;
   wire n186162;
   wire n186163;
   wire n186164;
   wire n186165;
   wire n186166;
   wire n186167;
   wire n186168;
   wire n186169;
   wire n186170;
   wire n186171;
   wire n186172;
   wire n186173;
   wire n186174;
   wire n186175;
   wire n186176;
   wire n186177;
   wire n186178;
   wire n186179;
   wire n186180;
   wire n186181;
   wire n186182;
   wire n186183;
   wire n186184;
   wire n186185;
   wire n186186;
   wire n186187;
   wire n186188;
   wire n186189;
   wire n186190;
   wire n186191;
   wire n186192;
   wire n186193;
   wire n186194;
   wire n186195;
   wire n186196;
   wire n186197;
   wire n186198;
   wire n186199;
   wire n186200;
   wire n186201;
   wire n186202;
   wire n186203;
   wire n186204;
   wire n186205;
   wire n186206;
   wire n186207;
   wire n186208;
   wire n186209;
   wire n186210;
   wire n186211;
   wire n186212;
   wire n186213;
   wire n186214;
   wire n186215;
   wire n186216;
   wire n186217;
   wire n186218;
   wire n186219;
   wire n186220;
   wire n186221;
   wire n186222;
   wire n186223;
   wire n186224;
   wire n186225;
   wire n186226;
   wire n186227;
   wire n186228;
   wire n186229;
   wire n186230;
   wire n186231;
   wire n186232;
   wire n186233;
   wire n186234;
   wire n186235;
   wire n186236;
   wire n186237;
   wire n186238;
   wire n186239;
   wire n186240;
   wire n186241;
   wire n186242;
   wire n186243;
   wire n186244;
   wire n186245;
   wire n186246;
   wire n186247;
   wire n186248;
   wire n186249;
   wire n186250;
   wire n186251;
   wire n186252;
   wire n186253;
   wire n186254;
   wire n186255;
   wire n186256;
   wire n186257;
   wire n186258;
   wire n186259;
   wire n186260;
   wire n186261;
   wire n186262;
   wire n186263;
   wire n186264;
   wire n186265;
   wire n186266;
   wire n186267;
   wire n186268;
   wire n186269;
   wire n186270;
   wire n186271;
   wire n186272;
   wire n186273;
   wire n186274;
   wire n186275;
   wire n186276;
   wire n186277;
   wire n186278;
   wire n186279;
   wire n186280;
   wire n186281;
   wire n186282;
   wire n186283;
   wire n186284;
   wire n186285;
   wire n186286;
   wire n186287;
   wire n186288;
   wire n186289;
   wire n186290;
   wire n186291;
   wire n186292;
   wire n186293;
   wire n186294;
   wire n186295;
   wire n186296;
   wire n186297;
   wire n186298;
   wire n186299;
   wire n186300;
   wire n186301;
   wire n186302;
   wire n186303;
   wire n186304;
   wire n186305;
   wire n186306;
   wire n186307;
   wire n186308;
   wire n186309;
   wire n186310;
   wire n186311;
   wire n186312;
   wire n186313;
   wire n186314;
   wire n186315;
   wire n186316;
   wire n186317;
   wire n186318;
   wire n186319;
   wire n186320;
   wire n186321;
   wire n186322;
   wire n186323;
   wire n186324;
   wire n186325;
   wire n186326;
   wire n186327;
   wire n186328;
   wire n186329;
   wire n186330;
   wire n186331;
   wire n186332;
   wire n186333;
   wire n186334;
   wire n186335;
   wire n186336;
   wire n186337;
   wire n186338;
   wire n186339;
   wire n186340;
   wire n186341;
   wire n186342;
   wire n186343;
   wire n186344;
   wire n186345;
   wire n186346;
   wire n186347;
   wire n186348;
   wire n186349;
   wire n186350;
   wire n186351;
   wire n186352;
   wire n186353;
   wire n186354;
   wire n186355;
   wire n186356;
   wire n186357;
   wire n186358;
   wire n186359;
   wire n186360;
   wire n186361;
   wire n186362;
   wire n186363;
   wire n186364;
   wire n186365;
   wire n186366;
   wire n186367;
   wire n186368;
   wire n186369;
   wire n186370;
   wire n186371;
   wire n186372;
   wire n186373;
   wire n186374;
   wire n186375;
   wire n186376;
   wire n186377;
   wire n186378;
   wire n186379;
   wire n186380;
   wire n186381;
   wire n186382;
   wire n186383;
   wire n186384;
   wire n186385;
   wire n186386;
   wire n186387;
   wire n186388;
   wire n186389;
   wire n186390;
   wire n186391;
   wire n186392;
   wire n186393;
   wire n186394;
   wire n186395;
   wire n186396;
   wire n186397;
   wire n186398;
   wire n186399;
   wire n186400;
   wire n186401;
   wire n186402;
   wire n186403;
   wire n186404;
   wire n186405;
   wire n186406;
   wire n186407;
   wire n186408;
   wire n186409;
   wire n186410;
   wire n186411;
   wire n186412;
   wire n186413;
   wire n186414;
   wire n186415;
   wire n186416;
   wire n186417;
   wire n186418;
   wire n186419;
   wire n186420;
   wire n186421;
   wire n186422;
   wire n186423;
   wire n186424;
   wire n186425;
   wire n186426;
   wire n186427;
   wire n186428;
   wire n186429;
   wire n186430;
   wire n186431;
   wire n186432;
   wire n186433;
   wire n186434;
   wire n186435;
   wire n186436;
   wire n186437;
   wire n186438;
   wire n186439;
   wire n186440;
   wire n186441;
   wire n186442;
   wire n186443;
   wire n186444;
   wire n186445;
   wire n186446;
   wire n186447;
   wire n186448;
   wire n186449;
   wire n186450;
   wire n186451;
   wire n186452;
   wire n186453;
   wire n186454;
   wire n186455;
   wire n186456;
   wire n186457;
   wire n186458;
   wire n186459;
   wire n186460;
   wire n186461;
   wire n186462;
   wire n186463;
   wire n186464;
   wire n186465;
   wire n186466;
   wire n186467;
   wire n186468;
   wire n186469;
   wire n186470;
   wire n186471;
   wire n186472;
   wire n186473;
   wire n186474;
   wire n186475;
   wire n186476;
   wire n186477;
   wire n186478;
   wire n186479;
   wire n186480;
   wire n186481;
   wire n186482;
   wire n186483;
   wire n186484;
   wire n186485;
   wire n186486;
   wire n186487;
   wire n186488;
   wire n186489;
   wire n186490;
   wire n186491;
   wire n186492;
   wire n186493;
   wire n186494;
   wire n186495;
   wire n186496;
   wire n186497;
   wire n186498;
   wire n186499;
   wire n186500;
   wire n186501;
   wire n186502;
   wire n186503;
   wire n186504;
   wire n186505;
   wire n186506;
   wire n186507;
   wire n186508;
   wire n186509;
   wire n186510;
   wire n186511;
   wire n186512;
   wire n186513;
   wire n186514;
   wire n186515;
   wire n186516;
   wire n186517;
   wire n186518;
   wire n186519;
   wire n186520;
   wire n186521;
   wire n186522;
   wire n186523;
   wire n186524;
   wire n186525;
   wire n186526;
   wire n186527;
   wire n186528;
   wire n186529;
   wire n186530;
   wire n186531;
   wire n186532;
   wire n186533;
   wire n186534;
   wire n186535;
   wire n186536;
   wire n186537;
   wire n186538;
   wire n186539;
   wire n186540;
   wire n186541;
   wire n186542;
   wire n186543;
   wire n186544;
   wire n186545;
   wire n186546;
   wire n186547;
   wire n186548;
   wire n186549;
   wire n186550;
   wire n186551;
   wire n186552;
   wire n186553;
   wire n186554;
   wire n186555;
   wire n186556;
   wire n186557;
   wire n186558;
   wire n186559;
   wire n186560;
   wire n186561;
   wire n186562;
   wire n186563;
   wire n186564;
   wire n186565;
   wire n186566;
   wire n186567;
   wire n186568;
   wire n186569;
   wire n186570;
   wire n186571;
   wire n186572;
   wire n186573;
   wire n186574;
   wire n186575;
   wire n186576;
   wire n186577;
   wire n186578;
   wire n186579;
   wire n186580;
   wire n186581;
   wire n186582;
   wire n186583;
   wire n186584;
   wire n186585;
   wire n186586;
   wire n186587;
   wire n186588;
   wire n186589;
   wire n186590;
   wire n186591;
   wire n186592;
   wire n186593;
   wire n186594;
   wire n186595;
   wire n186596;
   wire n186597;
   wire n186598;
   wire n186599;
   wire n186600;
   wire n186601;
   wire n186602;
   wire n186603;
   wire n186604;
   wire n186605;
   wire n186606;
   wire n186607;
   wire n186608;
   wire n186609;
   wire n186610;
   wire n186611;
   wire n186612;
   wire n186613;
   wire n186614;
   wire n186615;
   wire n186616;
   wire n186617;
   wire n186618;
   wire n186619;
   wire n186620;
   wire n186621;
   wire n186622;
   wire n186623;
   wire n186624;
   wire n186625;
   wire n186626;
   wire n186627;
   wire n186628;
   wire n186629;
   wire n186630;
   wire n186631;
   wire n186632;
   wire n186633;
   wire n186634;
   wire n186635;
   wire n186636;
   wire n186637;
   wire n186638;
   wire n186639;
   wire n186640;
   wire n186641;
   wire n186642;
   wire n186643;
   wire n186644;
   wire n186645;
   wire n186646;
   wire n186647;
   wire n186648;
   wire n186649;
   wire n186650;
   wire n186651;
   wire n186652;
   wire n186653;
   wire n186654;
   wire n186655;
   wire n186656;
   wire n186657;
   wire n186658;
   wire n186659;
   wire n186660;
   wire n186661;
   wire n186662;
   wire n186663;
   wire n186664;
   wire n186665;
   wire n186666;
   wire n186667;
   wire n186668;
   wire n186669;
   wire n186670;
   wire n186671;
   wire n186672;
   wire n186673;
   wire n186674;
   wire n186675;
   wire n186676;
   wire n186677;
   wire n186678;
   wire n186679;
   wire n186680;
   wire n186681;
   wire n186682;
   wire n186684;
   wire n186685;
   wire n186686;
   wire n186687;
   wire n186688;
   wire n186689;
   wire n186690;
   wire n186691;
   wire n186692;
   wire n186693;
   wire n186694;
   wire n186695;
   wire n186696;
   wire n186697;
   wire n186698;
   wire n186699;
   wire n186713;
   wire n186714;
   wire n186717;
   wire n186718;
   wire n186720;
   wire n186721;
   wire n186722;
   wire n186723;
   wire n186724;
   wire n186725;
   wire n186726;
   wire n186732;
   wire n211876;
   wire n211877;
   wire n211878;
   wire n211879;
   wire n211880;
   wire n211881;
   wire n211882;
   wire n211883;
   wire n211884;
   wire n211885;
   wire n211886;
   wire n211887;
   wire n211888;
   wire n211889;
   wire n211890;
   wire n211891;
   wire n211892;
   wire n211893;
   wire n211894;
   wire n211895;
   wire n211896;
   wire n211897;
   wire n211898;
   wire n211899;
   wire n211900;
   wire n211901;
   wire n211902;
   wire n211903;
   wire n211904;
   wire n211905;
   wire n211906;
   wire n211907;
   wire n211908;
   wire n211909;
   wire n211910;
   wire n211911;
   wire n211912;
   wire n211913;
   wire n211914;
   wire n211915;
   wire n211916;
   wire n211917;
   wire n211918;
   wire n211919;
   wire n211920;
   wire n211921;
   wire n211922;
   wire n211923;
   wire n211924;
   wire n211925;
   wire n211926;
   wire n211927;
   wire n211928;
   wire n211929;
   wire n211930;
   wire n211931;
   wire n211932;
   wire n211933;
   wire n211934;
   wire n211935;
   wire n211936;
   wire n211937;
   wire n211938;
   wire n211939;
   wire n211940;
   wire n211948;
   wire n211949;
   wire n211950;
   wire n211951;
   wire n211952;
   wire n211953;
   wire n211954;
   wire n211955;
   wire n211956;
   wire n211957;
   wire n211958;
   wire n211959;
   wire n211960;
   wire n211961;
   wire n211962;
   wire n211963;
   wire n211964;
   wire n211965;
   wire n211966;
   wire n211967;
   wire n211968;
   wire n211969;
   wire n211970;
   wire n211971;
   wire n211972;
   wire n211973;
   wire n211974;
   wire n211975;
   wire n211976;
   wire n211977;
   wire n211978;
   wire n211979;
   wire n211980;
   wire n211981;
   wire n211982;
   wire n211983;
   wire n211984;
   wire n211985;
   wire n211986;
   wire n211987;
   wire n211988;
   wire n211989;
   wire n211990;
   wire n211991;
   wire n211992;
   wire n211993;
   wire n211994;
   wire n211995;
   wire n211996;
   wire n211997;
   wire n211998;
   wire n211999;
   wire n212000;
   wire n212001;
   wire n212002;
   wire n212003;
   wire n212004;
   wire n212005;
   wire n212006;
   wire n212007;
   wire n212008;
   wire n212009;
   wire n212010;
   wire n212011;
   wire n212012;
   wire n212013;
   wire n212014;
   wire n212015;
   wire n212016;
   wire n212017;
   wire n212018;
   wire n212019;
   wire n212020;
   wire n212021;
   wire n212022;
   wire n212023;
   wire n212024;
   wire n212025;
   wire n212026;
   wire n212027;
   wire n212028;
   wire n212029;
   wire n212030;
   wire n212031;
   wire n212032;
   wire n212033;
   wire n212034;
   wire n212035;
   wire n212036;
   wire n212037;
   wire n212038;
   wire n212039;
   wire n212040;
   wire n212041;
   wire n212042;
   wire n212043;
   wire n212044;
   wire n212045;
   wire n212046;
   wire n212047;
   wire n212048;
   wire n212049;
   wire n212050;
   wire n212051;
   wire n212052;
   wire n212053;
   wire n212054;
   wire n212055;
   wire n212056;
   wire n212057;
   wire n212058;
   wire n212059;
   wire n212060;
   wire n212061;
   wire n212062;
   wire n212063;
   wire n212064;
   wire n212065;
   wire n212066;
   wire n212067;
   wire n212068;
   wire n212069;
   wire n212070;
   wire n212071;
   wire n212072;
   wire n212073;
   wire n212074;
   wire n212075;
   wire n212076;
   wire n212077;
   wire n212078;
   wire n212079;
   wire n212080;
   wire n212081;
   wire n212082;
   wire n212083;
   wire n212084;
   wire n212085;
   wire n212086;
   wire n212087;
   wire n212088;
   wire n212089;
   wire n212090;
   wire n212091;
   wire n212092;
   wire n212093;
   wire n212094;
   wire n212095;
   wire n212096;
   wire n212097;
   wire n212098;
   wire n212099;
   wire n212100;
   wire n212101;
   wire n212102;
   wire n212103;
   wire n212104;
   wire n212105;
   wire n212106;
   wire n212107;
   wire n212108;
   wire n212109;
   wire n212110;
   wire n212111;
   wire n212112;
   wire n212113;
   wire n212114;
   wire n212115;
   wire n212116;
   wire n212117;
   wire n212118;
   wire n212119;
   wire n212120;
   wire n212121;
   wire n212122;
   wire n212123;
   wire n212124;
   wire n212125;
   wire n212126;
   wire n212127;
   wire n212128;
   wire n212129;
   wire n212130;
   wire n212131;
   wire n212132;
   wire n212133;
   wire n212134;
   wire n212135;
   wire n212136;
   wire n212137;
   wire n212138;
   wire n212139;
   wire n212140;
   wire n212141;
   wire n212142;
   wire n212143;
   wire n212144;
   wire n212145;
   wire n212146;
   wire n212147;
   wire n212148;
   wire n212149;
   wire n212150;
   wire n212151;
   wire n212152;
   wire n212153;
   wire n212154;
   wire n212155;
   wire n212156;
   wire n212157;
   wire n212158;
   wire n212159;
   wire n212160;
   wire n212161;
   wire n212162;
   wire n212163;
   wire n212164;
   wire n212165;
   wire n212166;
   wire n212167;
   wire n212168;
   wire n212169;
   wire n212170;
   wire n212171;
   wire n212172;
   wire n212173;
   wire n212174;
   wire n212175;
   wire n212176;
   wire n212177;
   wire n212178;
   wire n212179;
   wire n212180;
   wire n212181;
   wire n212182;
   wire n212183;
   wire n212184;
   wire n212185;
   wire n212186;
   wire n212187;
   wire n212188;
   wire n212189;
   wire n212190;
   wire n212191;
   wire n212192;
   wire n212193;
   wire n212194;
   wire n212195;
   wire n212196;
   wire n212197;
   wire n212198;
   wire n212199;
   wire n212200;
   wire n212201;
   wire n212202;
   wire n212203;
   wire n212204;
   wire n212205;
   wire n212206;
   wire n212207;
   wire n212208;
   wire n212209;
   wire n212210;
   wire n212211;
   wire n212212;
   wire n212213;
   wire n212214;
   wire n212215;
   wire n212216;
   wire n212217;
   wire n212218;
   wire n212219;
   wire n212220;
   wire n212221;
   wire n212222;
   wire n212223;
   wire n212224;
   wire n212225;
   wire n212226;
   wire n212227;
   wire n212228;
   wire n212229;
   wire n212230;
   wire n212231;
   wire n212232;
   wire n212233;
   wire n212234;
   wire n212235;
   wire n212236;
   wire n212237;
   wire n212238;
   wire n212239;
   wire n212240;
   wire n212241;
   wire n212242;
   wire n212243;
   wire n212244;
   wire n212245;
   wire n212246;
   wire n212247;
   wire n212248;
   wire n212249;
   wire n212250;
   wire n212251;
   wire n212252;
   wire n212253;
   wire n212254;
   wire n212255;
   wire n212256;
   wire n212257;
   wire n212258;
   wire n212259;
   wire n212260;
   wire n212261;
   wire n212262;
   wire n212263;
   wire n212264;
   wire n212265;
   wire n212266;
   wire n212267;
   wire n212268;
   wire n212269;
   wire n212270;
   wire n212271;
   wire n212272;
   wire n212273;
   wire n212274;
   wire n212275;
   wire n212276;
   wire n212277;
   wire n212278;
   wire n212279;
   wire n212280;
   wire n212281;
   wire n212282;
   wire n212283;
   wire n212284;
   wire n212285;
   wire n212286;
   wire n212287;
   wire n212289;
   wire n212290;
   wire n212291;
   wire n212292;
   wire n212415;
   wire n212416;
   wire n212423;
   wire n212425;
   wire n212463;
   wire n212465;
   wire n212486;
   wire n212487;
   wire n212488;
   wire n212533;
   wire n212534;
   wire n212535;
   wire n212536;
   wire n212537;
   wire n212538;
   wire n212539;
   wire n212540;
   wire n212541;
   wire n212542;
   wire n212543;
   wire n212544;
   wire n212545;
   wire n212546;
   wire n212547;
   wire n212548;
   wire n212549;
   wire n212550;
   wire n212551;
   wire n212552;
   wire n212553;
   wire n212554;
   wire n212555;
   wire n212556;
   wire n212557;
   wire n212558;
   wire n212559;
   wire n212560;
   wire n212561;
   wire n212562;
   wire n212571;
   wire n212572;
   wire n212573;
   wire n212574;
   wire n212576;
   wire n212577;
   wire n212578;
   wire n212579;
   wire n212582;
   wire n212584;
   wire n212586;
   wire n212588;
   wire n212590;
   wire n212592;
   wire n212594;
   wire n212596;
   wire n212598;
   wire n212600;
   wire n212602;
   wire n212604;
   wire n212606;
   wire n212608;
   wire n212610;
   wire n212612;
   wire n212614;
   wire n212616;
   wire n212618;
   wire n212620;
   wire n212622;
   wire n212624;
   wire n212626;
   wire n212628;
   wire n212630;
   wire n212632;
   wire n212634;
   wire n212636;
   wire n212638;
   wire n212640;
   wire n212642;
   wire n212644;
   wire n212677;
   wire n212678;
   wire n212679;
   wire n212680;
   wire n212681;
   wire n212682;
   wire n212683;
   wire n212684;
   wire n212685;
   wire n212686;
   wire n212687;
   wire n212688;
   wire n212689;
   wire n212690;
   wire n212691;
   wire n212692;
   wire n212693;
   wire n212694;
   wire n212695;
   wire n212696;
   wire n212697;
   wire n212698;
   wire n212699;
   wire n212700;
   wire n212701;
   wire n212702;
   wire n212703;
   wire n212704;
   wire n212705;
   wire n212706;
   wire n212707;
   wire n212708;
   wire n212709;
   wire n212710;
   wire n212711;
   wire n212712;
   wire n212713;
   wire n212714;
   wire n212715;
   wire n212716;
   wire n212717;
   wire n212718;
   wire n212719;
   wire n212720;
   wire n212721;
   wire n212722;
   wire n212723;
   wire n212724;
   wire n212725;
   wire n212726;
   wire n212727;
   wire n212728;
   wire n212729;
   wire n212730;
   wire n212731;
   wire n212732;
   wire n212733;
   wire n212734;
   wire n212735;
   wire n212736;
   wire n212737;
   wire n212738;
   wire n212739;
   wire n212740;
   wire n212741;
   wire n212742;
   wire n212743;
   wire n212744;
   wire n212745;
   wire n212746;
   wire n212747;
   wire n212748;
   wire n212749;
   wire n212750;
   wire n212751;
   wire n212752;
   wire n212753;
   wire n212754;
   wire n212755;
   wire n212756;
   wire n212757;
   wire n212758;
   wire n212759;
   wire n212760;
   wire n212761;
   wire n212762;
   wire n212763;
   wire n212764;
   wire n212765;
   wire n212766;
   wire n212767;
   wire n212768;
   wire n212769;
   wire n212770;
   wire n212771;
   wire n212772;
   wire n212773;
   wire n212774;
   wire n212775;
   wire n212776;
   wire n212777;
   wire n212778;
   wire n212779;
   wire n212780;
   wire n212781;
   wire n212782;
   wire n212783;
   wire n212784;
   wire n212785;
   wire n212786;
   wire n212787;
   wire n212788;
   wire n243096;
   wire n243097;
   wire n243163;
   wire n243166;
   wire n243167;
   wire n244213;
   wire n244214;
   wire n244215;
   wire n244216;
   wire n244217;
   wire n244218;
   wire n244219;
   wire n244220;
   wire n244221;
   wire n244222;
   wire n244245;
   wire n244250;
   wire n244262;
   wire n244263;
   wire n244964;
   wire n244965;
   wire n244966;
   wire n244967;
   wire n244968;
   wire n244969;
   wire n244970;
   wire n244971;
   wire n244972;
   wire n244973;
   wire n244974;
   wire n244975;
   wire n244976;
   wire n244977;
   wire n244978;
   wire n244979;
   wire n244980;
   wire n244981;
   wire n244982;
   wire n244983;
   wire n244984;
   wire n244985;
   wire n244986;
   wire n244987;
   wire n244988;
   wire n244989;
   wire n244990;
   wire n244991;
   wire n244992;
   wire n244994;
   wire n244995;
   wire n244996;
   wire n244997;
   wire n244998;
   wire n244999;
   wire n245000;
   wire n245001;
   wire n245002;
   wire n245003;
   wire n245004;
   wire n245005;
   wire n245006;
   wire n245007;
   wire n245008;
   wire n245009;
   wire n245010;
   wire n245011;
   wire n245012;
   wire n245013;
   wire n245014;
   wire n245015;
   wire n245016;
   wire n245017;
   wire n245018;
   wire n245019;
   wire n245020;
   wire n245021;
   wire n245022;
   wire n245023;
   wire n245024;
   wire n245025;
   wire n245026;
   wire n245083;
   wire n245090;
   wire n245091;
   wire n245109;
   wire n245110;
   wire n245111;
   wire n245314;
   wire n245315;
   wire n245316;
   wire n245317;
   wire n245318;
   wire n245319;
   wire n245320;
   wire n245321;
   wire n245322;
   wire n245323;
   wire n245324;
   wire n245325;
   wire n245326;
   wire n245327;
   wire n245328;
   wire n245329;
   wire n245330;
   wire n245331;
   wire n245332;
   wire n245333;
   wire n245334;
   wire n245335;
   wire n245336;
   wire n245337;
   wire n245338;
   wire n245339;
   wire n245340;
   wire n245341;
   wire n245342;
   wire n245343;
   wire n245344;
   wire n245345;
   wire n245346;
   wire n245347;
   wire n245348;
   wire n245349;
   wire n245350;
   wire n245351;
   wire n245352;
   wire n245353;
   wire n245354;
   wire n245355;
   wire n245356;
   wire n245357;
   wire n245358;
   wire n245359;
   wire n245360;
   wire n245361;
   wire n245362;
   wire n245363;
   wire n245364;
   wire n245365;
   wire n245366;
   wire n245367;
   wire n245368;
   wire n245369;
   wire n245370;
   wire n245371;
   wire n245372;
   wire n245373;
   wire n245374;
   wire n245375;
   wire n245376;
   wire n245377;
   wire n245378;
   wire n245379;
   wire n245380;
   wire n245381;
   wire n245382;
   wire n245383;
   wire n245384;
   wire n245385;
   wire n245386;
   wire n245387;
   wire n245388;
   wire n245389;
   wire n245390;
   wire n245391;
   wire n245392;
   wire n245393;
   wire n245394;
   wire n245395;
   wire n245396;
   wire n245397;
   wire n245398;
   wire n245399;
   wire n245400;
   wire n245401;
   wire n245402;
   wire n245403;
   wire n245404;
   wire n245405;
   wire n245406;
   wire n245407;
   wire n245408;
   wire n245409;
   wire n245410;
   wire n245411;
   wire n245412;
   wire n245413;
   wire n245414;
   wire n245415;
   wire n245416;
   wire n245417;
   wire n245418;
   wire n245419;
   wire n245420;
   wire n245421;
   wire n245422;
   wire n245423;
   wire n245424;
   wire n245425;
   wire n245426;
   wire n245427;
   wire n245428;
   wire n245429;
   wire n245430;
   wire n245431;
   wire n245432;
   wire n245433;
   wire n245434;
   wire n245435;
   wire n245436;
   wire n245437;
   wire n245438;
   wire n245439;
   wire n245440;
   wire n245441;
   wire n245442;
   wire n245443;
   wire n245444;
   wire n245445;
   wire n245446;
   wire n245447;
   wire n245448;
   wire n245449;
   wire n245450;
   wire n245451;
   wire n245452;
   wire n245453;
   wire n245454;
   wire n245455;
   wire n245456;
   wire n245457;
   wire n245458;
   wire n245459;
   wire n245460;
   wire n245461;
   wire n245462;
   wire n245463;
   wire n245464;
   wire n245465;
   wire n245466;
   wire n245467;
   wire n245468;
   wire n245469;
   wire n245470;
   wire n245471;
   wire n245472;
   wire n245473;
   wire n245474;
   wire n245475;
   wire n245476;
   wire n245477;
   wire n245478;
   wire n245479;
   wire n245480;
   wire n245481;
   wire n245483;
   wire n245484;
   wire n245485;
   wire n245486;
   wire n245487;
   wire n245488;
   wire n245490;
   wire n245491;
   wire n245492;
   wire n245493;
   wire n245494;
   wire n245495;
   wire n245496;
   wire n245497;
   wire n245498;
   wire n245499;
   wire n245500;
   wire n245501;
   wire n245502;
   wire n245503;
   wire n245504;
   wire n245505;
   wire n245506;
   wire n245507;
   wire n245508;
   wire n245509;
   wire n245510;
   wire n245511;
   wire n245512;
   wire n245513;
   wire n245514;
   wire n245515;
   wire n245516;
   wire n245517;
   wire n245518;
   wire n245519;
   wire n245520;
   wire n245521;
   wire n245522;
   wire n245523;
   wire n245524;
   wire n245525;
   wire n245526;
   wire n245527;
   wire n245528;
   wire n245529;
   wire n245530;
   wire n245531;
   wire n245532;
   wire n245533;
   wire n245534;
   wire n245535;
   wire n245536;
   wire n245537;
   wire n245538;
   wire n245539;
   wire n245540;
   wire n245541;
   wire n245542;
   wire n245543;
   wire n245544;
   wire n245545;
   wire n245546;
   wire n245547;
   wire n245548;
   wire n245549;
   wire n245550;
   wire n245551;
   wire n245552;
   wire n245553;
   wire n245554;
   wire n245555;
   wire n245556;
   wire n245557;
   wire n245558;
   wire n245559;
   wire n245560;
   wire n245561;
   wire n245562;
   wire n245563;
   wire n245564;
   wire n245565;
   wire n245566;
   wire n245567;
   wire n245568;
   wire n245569;
   wire n245570;
   wire n245571;
   wire n245572;
   wire n245573;
   wire n245574;
   wire n245575;
   wire n245576;
   wire n245577;
   wire n245578;
   wire n245579;
   wire n245580;
   wire n245581;
   wire n245582;
   wire n245583;
   wire n245584;
   wire n245585;
   wire n245586;
   wire n245587;
   wire n245588;
   wire n245589;
   wire n245590;
   wire n245591;
   wire n245592;
   wire n245593;
   wire n245594;
   wire n245595;
   wire n245596;
   wire n245597;
   wire n245598;
   wire n245599;
   wire n245600;
   wire n245601;
   wire n245602;
   wire n245603;
   wire n245604;
   wire n245605;
   wire n245606;
   wire n245607;
   wire n245608;
   wire n245609;
   wire n245610;
   wire n245611;
   wire n245612;
   wire n245613;
   wire n245614;
   wire n245615;
   wire n245616;
   wire n245617;
   wire n245618;
   wire n245619;
   wire n245620;
   wire n245621;
   wire n245622;
   wire n245623;
   wire n245624;
   wire n245625;
   wire n245626;
   wire n245627;
   wire n245628;
   wire n245629;
   wire n245630;
   wire n245631;
   wire n245632;
   wire n245633;
   wire n245634;
   wire n245635;
   wire n245636;
   wire n245637;
   wire n245638;
   wire n245639;
   wire n245640;
   wire n245641;
   wire n245642;
   wire n245643;
   wire n245644;
   wire n245645;
   wire n245646;
   wire n245647;
   wire n245648;
   wire n245649;
   wire n245650;
   wire n245651;
   wire n245652;
   wire n245653;
   wire n245654;
   wire n245655;
   wire n245656;
   wire n245657;
   wire n245658;
   wire n245659;
   wire n245660;
   wire n245661;
   wire n245662;
   wire n245663;
   wire n245664;
   wire n245665;
   wire n245666;
   wire n245667;
   wire n245668;
   wire n245669;
   wire n245670;
   wire n245671;
   wire n245672;
   wire n245673;
   wire n245674;
   wire n245675;
   wire n245676;
   wire n245677;
   wire n245678;
   wire n245679;
   wire n245680;
   wire n245681;
   wire n245682;
   wire n245683;
   wire n245684;
   wire n245685;
   wire n245686;
   wire n245687;
   wire n245688;
   wire n245689;
   wire n245690;
   wire n245691;
   wire n245692;
   wire n245693;
   wire n245694;
   wire n245695;
   wire n245696;
   wire n245697;
   wire n245698;
   wire n245699;
   wire n245700;
   wire n245701;
   wire n245702;
   wire n245703;
   wire n245704;
   wire n245705;
   wire n245706;
   wire n245707;
   wire n245708;
   wire n245709;
   wire n245710;
   wire n245711;
   wire n245712;
   wire n245713;
   wire n245714;
   wire n245715;
   wire n245716;
   wire n245717;
   wire n245718;
   wire n245719;
   wire n245720;
   wire n245721;
   wire n245722;
   wire n245723;
   wire n245724;
   wire n245725;
   wire n245726;
   wire n245727;
   wire n245728;
   wire n245729;
   wire n245730;
   wire n245731;
   wire n245732;
   wire n245733;
   wire n245734;
   wire n245735;
   wire n245736;
   wire n245737;
   wire n245738;
   wire n245739;
   wire n245740;
   wire n245741;
   wire n245742;
   wire n245743;
   wire n245744;
   wire n245745;
   wire n245746;
   wire n245747;
   wire n245748;
   wire n245749;
   wire n245750;
   wire n245751;
   wire n245752;
   wire n245753;
   wire n245754;
   wire n245755;
   wire n245756;
   wire n245757;
   wire n245758;
   wire n245759;
   wire n245760;
   wire n245761;
   wire n245762;
   wire n245763;
   wire n245764;
   wire n245765;
   wire n245766;
   wire n245767;
   wire n245768;
   wire n245769;
   wire n245770;
   wire n245771;
   wire n245772;
   wire n245773;
   wire n245774;
   wire n245775;
   wire n245776;
   wire n245777;
   wire n245778;
   wire n245779;
   wire n245780;
   wire n245781;
   wire n245782;
   wire n245783;
   wire n245784;
   wire n245785;
   wire n245786;
   wire n245787;
   wire n245788;
   wire n245789;
   wire n245790;
   wire n245791;
   wire n245792;
   wire n245793;
   wire n245794;
   wire n245795;
   wire n245796;
   wire n245797;
   wire n245798;
   wire n245799;
   wire n245800;
   wire n245801;
   wire n245802;
   wire n245803;
   wire n245804;
   wire n245805;
   wire n245806;
   wire n245807;
   wire n245808;
   wire n245809;
   wire n245810;
   wire n245811;
   wire n245812;
   wire n245813;
   wire n245814;
   wire n245815;
   wire n245816;
   wire n245817;
   wire n245818;
   wire n245819;
   wire n245820;
   wire n245821;
   wire n245822;
   wire n245823;
   wire n245824;
   wire n245825;
   wire n245826;
   wire n245827;
   wire n245828;
   wire n245829;
   wire n245830;
   wire n245831;
   wire n245832;
   wire n245833;
   wire n245834;
   wire n245835;
   wire n245836;
   wire n245837;
   wire n245838;
   wire n245839;
   wire n245840;
   wire n245841;
   wire n245842;
   wire n245843;
   wire n245844;
   wire n245845;
   wire n245846;
   wire n245847;
   wire n245848;
   wire n245849;
   wire n245850;
   wire n245851;
   wire n245852;
   wire n245853;
   wire n245854;
   wire n245855;
   wire n245856;
   wire n245857;
   wire n245858;
   wire n245859;
   wire n245860;
   wire n245861;
   wire n245862;
   wire n245863;
   wire n245864;
   wire n245865;
   wire n245866;
   wire n245867;
   wire n245868;
   wire n245869;
   wire n245870;
   wire n245871;
   wire n245872;
   wire n245873;
   wire n245874;
   wire n245875;
   wire n245876;
   wire n245877;
   wire n245878;
   wire n245879;
   wire n245880;
   wire n245881;
   wire n245882;
   wire n245883;
   wire n245884;
   wire n245885;
   wire n245886;
   wire n245887;
   wire n245888;
   wire n245889;
   wire n245890;
   wire n245891;
   wire n245892;
   wire n245893;
   wire n245894;
   wire n245895;
   wire n245896;
   wire n245897;
   wire n245898;
   wire n245899;
   wire n245900;
   wire n245901;
   wire n245902;
   wire n245903;
   wire n245904;
   wire n245905;
   wire n245906;
   wire n245908;
   wire n245909;
   wire n245911;
   wire n245912;
   wire n245914;
   wire n245915;
   wire n245917;
   wire n245918;
   wire n245920;
   wire n245921;
   wire n245922;
   wire n245923;
   wire n245924;
   wire n245925;
   wire n245926;
   wire n245927;
   wire n245928;
   wire n245929;
   wire n245930;
   wire n245931;
   wire n245932;
   wire n245933;
   wire n245934;
   wire n245935;
   wire n245936;
   wire n245937;
   wire n245938;
   wire n245939;
   wire n245940;
   wire n245941;
   wire n245942;
   wire n245944;
   wire n245945;
   wire n245946;
   wire n245947;
   wire n245948;
   wire n245949;
   wire n245950;
   wire n245951;
   wire n245952;
   wire n245953;
   wire n245954;
   wire n245955;
   wire n245956;
   wire n245957;
   wire n245958;
   wire n245959;
   wire n245960;
   wire n245961;
   wire n245962;
   wire n245963;
   wire n245964;
   wire n245965;
   wire n245966;
   wire n245967;
   wire n245968;
   wire n245970;
   wire n245971;
   wire n245972;
   wire n245973;
   wire n245974;
   wire n245975;
   wire n245976;
   wire n245977;
   wire n245978;
   wire n245979;
   wire n245980;
   wire n245981;
   wire n245982;
   wire n245983;
   wire n245984;
   wire n245985;
   wire n245986;
   wire n245987;
   wire n245988;
   wire n245989;
   wire n245990;
   wire n245991;
   wire n245992;
   wire n245993;
   wire n245994;
   wire n245995;
   wire n245996;
   wire n245997;
   wire n245998;
   wire n245999;
   wire n246000;
   wire n246001;
   wire n246002;
   wire n246003;
   wire n246004;
   wire n246005;
   wire n246006;
   wire n246007;
   wire n246008;
   wire n246009;
   wire n246010;
   wire n246011;
   wire n246012;
   wire n246013;
   wire n246014;
   wire n246015;
   wire n246016;
   wire n246017;
   wire n246018;
   wire n246019;
   wire n246020;
   wire n246021;
   wire n246022;
   wire n246023;
   wire n246024;
   wire n246025;
   wire n246026;
   wire n246027;
   wire n246028;
   wire n246029;
   wire n246030;
   wire n246031;
   wire n246032;
   wire n246033;
   wire n246034;
   wire n246035;
   wire n246036;
   wire n246037;
   wire n246038;
   wire n246039;
   wire n246040;
   wire n246041;
   wire n246042;
   wire n246043;
   wire n246044;
   wire n246045;
   wire n246046;
   wire n246047;
   wire n246048;
   wire n246049;
   wire n246050;
   wire n246051;
   wire n246052;
   wire n246053;
   wire n246054;
   wire n246055;
   wire n246056;
   wire n246057;
   wire n246058;
   wire n246059;
   wire n246060;
   wire n246061;
   wire n246062;
   wire n246063;
   wire n246064;
   wire n246065;
   wire n246066;
   wire n246067;
   wire n246068;
   wire n246069;
   wire n246070;
   wire n246071;
   wire n246072;
   wire n246073;
   wire n246074;
   wire n246075;
   wire n246076;
   wire n246077;
   wire n246078;
   wire n246079;
   wire n246080;
   wire n246081;
   wire n246082;
   wire n246083;
   wire n246084;
   wire n246085;
   wire n246086;
   wire n246087;
   wire n246088;
   wire n246089;
   wire n246090;
   wire n246091;
   wire n246092;
   wire n246093;
   wire n246094;
   wire n246095;
   wire n246096;
   wire n246097;
   wire n246098;
   wire n246099;
   wire n246100;
   wire n246101;
   wire n246102;
   wire n246103;
   wire n246104;
   wire n246105;
   wire n246106;
   wire n246107;
   wire n246108;
   wire n246109;
   wire n246110;
   wire n246111;
   wire n246112;
   wire n246113;
   wire n246114;
   wire n246115;
   wire n246116;
   wire n246117;
   wire n246118;
   wire n246119;
   wire n246120;
   wire n246121;
   wire n246122;
   wire n246123;
   wire n246124;
   wire n246125;
   wire n246126;
   wire n246127;
   wire n246128;
   wire n246129;
   wire n246130;
   wire n246131;
   wire n246132;
   wire n246133;
   wire n246134;
   wire n246135;
   wire n246136;
   wire n246137;
   wire n246138;
   wire n246139;
   wire n246140;
   wire n246141;
   wire n246142;
   wire n246143;
   wire n246144;
   wire n246145;
   wire n246146;
   wire n246147;
   wire n246148;
   wire n246149;
   wire n246150;
   wire n246151;
   wire n246152;
   wire n246153;
   wire n246154;
   wire n246155;
   wire n246156;
   wire n246157;
   wire n246158;
   wire n246159;
   wire n246160;
   wire n246161;
   wire n246162;
   wire n246163;
   wire n246164;
   wire n246165;
   wire n246166;
   wire n246167;
   wire n246168;
   wire n246169;
   wire n246170;
   wire n246171;
   wire n246172;
   wire n246173;
   wire n246174;
   wire n246175;
   wire n246176;
   wire n246177;
   wire n246178;
   wire n246179;
   wire n246180;
   wire n246181;
   wire n246182;
   wire n246183;
   wire n246184;
   wire n246185;
   wire n246186;
   wire n246187;
   wire n246188;
   wire n246189;
   wire n246190;
   wire n246191;
   wire n246192;
   wire n246193;
   wire n246194;
   wire n246195;
   wire n246196;
   wire n246197;
   wire n246198;
   wire n246200;
   wire n246201;
   wire n246202;
   wire n246203;
   wire n246204;
   wire n246205;
   wire n246206;
   wire n246207;
   wire n246208;
   wire n246209;
   wire n246210;
   wire n246211;
   wire n246212;
   wire n246213;
   wire n246214;
   wire n246215;
   wire n246216;
   wire n246217;
   wire n246218;
   wire n246219;
   wire n246220;
   wire n246221;
   wire n246222;
   wire n246223;
   wire n246224;
   wire n246225;
   wire n246226;
   wire n246227;
   wire n246228;
   wire n246229;
   wire n246230;
   wire n246231;
   wire n246232;
   wire n246233;
   wire n246234;
   wire n246235;
   wire n246236;
   wire n246237;
   wire n246238;
   wire n246239;
   wire n246240;
   wire n246241;
   wire n246242;
   wire n246243;
   wire n246244;
   wire n246245;
   wire n246246;
   wire n246247;
   wire n246248;
   wire n246249;
   wire n246250;
   wire n246251;
   wire n246252;
   wire n246253;
   wire n246254;
   wire n246255;
   wire n246256;
   wire n246257;
   wire n246258;
   wire n246259;
   wire n246260;
   wire n246261;
   wire n246262;
   wire n246263;
   wire n246264;
   wire n246265;
   wire n246266;
   wire n246267;
   wire n246268;
   wire n246269;
   wire n246270;
   wire n246271;
   wire n246272;
   wire n246273;
   wire n246274;
   wire n246275;
   wire n246276;
   wire n246277;
   wire n246278;
   wire n246279;
   wire n246280;
   wire n246281;
   wire n246282;
   wire n246283;
   wire n246284;
   wire n246285;
   wire n246286;
   wire n246287;
   wire n246288;
   wire n246289;
   wire n246290;
   wire n246291;
   wire n246292;
   wire n246293;
   wire n246294;
   wire n246295;
   wire n246296;
   wire n246297;
   wire n246298;
   wire n246299;
   wire n246300;
   wire n246301;
   wire n246302;
   wire n246303;
   wire n246304;
   wire n246305;
   wire n246306;
   wire n246307;
   wire n246308;
   wire n246309;
   wire n246310;
   wire n246311;
   wire n246312;
   wire n246313;
   wire n246314;
   wire n246315;
   wire n246316;
   wire n246317;
   wire n246318;
   wire n246319;
   wire n246320;
   wire n246321;
   wire n246322;
   wire n246323;
   wire n246324;
   wire n246325;
   wire n246326;
   wire n246327;
   wire n246328;
   wire n246329;
   wire n246330;
   wire n246331;
   wire n246332;
   wire n246333;
   wire n246334;
   wire n246335;
   wire n246336;
   wire n246337;
   wire n246338;
   wire n246339;
   wire n246340;
   wire n246341;
   wire n246342;
   wire n246343;
   wire n246344;
   wire n246345;
   wire n246346;
   wire n246347;
   wire n246348;
   wire n246349;
   wire n246350;
   wire n246351;
   wire n246352;
   wire n246353;
   wire n246354;
   wire n246355;
   wire n246356;
   wire n246357;
   wire n246358;
   wire n246359;
   wire n246360;
   wire n246361;
   wire n246362;
   wire n246363;
   wire n246364;
   wire n246365;
   wire n246366;
   wire n246367;
   wire n246368;
   wire n246369;
   wire n246370;
   wire n246371;
   wire n246372;
   wire n246373;
   wire n246374;
   wire n246375;
   wire n246376;
   wire n246377;
   wire n246378;
   wire n246379;
   wire n246380;
   wire n246381;
   wire n246382;
   wire n246383;
   wire n246384;
   wire n246385;
   wire n246386;
   wire n246387;
   wire n246388;
   wire n246389;
   wire n246390;
   wire n246391;
   wire n246392;
   wire n246393;
   wire n246394;
   wire n246395;
   wire n246396;
   wire n246397;
   wire n246398;
   wire n246399;
   wire n246400;
   wire n246401;
   wire n246402;
   wire n246403;
   wire n246404;
   wire n246405;
   wire n246406;
   wire n246407;
   wire n246408;
   wire n246409;
   wire n246410;
   wire n246411;
   wire n246412;
   wire n246413;
   wire n246414;
   wire n246415;
   wire n246416;
   wire n246417;
   wire n246418;
   wire n246419;
   wire n246420;
   wire n246421;
   wire n246422;
   wire n246423;
   wire n246424;
   wire n246425;
   wire n246426;
   wire n246427;
   wire n246428;
   wire n246429;
   wire n246430;
   wire n246431;
   wire n246432;
   wire n246433;
   wire n246434;
   wire n246435;
   wire n246436;
   wire n246437;
   wire n246438;
   wire n246439;
   wire n246440;
   wire n246441;
   wire n246442;
   wire n246443;
   wire n246444;
   wire n246445;
   wire n246446;
   wire n246447;
   wire n246448;
   wire n246449;
   wire n246450;
   wire n246451;
   wire n246452;
   wire n246453;
   wire n246454;
   wire n246455;
   wire n246456;
   wire n246457;
   wire n246458;
   wire n246459;
   wire n246460;
   wire n246461;
   wire n246462;
   wire n246463;
   wire n246464;
   wire n246465;
   wire n246466;
   wire n246467;
   wire n246468;
   wire n246469;
   wire n246470;
   wire n246471;
   wire n246472;
   wire n246473;
   wire n246474;
   wire n246475;
   wire n246476;
   wire n246477;
   wire n246478;
   wire n246479;
   wire n246480;
   wire n246481;
   wire n246482;
   wire n246483;
   wire n246484;
   wire n246485;
   wire n246486;
   wire n246487;
   wire n246488;
   wire n246489;
   wire n246490;
   wire n246491;
   wire n246492;
   wire n246493;
   wire n246494;
   wire n246495;
   wire n246496;
   wire n246497;
   wire n246498;
   wire n246499;
   wire n246500;
   wire n246501;
   wire n246502;
   wire n246503;
   wire n246504;
   wire n246505;
   wire n246506;
   wire n246507;
   wire n246508;
   wire n246509;
   wire n246510;
   wire n246511;
   wire n246512;
   wire n246513;
   wire n246514;
   wire n246515;
   wire n246516;
   wire n246517;
   wire n246518;
   wire n246519;
   wire n246520;
   wire n246521;
   wire n246522;
   wire n246523;
   wire n246524;
   wire n246525;
   wire n246526;
   wire n246527;
   wire n246528;
   wire n246529;
   wire n246530;
   wire n246531;
   wire n246532;
   wire n246533;
   wire n246534;
   wire n246535;
   wire n246536;
   wire n246537;
   wire n246538;
   wire n246539;
   wire n246540;
   wire n246541;
   wire n246542;
   wire n246543;
   wire n246544;
   wire n246545;
   wire n246546;
   wire n246547;
   wire n246548;
   wire n246549;
   wire n246550;
   wire n246551;
   wire n246552;
   wire n246553;
   wire n246554;
   wire n246555;
   wire n246556;
   wire n246557;
   wire n246558;
   wire n246559;
   wire n246560;
   wire n246561;
   wire n246562;
   wire n246563;
   wire n246564;
   wire n246565;
   wire n246566;
   wire n246567;
   wire n246568;
   wire n246569;
   wire n246570;
   wire n246571;
   wire n246572;
   wire n246573;
   wire n246574;
   wire n246575;
   wire n246576;
   wire n246577;
   wire n246578;
   wire n246579;
   wire n246580;
   wire n246581;
   wire n246582;
   wire n246583;
   wire n246584;
   wire n246585;
   wire n246586;
   wire n246587;
   wire n246588;
   wire n246589;
   wire n246590;
   wire n246591;
   wire n246592;
   wire n246593;
   wire n246594;
   wire n246595;
   wire n246596;
   wire n246597;
   wire n246598;
   wire n246599;
   wire n246600;
   wire n246601;
   wire n246602;
   wire n246603;
   wire n246604;
   wire n246606;
   wire n246607;
   wire n246608;
   wire n246609;
   wire n246610;
   wire n246611;
   wire n246612;
   wire n246613;
   wire n246614;
   wire n246615;
   wire n246617;
   wire n246618;
   wire n246619;
   wire n246620;
   wire n246621;
   wire n246623;
   wire n246624;
   wire n246625;
   wire n246627;
   wire n246628;
   wire n246629;
   wire n246631;
   wire n246632;
   wire n246633;
   wire n246635;
   wire n246636;
   wire n246637;
   wire n246638;
   wire n246639;
   wire n246640;
   wire n246641;
   wire n246642;
   wire n246643;
   wire n246644;
   wire n246645;
   wire n246646;
   wire n246647;
   wire n246648;
   wire n246649;
   wire n246650;
   wire n246651;
   wire n246652;
   wire n246653;
   wire n246654;
   wire n246655;
   wire n246656;
   wire n246657;
   wire n246658;
   wire n246659;
   wire n246660;
   wire n246661;
   wire n246662;
   wire n246663;
   wire n246664;
   wire n246665;
   wire n246666;
   wire n246667;
   wire n246668;
   wire n246669;
   wire n246670;
   wire n246671;
   wire n246672;
   wire n246673;
   wire n246674;
   wire n246675;
   wire n246676;
   wire n246677;
   wire n246678;
   wire n246679;
   wire n246680;
   wire n246681;
   wire n246682;
   wire n246683;
   wire n246684;
   wire n246685;
   wire n246686;
   wire n246687;
   wire n246688;
   wire n246689;
   wire n246690;
   wire n246691;
   wire n246692;
   wire n246693;
   wire n246694;
   wire n246695;
   wire n246696;
   wire n246697;
   wire n246698;
   wire n246699;
   wire n246700;
   wire n246701;
   wire n246702;
   wire n246703;
   wire n246704;
   wire n246705;
   wire n246706;
   wire n246707;
   wire n246708;
   wire n246709;
   wire n246710;
   wire n246711;
   wire n246712;
   wire n246713;
   wire n246714;
   wire n246715;
   wire n246716;
   wire n246717;
   wire n246718;
   wire n246719;
   wire n246720;
   wire n246721;
   wire n246722;
   wire n246723;
   wire n246724;
   wire n246725;
   wire n246726;
   wire n246727;
   wire n246728;
   wire n246729;
   wire n246730;
   wire n246731;
   wire n246732;
   wire n246733;
   wire n246734;
   wire n246735;
   wire n246736;
   wire n246737;
   wire n246738;
   wire n246739;
   wire n246740;
   wire n246741;
   wire n246742;
   wire n246743;
   wire n246745;
   wire n246746;
   wire n246747;
   wire n246748;
   wire n246749;
   wire n246750;
   wire n246751;
   wire n246752;
   wire n246753;
   wire n246754;
   wire n246755;
   wire n246756;
   wire n246757;
   wire n246758;
   wire n246759;
   wire n246760;
   wire n246761;
   wire n246762;
   wire n246763;
   wire n246764;
   wire n246765;
   wire n246766;
   wire n246767;
   wire n246768;
   wire n246769;
   wire n246770;
   wire n246771;
   wire n246772;
   wire n246773;
   wire n246774;
   wire n246775;
   wire n246776;
   wire n246777;
   wire n246778;
   wire n246779;
   wire n246780;
   wire n246781;
   wire n246782;
   wire n246783;
   wire n246784;
   wire n246785;
   wire n246786;
   wire n246787;
   wire n246788;
   wire n246789;
   wire n246790;
   wire n246791;
   wire n246792;
   wire n246793;
   wire n246794;
   wire n246795;
   wire n246796;
   wire n246797;
   wire n246798;
   wire n246799;
   wire n246800;
   wire n246801;
   wire n246802;
   wire n246803;
   wire n246804;
   wire n246805;
   wire n246806;
   wire n246807;
   wire n246808;
   wire n246809;
   wire n246810;
   wire n246811;
   wire n246812;
   wire n246813;
   wire n246814;
   wire n246815;
   wire n246816;
   wire n246817;
   wire n246818;
   wire n246819;
   wire n246820;
   wire n246821;
   wire n246822;
   wire n246823;
   wire n246824;
   wire n246825;
   wire n246826;
   wire n246827;
   wire n246828;
   wire n246829;
   wire n246830;
   wire n246831;
   wire n246832;
   wire n246833;
   wire n246834;
   wire n246835;
   wire n246836;
   wire n246837;
   wire n246838;
   wire n246839;
   wire n246840;
   wire n246841;
   wire n246842;
   wire n246843;
   wire n246844;
   wire n246845;
   wire n246846;
   wire n246847;
   wire n246848;
   wire n246849;
   wire n246850;
   wire n246851;
   wire n246852;
   wire n246853;
   wire n246854;
   wire n246855;
   wire n246856;
   wire n246857;
   wire n246858;
   wire n246859;
   wire n246860;
   wire n246861;
   wire n246862;
   wire n246863;
   wire n246864;
   wire n246865;
   wire n246866;
   wire n246867;
   wire n246868;
   wire n246869;
   wire n246870;
   wire n246871;
   wire n246872;
   wire n246873;
   wire n246874;
   wire n246875;
   wire n246876;
   wire n246877;
   wire n246878;
   wire n246879;
   wire n246880;
   wire n246881;
   wire n246882;
   wire n246883;
   wire n246884;
   wire n246885;
   wire n246886;
   wire n246887;
   wire n246888;
   wire n246889;
   wire n246890;
   wire n246891;
   wire n246892;
   wire n246893;
   wire n246894;
   wire n246895;
   wire n246896;
   wire n246897;
   wire n246898;
   wire n246899;
   wire n246900;
   wire n246901;
   wire n246902;
   wire n246903;
   wire n246904;
   wire n246905;
   wire n246906;
   wire n246907;
   wire n246908;
   wire n246909;
   wire n246910;
   wire n246911;
   wire n246912;
   wire n246913;
   wire n246914;
   wire n246915;
   wire n246916;
   wire n246917;
   wire n246918;
   wire n246919;
   wire n246920;
   wire n246921;
   wire n246922;
   wire n246923;
   wire n246924;
   wire n246925;
   wire n246926;
   wire n246927;
   wire n246928;
   wire n246929;
   wire n246930;
   wire n246931;
   wire n246932;
   wire n246933;
   wire n246934;
   wire n246935;
   wire n246936;
   wire n246937;
   wire n246938;
   wire n246939;
   wire n246940;
   wire n246941;
   wire n246942;
   wire n246943;
   wire n246944;
   wire n246945;
   wire n246946;
   wire n246947;
   wire n246948;
   wire n246949;
   wire n246950;
   wire n246951;
   wire n246952;
   wire n246953;
   wire n246954;
   wire n246955;
   wire n246956;
   wire n246957;
   wire n246958;
   wire n246959;
   wire n246960;
   wire n246961;
   wire n246962;
   wire n246963;
   wire n246964;
   wire n246965;
   wire n246966;
   wire n246967;
   wire n246968;
   wire n246969;
   wire n246970;
   wire n246971;
   wire n246972;
   wire n246973;
   wire n246974;
   wire n246975;
   wire n246976;
   wire n246977;
   wire n246978;
   wire n246979;
   wire n246980;
   wire n246981;
   wire n246982;
   wire n246983;
   wire n246984;
   wire n246985;
   wire n246986;
   wire n246987;
   wire n246988;
   wire n246989;
   wire n246990;
   wire n246991;
   wire n246992;
   wire n246993;
   wire n246994;
   wire n246995;
   wire n246996;
   wire n246997;
   wire n246998;
   wire n246999;
   wire n247000;
   wire n247001;
   wire n247002;
   wire n247003;
   wire n247004;
   wire n247005;
   wire n247006;
   wire n247007;
   wire n247008;
   wire n247009;
   wire n247010;
   wire n247011;
   wire n247012;
   wire n247013;
   wire n247014;
   wire n247015;
   wire n247016;
   wire n247017;
   wire n247018;
   wire n247019;
   wire n247020;
   wire n247021;
   wire n247022;
   wire n247023;
   wire n247024;
   wire n247025;
   wire n247026;
   wire n247027;
   wire n247028;
   wire n247029;
   wire n247030;
   wire n247031;
   wire n247032;
   wire n247033;
   wire n247034;
   wire n247035;
   wire n247036;
   wire n247037;
   wire n247038;
   wire n247039;
   wire n247040;
   wire n247041;
   wire n247042;
   wire n247043;
   wire n247044;
   wire n247045;
   wire n247046;
   wire n247047;
   wire n247048;
   wire n247049;
   wire n247050;
   wire n247051;
   wire n247052;
   wire n247053;
   wire n247054;
   wire n247055;
   wire n247056;
   wire n247057;
   wire n247059;
   wire n247060;
   wire n247061;
   wire n247062;
   wire n247063;
   wire n247064;
   wire n247065;
   wire n247066;
   wire n247067;
   wire n247069;
   wire n247070;
   wire n247071;
   wire n247072;
   wire n247073;
   wire n247074;
   wire n247076;
   wire n247077;
   wire n247078;
   wire n247079;
   wire n247080;
   wire n247081;
   wire n247082;
   wire n247083;
   wire n247084;
   wire n247085;
   wire n247086;
   wire n247087;
   wire n247088;
   wire n247089;
   wire n247090;
   wire n247091;
   wire n247092;
   wire n247094;
   wire n247095;
   wire n247096;
   wire n247097;
   wire n247098;
   wire n247099;
   wire n247101;
   wire n247102;
   wire n247103;
   wire n247104;
   wire n247105;
   wire n247107;
   wire n247109;
   wire n247110;
   wire n247111;
   wire n247112;
   wire n247113;
   wire n247114;
   wire n247115;
   wire n247116;
   wire n247117;
   wire n247118;
   wire n247119;
   wire n247120;
   wire n247121;
   wire n247122;
   wire n247123;
   wire n247124;
   wire n247125;
   wire n247126;
   wire n247127;
   wire n247128;
   wire n247129;
   wire n247130;
   wire n247131;
   wire n247132;
   wire n247133;
   wire n247134;
   wire n247135;
   wire n247136;
   wire n247137;
   wire n247138;
   wire n247139;
   wire n247140;
   wire n247141;
   wire n247142;
   wire n247143;
   wire n247144;
   wire n247145;
   wire n247146;
   wire n247147;
   wire n247148;
   wire n247149;
   wire n247150;
   wire n247151;
   wire n247152;
   wire n247153;
   wire n247154;
   wire n247156;
   wire n247157;
   wire n247158;
   wire n247159;
   wire n247160;
   wire n247161;
   wire n247162;
   wire n247163;
   wire n247164;
   wire n247165;
   wire n247166;
   wire n247167;
   wire n247168;
   wire n247169;
   wire n247170;
   wire n247171;
   wire n247172;
   wire n247173;
   wire n247174;
   wire n247175;
   wire n247176;
   wire n247177;
   wire n247178;
   wire n247179;
   wire n247180;
   wire n247181;
   wire n247182;
   wire n247184;
   wire n247185;
   wire n247186;
   wire n247187;
   wire n247188;
   wire n247189;
   wire n247190;
   wire n247191;
   wire n247192;
   wire n247193;
   wire n247194;
   wire n247195;
   wire n247196;
   wire n247197;
   wire n247198;
   wire n247199;
   wire n247200;
   wire n247201;
   wire n247202;
   wire n247204;
   wire n247205;
   wire n247206;
   wire n247207;
   wire n247208;
   wire n247209;
   wire n247210;
   wire n247211;
   wire n247212;
   wire n247213;
   wire n247214;
   wire n247215;
   wire n247216;
   wire n247217;
   wire n247218;
   wire n247219;
   wire n247220;
   wire n247221;
   wire n247222;
   wire n247223;
   wire n247224;
   wire n247225;
   wire n247226;
   wire n247227;
   wire n247228;
   wire n247229;
   wire n247230;
   wire n247231;
   wire n247232;
   wire n247233;
   wire n247234;
   wire n247235;
   wire n247236;
   wire n247237;
   wire n247238;
   wire n247239;
   wire n247241;
   wire n247242;
   wire n247243;
   wire n247244;
   wire n247245;
   wire n247246;
   wire n247247;
   wire n247248;
   wire n247249;
   wire n247250;
   wire n247251;
   wire n247252;
   wire n247253;
   wire n247254;
   wire n247255;
   wire n247256;
   wire n247257;
   wire n247258;
   wire n247259;
   wire n247260;
   wire n247261;
   wire n247262;
   wire n247263;
   wire n247264;
   wire n247265;
   wire n247266;
   wire n247267;
   wire n247268;
   wire n247269;
   wire n247270;
   wire n247271;
   wire n247273;
   wire n247274;
   wire n247275;
   wire n247276;
   wire n247277;
   wire n247278;
   wire n247279;
   wire n247280;
   wire n247281;
   wire n247282;
   wire n247283;
   wire n247284;
   wire n247285;
   wire n247286;
   wire n247288;
   wire n247289;
   wire n247290;
   wire n247291;
   wire n247292;
   wire n247293;
   wire n247294;
   wire n247295;
   wire n247296;
   wire n247297;
   wire n247298;
   wire n247299;
   wire n247300;
   wire n247301;
   wire n247302;
   wire n247304;
   wire n247305;
   wire n247306;
   wire n247307;
   wire n247308;
   wire n247309;
   wire n247310;
   wire n247311;
   wire n247312;
   wire n247313;
   wire n247314;
   wire n247315;
   wire n247317;
   wire n247318;
   wire n247319;
   wire n247320;
   wire n247321;
   wire n247322;
   wire n247323;
   wire n247324;
   wire n247325;
   wire n247326;
   wire n247327;
   wire n247328;
   wire n247329;
   wire n247330;
   wire n247331;
   wire n247332;
   wire n247333;
   wire n247334;
   wire n247335;
   wire n247336;
   wire n247337;
   wire n247338;
   wire n247339;
   wire n247340;
   wire n247341;
   wire n247342;
   wire n247343;
   wire n247344;
   wire n247345;
   wire n247346;
   wire n247347;
   wire n247348;
   wire n247349;
   wire n247350;
   wire n247351;
   wire n247352;
   wire n247354;
   wire n247355;
   wire n247356;
   wire n247357;
   wire n247358;
   wire n247359;
   wire n247360;
   wire n247361;
   wire n247362;
   wire n247363;
   wire n247364;
   wire n247365;
   wire n247366;
   wire n247367;
   wire n247368;
   wire n247369;
   wire n247370;
   wire n247371;
   wire n247372;
   wire n247373;
   wire n247374;
   wire n247375;
   wire n247376;
   wire n247377;
   wire n247378;
   wire n247379;
   wire n247380;
   wire n247381;
   wire n247382;
   wire n247383;
   wire n247384;
   wire n247385;
   wire n247386;
   wire n247387;
   wire n247388;
   wire n247389;
   wire n247390;
   wire n247391;
   wire n247392;
   wire n247393;
   wire n247395;
   wire n247396;
   wire n247397;
   wire n247398;
   wire n247400;
   wire n247401;
   wire n247402;
   wire n247403;
   wire n247404;
   wire n247405;
   wire n247406;
   wire n247407;
   wire n247409;
   wire n247410;
   wire n247411;
   wire n247412;
   wire n247413;
   wire n247414;
   wire n247415;
   wire n247416;
   wire n247418;
   wire n247419;
   wire n247420;
   wire n247421;
   wire n247422;
   wire n247423;
   wire n247424;
   wire n247425;
   wire n247426;
   wire n247427;
   wire n247428;
   wire n247429;
   wire n247431;
   wire n247432;
   wire n247433;
   wire n247434;
   wire n247435;
   wire n247436;
   wire n247437;
   wire n247438;
   wire n247439;
   wire n247440;
   wire n247441;
   wire n247442;
   wire n247443;
   wire n247444;
   wire n247445;
   wire n247446;
   wire n247447;
   wire n247448;
   wire n247449;
   wire n247450;
   wire n247451;
   wire n247453;
   wire n247454;
   wire n247455;
   wire n247456;
   wire n247457;
   wire n247458;
   wire n247459;
   wire n247460;
   wire n247461;
   wire n247462;
   wire n247463;
   wire n247464;
   wire n247465;
   wire n247466;
   wire n247467;
   wire n247468;
   wire n247469;
   wire n247470;
   wire n247471;
   wire n247472;
   wire n247473;
   wire n247474;
   wire n247475;
   wire n247476;
   wire n247477;
   wire n247478;
   wire n247479;
   wire n247480;
   wire n247481;
   wire n247482;
   wire n247483;
   wire n247484;
   wire n247485;
   wire n247486;
   wire n247487;
   wire n247489;
   wire n247490;
   wire n247491;
   wire n247492;
   wire n247493;
   wire n247494;
   wire n247495;
   wire n247496;
   wire n247497;
   wire n247498;
   wire n247499;
   wire n247500;
   wire n247501;
   wire n247502;
   wire n247503;
   wire n247504;
   wire n247505;
   wire n247506;
   wire n247507;
   wire n247508;
   wire n247509;
   wire n247511;
   wire n247512;
   wire n247513;
   wire n247514;
   wire n247515;
   wire n247516;
   wire n247517;
   wire n247518;
   wire n247519;
   wire n247520;
   wire n247521;
   wire n247522;
   wire n247523;
   wire n247524;
   wire n247525;
   wire n247526;
   wire n247527;
   wire n247528;
   wire n247529;
   wire n247530;
   wire n247531;
   wire n247533;
   wire n247534;
   wire n247535;
   wire n247536;
   wire n247537;
   wire n247538;
   wire n247539;
   wire n247540;
   wire n247541;
   wire n247542;
   wire n247543;
   wire n247544;
   wire n247545;
   wire n247546;
   wire n247547;
   wire n247548;
   wire n247549;
   wire n247550;
   wire n247551;
   wire n247552;
   wire n247553;
   wire n247554;
   wire n247555;
   wire n247556;
   wire n247557;
   wire n247558;
   wire n247559;
   wire n247560;
   wire n247561;
   wire n247562;
   wire n247563;
   wire n247564;
   wire n247565;
   wire n247566;
   wire n247567;
   wire n247568;
   wire n247569;
   wire n247570;
   wire n247571;
   wire n247572;
   wire n247573;
   wire n247574;
   wire n247575;
   wire n247576;
   wire n247577;
   wire n247578;
   wire n247579;
   wire n247580;
   wire n247581;
   wire n247582;
   wire n247583;
   wire n247584;
   wire n247585;
   wire n247586;
   wire n247587;
   wire n247588;
   wire n247589;
   wire n247590;
   wire n247591;
   wire n247592;
   wire n247593;
   wire n247594;
   wire n247595;
   wire n247596;
   wire n247597;
   wire n247598;
   wire n247599;
   wire n247600;
   wire n247601;
   wire n247602;
   wire n247603;
   wire n247604;
   wire n247611;
   wire n247612;
   wire n247613;
   wire n247614;
   wire n247621;
   wire n247622;
   wire n247623;
   wire n247624;
   wire n247632;
   wire n247633;
   wire n247634;
   wire n247635;
   wire n247642;
   wire n247643;
   wire n247644;
   wire n247645;
   wire n247646;
   wire n247647;
   wire n247648;
   wire n247649;
   wire n247656;
   wire n247657;
   wire n247658;
   wire n247659;
   wire n247667;
   wire n247668;
   wire n247669;
   wire n247670;
   wire n247678;
   wire n247679;
   wire n247680;
   wire n247681;
   wire n247688;
   wire n247689;
   wire n247690;
   wire n247691;
   wire n247692;
   wire n247693;
   wire n247694;
   wire n247695;
   wire n247696;
   wire n247697;
   wire n247698;
   wire n247699;
   wire n247700;
   wire n247701;
   wire n247702;
   wire n247703;
   wire n247704;
   wire n247705;
   wire n247706;
   wire n247707;
   wire n247708;
   wire n247709;
   wire n247710;
   wire n247711;
   wire n247712;
   wire n247713;
   wire n247714;
   wire n247715;
   wire n247716;
   wire n247717;
   wire n247718;
   wire n247719;
   wire n247720;
   wire n247721;
   wire n247722;
   wire n247723;
   wire n247724;
   wire n247725;
   wire n247726;
   wire n247727;
   wire n247728;
   wire n247729;
   wire n247730;
   wire n247731;
   wire n247732;
   wire n247733;
   wire n247734;
   wire n247735;
   wire n247736;
   wire n247737;
   wire n247738;
   wire n247739;
   wire n247740;
   wire n247741;
   wire n247742;
   wire n247743;
   wire n247744;
   wire n247745;
   wire n247746;
   wire n247747;
   wire n247748;
   wire n247749;
   wire n247750;
   wire n247751;
   wire n247752;
   wire n247753;
   wire n247754;
   wire n247755;
   wire n247756;
   wire n247757;
   wire n247758;
   wire n247759;
   wire n247760;
   wire n247761;
   wire n247762;
   wire n247763;
   wire n247764;
   wire n247765;
   wire n247766;
   wire n247767;
   wire n247768;
   wire n247769;
   wire n247770;
   wire n247771;
   wire n247772;
   wire n247773;
   wire n247774;
   wire n247775;
   wire n247776;
   wire n247777;
   wire n247778;
   wire n247779;
   wire n247780;
   wire n247781;
   wire n247782;
   wire n247783;
   wire n247784;
   wire n247785;
   wire n247786;
   wire n247787;
   wire n247788;
   wire n247789;
   wire n247790;
   wire n247791;
   wire n247792;
   wire n247793;
   wire n247794;
   wire n247795;
   wire n247796;
   wire n247797;
   wire n247798;
   wire n247799;
   wire n247800;
   wire n247801;
   wire n247802;
   wire n247803;
   wire n247804;
   wire n247805;
   wire n247806;
   wire n247807;
   wire n247808;
   wire n247809;
   wire n247810;
   wire n247811;
   wire n247812;
   wire n247813;
   wire n247814;
   wire n247815;
   wire n247816;
   wire n247817;
   wire n247818;
   wire n247819;
   wire n247820;
   wire n247821;
   wire n247822;
   wire n247823;
   wire n247824;
   wire n247825;
   wire n247826;
   wire n247827;
   wire n247828;
   wire n247829;
   wire n247830;
   wire n247831;
   wire n247832;
   wire n247833;
   wire n247834;
   wire n247835;
   wire n247836;
   wire n247837;
   wire n247838;
   wire n247839;
   wire n247840;
   wire n247841;
   wire n247842;
   wire n247843;
   wire n247844;
   wire n247845;
   wire n247846;
   wire n247847;
   wire n247848;
   wire n247849;
   wire n247850;
   wire n247851;
   wire n247852;
   wire n247853;
   wire n247854;
   wire n247855;
   wire n247856;
   wire n247857;
   wire n247858;
   wire n247859;
   wire n247860;
   wire n247861;
   wire n247862;
   wire n247863;
   wire n247864;
   wire n247865;
   wire n247866;
   wire n247867;
   wire n247868;
   wire n247869;
   wire n247870;
   wire n247871;
   wire n247872;
   wire n247873;
   wire n247874;
   wire n247875;
   wire n247876;
   wire n247877;
   wire n247878;
   wire n247879;
   wire n247880;
   wire n247881;
   wire n247882;
   wire n247883;
   wire n247884;
   wire n247885;
   wire n247886;
   wire n247887;
   wire n247888;
   wire n247889;
   wire n247890;
   wire n247891;
   wire n247892;
   wire n247893;
   wire n247894;
   wire n247895;
   wire n247896;
   wire n247897;
   wire n247898;
   wire n247899;
   wire n247900;
   wire n247901;
   wire n247902;
   wire n247903;
   wire n247904;
   wire n247905;
   wire n247906;
   wire n247907;
   wire n247908;
   wire n247909;
   wire n247910;
   wire n247911;
   wire n247912;
   wire n247913;
   wire n247914;
   wire n247915;
   wire n247916;
   wire n247917;
   wire n247918;
   wire n247919;
   wire n247920;
   wire n247921;
   wire n247922;
   wire n247923;
   wire n247924;
   wire n247925;
   wire n247926;
   wire n247927;
   wire n247928;
   wire n247929;
   wire n247930;
   wire n247931;
   wire n247932;
   wire n247933;
   wire n247934;
   wire n247935;
   wire n247936;
   wire n247937;
   wire n247938;
   wire n247939;
   wire n247940;
   wire n247941;
   wire n247942;
   wire n247943;
   wire n247944;
   wire n247945;
   wire n247946;
   wire n247947;
   wire n247948;
   wire n247949;
   wire n247950;
   wire n247951;
   wire n247952;
   wire n247953;
   wire n247954;
   wire n247955;
   wire n247956;
   wire n247957;
   wire n247958;
   wire n247959;
   wire n247960;
   wire n247961;
   wire n247962;
   wire n247963;
   wire n247964;
   wire n247965;
   wire n247966;
   wire n247967;
   wire n247968;
   wire n247969;
   wire n247970;
   wire n247971;
   wire n247972;
   wire n247973;
   wire n247974;
   wire n247975;
   wire n247976;
   wire n247977;
   wire n247978;
   wire n247979;
   wire n247980;
   wire n247981;
   wire n247982;
   wire n247983;
   wire n247984;
   wire n247985;
   wire n247986;
   wire n247987;
   wire n247988;
   wire n247989;
   wire n247990;
   wire n247991;
   wire n247992;
   wire n247993;
   wire n247994;
   wire n247995;
   wire n247996;
   wire n247997;
   wire n247998;
   wire n247999;
   wire n248000;
   wire n248001;
   wire n248002;
   wire n248003;
   wire n248004;
   wire n248005;
   wire n248006;
   wire n248007;
   wire n248008;
   wire n248009;
   wire n248010;
   wire n248011;
   wire n248012;
   wire n248013;
   wire n248014;
   wire n248015;
   wire n248016;
   wire n248017;
   wire n248018;
   wire n248019;
   wire n248020;
   wire n248021;
   wire n248022;
   wire n248023;
   wire n248024;
   wire n248025;
   wire n248026;
   wire n248027;
   wire n248028;
   wire n248029;
   wire n248030;
   wire n248031;
   wire n248032;
   wire n248033;
   wire n248034;
   wire n248035;
   wire n248036;
   wire n248037;
   wire n248038;
   wire n248039;
   wire n248040;
   wire n248041;
   wire n248042;
   wire n248043;
   wire n248044;
   wire n248045;
   wire n248046;
   wire n248047;
   wire n248048;
   wire n248049;
   wire n248050;
   wire n248051;
   wire n248052;
   wire n248053;
   wire n248054;
   wire n248055;
   wire n248056;
   wire n248057;
   wire n248058;
   wire n248059;
   wire n248060;
   wire n248061;
   wire n248062;
   wire n248063;
   wire n248064;
   wire n248065;
   wire n248066;
   wire n248067;
   wire n248068;
   wire n248069;
   wire n248070;
   wire n248071;
   wire n248072;
   wire n248073;
   wire n248074;
   wire n248075;
   wire n248076;
   wire n248077;
   wire n248078;
   wire n248079;
   wire n248080;
   wire n248081;
   wire n248082;
   wire n248083;
   wire n248084;
   wire n248085;
   wire n248086;
   wire n248087;
   wire n248088;
   wire n248089;
   wire n248090;
   wire n248091;
   wire n248092;
   wire n248093;
   wire n248094;
   wire n248095;
   wire n248096;
   wire n248097;
   wire n248098;
   wire n248099;
   wire n248100;
   wire n248101;
   wire n248102;
   wire n248103;
   wire n248104;
   wire n248105;
   wire n248106;
   wire n248107;
   wire n248108;
   wire n248109;
   wire n248110;
   wire n248111;
   wire n248112;
   wire n248113;
   wire n248114;
   wire n248115;
   wire n248116;
   wire n248117;
   wire n248118;
   wire n248119;
   wire n248120;
   wire n248121;
   wire n248122;
   wire n248123;
   wire n248124;
   wire n248125;
   wire n248126;
   wire n248127;
   wire n248128;
   wire n248129;
   wire n248130;
   wire n248131;
   wire n248132;
   wire n248133;
   wire n248134;
   wire n248135;
   wire n248136;
   wire n248137;
   wire n248138;
   wire n248139;
   wire n248140;
   wire n248141;
   wire n248142;
   wire n248143;
   wire n248144;
   wire n248145;
   wire n248146;
   wire n248147;
   wire n248148;
   wire n248149;
   wire n248150;
   wire n248151;
   wire n248152;
   wire n248153;
   wire n248154;
   wire n248155;
   wire n248156;
   wire n248157;
   wire n248158;
   wire n248159;
   wire n248160;
   wire n248161;
   wire n248162;
   wire n248163;
   wire n248164;
   wire n248165;
   wire n248166;
   wire n248167;
   wire n248168;
   wire n248169;
   wire n248170;
   wire n248171;
   wire n248172;
   wire n248173;
   wire n248174;
   wire n248175;
   wire n248176;
   wire n248177;
   wire n248178;
   wire n248179;
   wire n248180;
   wire n248181;
   wire n248182;
   wire n248183;
   wire n248184;
   wire n248185;
   wire n248186;
   wire n248187;
   wire n248188;
   wire n248189;
   wire n248190;
   wire n248191;
   wire n248192;
   wire n248193;
   wire n248194;
   wire n248195;
   wire n248196;
   wire n248197;
   wire n248198;
   wire n248199;
   wire n248200;
   wire n248201;
   wire n248202;
   wire n248203;
   wire n248204;
   wire n248205;
   wire n248206;
   wire n248207;
   wire n248208;
   wire n248209;
   wire n248210;
   wire n248211;
   wire n248212;
   wire n248213;
   wire n248214;
   wire n248215;
   wire n248216;
   wire n248217;
   wire n248218;
   wire n248219;
   wire n248220;
   wire n248221;
   wire n248222;
   wire n248223;
   wire n248224;
   wire n248225;
   wire n248226;
   wire n248227;
   wire n248228;
   wire n248229;
   wire n248230;
   wire n248231;
   wire n248232;
   wire n248233;
   wire n248234;
   wire n248235;
   wire n248236;
   wire n248237;
   wire n248238;
   wire n248239;
   wire n248240;
   wire n248241;
   wire n248242;
   wire n248243;
   wire n248244;
   wire n248245;
   wire n248246;
   wire n248247;
   wire n248248;
   wire n248249;
   wire n248250;
   wire n248251;
   wire n248252;
   wire n248253;
   wire n248254;
   wire n248255;
   wire n248256;
   wire n248257;
   wire n248258;
   wire n248259;
   wire n248260;
   wire n248261;
   wire n248262;
   wire n248263;
   wire n248264;
   wire n248265;
   wire n248266;
   wire n248267;
   wire n248268;
   wire n248269;
   wire n248270;
   wire n248271;
   wire n248272;
   wire n248273;
   wire n248274;
   wire n248275;
   wire n248276;
   wire n248277;
   wire n248278;
   wire n248279;
   wire n248280;
   wire n248281;
   wire n248282;
   wire n248283;
   wire n248284;
   wire n248285;
   wire n248286;
   wire n248287;
   wire n248288;
   wire n248289;
   wire n248290;
   wire n248291;
   wire n248292;
   wire n248293;
   wire n248294;
   wire n248295;
   wire n248296;
   wire n248297;
   wire n248298;
   wire n248299;
   wire n248300;
   wire n248301;
   wire n248302;
   wire n248303;
   wire n248304;
   wire n248305;
   wire n248306;
   wire n248307;
   wire n248308;
   wire n248309;
   wire n248310;
   wire n248311;
   wire n248312;
   wire n248313;
   wire n248314;
   wire n248315;
   wire n248316;
   wire n248317;
   wire n248318;
   wire n248319;
   wire n248320;
   wire n248321;
   wire n248322;
   wire n248323;
   wire n248324;
   wire n248325;
   wire n248326;
   wire n248327;
   wire n248328;
   wire n248329;
   wire n248330;
   wire n248331;
   wire n248332;
   wire n248333;
   wire n248334;
   wire n248335;
   wire n248336;
   wire n248337;
   wire n248338;
   wire n248339;
   wire n248340;
   wire n248341;
   wire n248342;
   wire n248343;
   wire n248344;
   wire n248345;
   wire n248346;
   wire n248347;
   wire n248348;
   wire n248349;
   wire n248350;
   wire n248351;
   wire n248352;
   wire n248353;
   wire n248354;
   wire n248355;
   wire n248356;
   wire n248357;
   wire n248358;
   wire n248359;
   wire n248360;
   wire n248361;
   wire n248362;
   wire n248363;
   wire n248364;
   wire n248365;
   wire n248366;
   wire n248367;
   wire n248368;
   wire n248369;
   wire n248370;
   wire n248371;
   wire n248372;
   wire n248373;
   wire n248374;
   wire n248375;
   wire n248376;
   wire n248377;
   wire n248378;
   wire n248379;
   wire n248380;
   wire n248381;
   wire n248382;
   wire n248383;
   wire n248384;
   wire n248385;
   wire n248386;
   wire n248387;
   wire n248388;
   wire n248389;
   wire n248390;
   wire n248391;
   wire n248392;
   wire n248393;
   wire n248394;
   wire n248395;
   wire n248396;
   wire n248397;
   wire n248398;
   wire n248399;
   wire n248400;
   wire n248401;
   wire n248402;
   wire n248403;
   wire n248404;
   wire n248405;
   wire n248406;
   wire n248407;
   wire n248408;
   wire n248409;
   wire n248410;
   wire n248411;
   wire n248412;
   wire n248413;
   wire n248414;
   wire n248415;
   wire n248416;
   wire n248417;
   wire n248418;
   wire n248419;
   wire n248420;
   wire n248421;
   wire n248422;
   wire n248423;
   wire n248424;
   wire n248425;
   wire n248426;
   wire n248427;
   wire n248428;
   wire n248429;
   wire n248430;
   wire n248431;
   wire n248432;
   wire n248433;
   wire n248434;
   wire n248435;
   wire n248436;
   wire n248437;
   wire n248438;
   wire n248439;
   wire n248440;
   wire n248441;
   wire n248442;
   wire n248443;
   wire n248444;
   wire n248445;
   wire n248446;
   wire n248447;
   wire n248448;
   wire n248449;
   wire n248450;
   wire n248451;
   wire n248452;
   wire n248453;
   wire n248454;
   wire n248455;
   wire n248456;
   wire n248457;
   wire n248458;
   wire n248459;
   wire n248460;
   wire n248461;
   wire n248462;
   wire n248463;
   wire n248464;
   wire n248465;
   wire n248466;
   wire n248467;
   wire n248468;
   wire n248469;
   wire n248470;
   wire n248471;
   wire n248472;
   wire n248473;
   wire n248474;
   wire n248475;
   wire n248476;
   wire n248477;
   wire n248478;
   wire n248479;
   wire n248480;
   wire n248481;
   wire n248482;
   wire n248483;
   wire n248484;
   wire n248485;
   wire n248486;
   wire n248487;
   wire n248488;
   wire n248489;
   wire n248490;
   wire n248491;
   wire n248492;
   wire n248493;
   wire n248494;
   wire n248495;
   wire n248496;
   wire n248497;
   wire n248498;
   wire n248499;
   wire n248500;
   wire n248501;
   wire n248502;
   wire n248503;
   wire n248504;
   wire n248505;
   wire n248506;
   wire n248507;
   wire n248508;
   wire n248509;
   wire n248510;
   wire n248511;
   wire n248512;
   wire n248513;
   wire n248514;
   wire n248515;
   wire n248516;
   wire n248517;
   wire n248518;
   wire n248519;
   wire n248520;
   wire n248521;
   wire n248522;
   wire n248523;
   wire n248524;
   wire n248525;
   wire n248526;
   wire n248527;
   wire n248528;
   wire n248529;
   wire n248530;
   wire n248531;
   wire n248532;
   wire n248533;
   wire n248534;
   wire n248535;
   wire n248536;
   wire n248537;
   wire n248538;
   wire n248539;
   wire n248540;
   wire n248541;
   wire n248542;
   wire n248543;
   wire n248544;
   wire n248545;
   wire n248546;
   wire n248547;
   wire n248548;
   wire n248549;
   wire n248550;
   wire n248551;
   wire n248552;
   wire n248553;
   wire n248554;
   wire n248555;
   wire n248556;
   wire n248557;
   wire n248558;
   wire n248559;
   wire n248560;
   wire n248561;
   wire n248562;
   wire n248563;
   wire n248564;
   wire n248565;
   wire n248566;
   wire n248567;
   wire n248568;
   wire n248569;
   wire n248570;
   wire n248571;
   wire n248572;
   wire n248573;
   wire n248574;
   wire n248575;
   wire n248576;
   wire n248577;
   wire n248578;
   wire n248579;
   wire n248580;
   wire n248581;
   wire n248582;
   wire n248583;
   wire n248584;
   wire n248585;
   wire n248586;
   wire n248587;
   wire n248588;
   wire n248589;
   wire n248590;
   wire n248591;
   wire n248592;
   wire n248593;
   wire n248594;
   wire n248595;
   wire n248596;
   wire n248597;
   wire n248598;
   wire n248599;
   wire n248600;
   wire n248601;
   wire n248602;
   wire n248603;
   wire n248604;
   wire n248605;
   wire n248606;
   wire n248607;
   wire n248608;
   wire n248609;
   wire n248610;
   wire n248611;
   wire n248612;
   wire n248613;
   wire n248614;
   wire n248615;
   wire n248616;
   wire n248617;
   wire n248618;
   wire n248619;
   wire n248620;
   wire n248621;
   wire n248622;
   wire n248623;
   wire n248624;
   wire n248625;
   wire n248626;
   wire n248627;
   wire n248628;
   wire n248629;
   wire n248630;
   wire n248631;
   wire n248632;
   wire n248633;
   wire n248634;
   wire n248635;
   wire n248636;
   wire n248637;
   wire n248638;
   wire n248639;
   wire n248640;
   wire n248641;
   wire n248642;
   wire n248643;
   wire n248644;
   wire n248645;
   wire n248646;
   wire n248647;
   wire n248648;
   wire n248649;
   wire n248650;
   wire n248651;
   wire n248652;
   wire n248653;
   wire n248654;
   wire n248655;
   wire n248656;
   wire n248657;
   wire n248658;
   wire n248659;
   wire n248660;
   wire n248661;
   wire n248662;
   wire n248663;
   wire n248664;
   wire n248665;
   wire n248666;
   wire n248667;
   wire n248668;
   wire n248669;
   wire n248670;
   wire n248671;
   wire n248672;
   wire n248673;
   wire n248674;
   wire n248675;
   wire n248676;
   wire n248677;
   wire n248678;
   wire n248679;
   wire n248680;
   wire n248681;
   wire n248682;
   wire n248683;
   wire n248684;
   wire n248685;
   wire n248686;
   wire n248687;
   wire n248688;
   wire n248689;
   wire n248690;
   wire n248691;
   wire n248692;
   wire n248693;
   wire n248694;
   wire n248695;
   wire n248696;
   wire n248697;
   wire n248698;
   wire n248699;
   wire n248700;
   wire n248701;
   wire n248702;
   wire n248703;
   wire n248704;
   wire n248705;
   wire n248706;
   wire n248707;
   wire n248708;
   wire n248709;
   wire n248710;
   wire n248711;
   wire n248712;
   wire n248713;
   wire n248714;
   wire n248715;
   wire n248716;
   wire n248717;
   wire n248718;
   wire n248719;
   wire n248720;
   wire n248721;
   wire n248722;
   wire n248723;
   wire n248724;
   wire n248725;
   wire n248726;
   wire n248727;
   wire n248728;
   wire n248729;
   wire n248730;
   wire n248731;
   wire n248732;
   wire n248733;
   wire n248734;
   wire n248735;
   wire n248736;
   wire n248737;
   wire n248738;
   wire n248739;
   wire n248740;
   wire n248741;
   wire n248742;
   wire n248743;
   wire n248744;
   wire n248745;
   wire n248746;
   wire n248747;
   wire n248748;
   wire n248749;
   wire n248750;
   wire n248751;
   wire n248752;
   wire n248753;
   wire n248754;
   wire n248755;
   wire n248756;
   wire n248757;
   wire n248758;
   wire n248759;
   wire n248760;
   wire n248761;
   wire n248762;
   wire n248763;
   wire n248764;
   wire n248765;
   wire n248766;
   wire n248767;
   wire n248768;
   wire n248769;
   wire n248770;
   wire n248771;
   wire n248772;
   wire n248773;
   wire n248774;
   wire n248775;
   wire n248776;
   wire n248777;
   wire n248778;
   wire n248779;
   wire n248780;
   wire n248781;
   wire n248782;
   wire n248783;
   wire n248784;
   wire n248785;
   wire n248786;
   wire n248787;
   wire n248788;
   wire n248789;
   wire n248790;
   wire n248791;
   wire n248792;
   wire n248793;
   wire n248794;
   wire n248795;
   wire n248796;
   wire n248797;
   wire n248798;
   wire n248799;
   wire n248800;
   wire n248801;
   wire n248802;
   wire n248803;
   wire n248804;
   wire n248805;
   wire n248806;
   wire n248807;
   wire n248808;
   wire n248809;
   wire n248810;
   wire n248811;
   wire n248812;
   wire n248813;
   wire n248814;
   wire n248815;
   wire n248816;
   wire n248817;
   wire n248818;
   wire n248819;
   wire n248820;
   wire n248821;
   wire n248822;
   wire n248823;
   wire n248824;
   wire n248825;
   wire n248826;
   wire n248827;
   wire n248828;
   wire n248829;
   wire n248830;
   wire n248831;
   wire n248832;
   wire n248833;
   wire n248834;
   wire n248835;
   wire n248836;
   wire n248837;
   wire n248838;
   wire n248839;
   wire n248840;
   wire n248841;
   wire n248842;
   wire n248843;
   wire n248844;
   wire n248845;
   wire n248854;
   wire n248855;
   wire n248856;
   wire n248857;
   wire n248866;
   wire n248867;
   wire n248868;
   wire n248869;
   wire n248878;
   wire n248879;
   wire n248880;
   wire n248881;
   wire n248890;
   wire n248891;
   wire n248892;
   wire n248893;
   wire n248894;
   wire n248895;
   wire n248896;
   wire n248897;
   wire n248906;
   wire n248907;
   wire n248908;
   wire n248909;
   wire n248918;
   wire n248919;
   wire n248920;
   wire n248921;
   wire n248930;
   wire n248931;
   wire n248932;
   wire n248933;
   wire n248942;
   wire n248943;
   wire n248944;
   wire n248945;
   wire n248946;
   wire n248947;
   wire n248948;
   wire n248949;
   wire n248950;
   wire n248951;
   wire n248952;
   wire n248953;
   wire n248954;
   wire n248955;
   wire n248956;
   wire n248957;
   wire n248958;
   wire n248959;
   wire n248960;
   wire n248961;
   wire n248962;
   wire n248963;
   wire n248964;
   wire n248965;
   wire n248966;
   wire n248967;
   wire n248968;
   wire n248969;
   wire n248970;
   wire n248971;
   wire n248972;
   wire n248973;
   wire n248974;
   wire n248975;
   wire n248976;
   wire n248977;
   wire n248978;
   wire n248980;
   wire n248981;
   wire n248982;
   wire n248983;
   wire n248984;
   wire n248985;
   wire n248986;
   wire n248987;
   wire n248988;
   wire n248989;
   wire n248990;
   wire n248991;
   wire n248992;
   wire n248993;
   wire n248994;
   wire n248995;
   wire n248996;
   wire n248997;
   wire n248998;
   wire n248999;
   wire n249000;
   wire n249001;
   wire n249002;
   wire n249003;
   wire n249004;
   wire n249005;
   wire n249006;
   wire n249007;
   wire n249008;
   wire n249009;
   wire n249010;
   wire n249011;
   wire n249012;
   wire n249013;
   wire n249014;
   wire n249015;
   wire n249016;
   wire n249017;
   wire n249018;
   wire n249019;
   wire n249020;
   wire n249021;
   wire n249022;
   wire n249023;
   wire n249024;
   wire n249025;
   wire n249026;
   wire n249027;
   wire n249028;
   wire n249029;
   wire n249030;
   wire n249031;
   wire n249032;
   wire n249033;
   wire n249034;
   wire n249035;
   wire n249036;
   wire n249037;
   wire n249038;
   wire n249039;
   wire n249040;
   wire n249041;
   wire n249042;
   wire n249043;
   wire n249044;
   wire n249045;
   wire n249046;
   wire n249047;
   wire n249048;
   wire n249049;
   wire n249051;
   wire n249052;
   wire n249053;
   wire n249055;
   wire n249056;
   wire n249057;
   wire n249058;
   wire n249060;
   wire n249061;
   wire n249062;
   wire n249063;
   wire n249064;
   wire n249065;
   wire n249066;
   wire n249067;
   wire n249068;
   wire n249069;
   wire n249070;
   wire n249071;
   wire n249072;
   wire n249073;
   wire n249074;
   wire n249075;
   wire n249077;
   wire n249078;
   wire n249079;
   wire n249080;
   wire n249081;
   wire n249082;
   wire n249083;
   wire n249084;
   wire n249085;
   wire n249086;
   wire n249087;
   wire n249088;
   wire n249089;
   wire n249090;
   wire n249091;
   wire n249092;
   wire n249093;
   wire n249094;
   wire n249095;
   wire n249096;
   wire n249097;
   wire n249098;
   wire n249099;
   wire n249100;
   wire n249101;
   wire n249102;
   wire n249103;
   wire n249104;
   wire n249105;
   wire n249106;
   wire n249107;
   wire n249108;
   wire n249109;
   wire n249110;
   wire n249111;
   wire n249112;
   wire n249113;
   wire n249114;
   wire n249115;
   wire n249116;
   wire n249117;
   wire n249118;
   wire n249119;
   wire n249120;
   wire n249121;
   wire n249122;
   wire n249123;
   wire n249124;
   wire n249125;
   wire n249126;
   wire n249127;
   wire n249128;
   wire n249129;
   wire n249130;
   wire n249131;
   wire n249132;
   wire n249133;
   wire n249134;
   wire n249135;
   wire n249136;
   wire n249137;
   wire n249138;
   wire n249140;
   wire n249141;
   wire n249142;
   wire n249143;
   wire n249144;
   wire n249145;
   wire n249146;
   wire n249147;
   wire n249148;
   wire n249149;
   wire n249150;
   wire n249151;
   wire n249152;
   wire n249153;
   wire n249154;
   wire n249155;
   wire n249156;
   wire n249157;
   wire n249158;
   wire n249159;
   wire n249160;
   wire n249161;
   wire n249162;
   wire n249163;
   wire n249164;
   wire n249165;
   wire n249166;
   wire n249167;
   wire n249168;
   wire n249169;
   wire n249170;
   wire n249171;
   wire n249172;
   wire n249173;
   wire n249174;
   wire n249175;
   wire n249176;
   wire n249177;
   wire n249178;
   wire n249179;
   wire n249181;
   wire n249182;
   wire n249183;
   wire n249184;
   wire n249185;
   wire n249186;
   wire n249187;
   wire n249188;
   wire n249189;
   wire n249190;
   wire n249191;
   wire n249192;
   wire n249193;
   wire n249194;
   wire n249195;
   wire n249196;
   wire n249197;
   wire n249198;
   wire n249199;
   wire n249200;
   wire n249201;
   wire n249202;
   wire n249203;
   wire n249204;
   wire n249205;
   wire n249206;
   wire n249207;
   wire n249208;
   wire n249209;
   wire n249210;
   wire n249211;
   wire n249212;
   wire n249213;
   wire n249214;
   wire n249215;
   wire n249216;
   wire n249217;
   wire n249218;
   wire n249219;
   wire n249220;
   wire n249221;
   wire n249222;
   wire n249223;
   wire n249224;
   wire n249225;
   wire n249226;
   wire n249227;
   wire n249228;
   wire n249229;
   wire n249230;
   wire n249231;
   wire n249232;
   wire n249233;
   wire n249234;
   wire n249235;
   wire n249236;
   wire n249237;
   wire n249238;
   wire n249239;
   wire n249240;
   wire n249241;
   wire n249242;
   wire n249244;
   wire n249246;
   wire n249247;
   wire n249248;
   wire n249249;
   wire n249250;
   wire n249251;
   wire n249252;
   wire n249253;
   wire n249254;
   wire n249255;
   wire n249256;
   wire n249257;
   wire n249258;
   wire n249259;
   wire n249260;
   wire n249261;
   wire n249262;
   wire n249263;
   wire n249264;
   wire n249265;
   wire n249266;
   wire n249267;
   wire n249268;
   wire n249269;
   wire n249270;
   wire n249271;
   wire n249272;
   wire n249273;
   wire n249274;
   wire n249275;
   wire n249276;
   wire n249277;
   wire n249278;
   wire n249279;
   wire n249280;
   wire n249281;
   wire n249282;
   wire n249283;
   wire n249284;
   wire n249285;
   wire n249286;
   wire n249287;
   wire n249288;
   wire n249289;
   wire n249290;
   wire n249291;
   wire n249292;
   wire n249293;
   wire n249294;
   wire n249295;
   wire n249296;
   wire n249297;
   wire n249298;
   wire n249299;
   wire n249300;
   wire n249301;
   wire n249302;
   wire n249303;
   wire n249304;
   wire n249305;
   wire n249306;
   wire n249307;
   wire n249308;
   wire n249309;
   wire n249310;
   wire n249311;
   wire n249312;
   wire n249313;
   wire n249314;
   wire n249315;
   wire n249316;
   wire n249317;
   wire n249318;
   wire n249319;
   wire n249320;
   wire n249321;
   wire n249322;
   wire n249323;
   wire n249324;
   wire n249325;
   wire n249326;
   wire n249327;
   wire n249328;
   wire n249329;
   wire n249330;
   wire n249331;
   wire n249332;
   wire n249333;
   wire n249334;
   wire n249335;
   wire n249336;
   wire n249337;
   wire n249338;
   wire n249339;
   wire n249340;
   wire n249341;
   wire n249342;
   wire n249343;
   wire n249344;
   wire n249345;
   wire n249346;
   wire n249347;
   wire n249348;
   wire n249349;
   wire n249350;
   wire n249351;
   wire n249352;
   wire n249353;
   wire n249354;
   wire n249355;
   wire n249356;
   wire n249357;
   wire n249358;
   wire n249359;
   wire n249360;
   wire n249361;
   wire n249362;
   wire n249363;
   wire n249364;
   wire n249365;
   wire n249366;
   wire n249367;
   wire n249368;
   wire n249369;
   wire n249370;
   wire n249371;
   wire n249372;
   wire n249373;
   wire n249374;
   wire n249375;
   wire n249376;
   wire n249377;
   wire n249378;
   wire n249379;
   wire n249380;
   wire n249381;
   wire n249382;
   wire n249383;
   wire n249384;
   wire n249385;
   wire n249386;
   wire n249387;
   wire n249388;
   wire n249389;
   wire n249390;
   wire n249391;
   wire n249392;
   wire n249393;
   wire n249394;
   wire n249395;
   wire n249396;
   wire n249397;
   wire n249398;
   wire n249399;
   wire n249400;
   wire n249401;
   wire n249402;
   wire n249403;
   wire n249404;
   wire n249405;
   wire n249406;
   wire n249407;
   wire n249408;
   wire n249409;
   wire n249410;
   wire n249411;
   wire n249412;
   wire n249413;
   wire n249414;
   wire n249415;
   wire n249416;
   wire n249417;
   wire n249418;
   wire n249419;
   wire n249420;
   wire n249421;
   wire n249422;
   wire n249423;
   wire n249424;
   wire n249425;
   wire n249426;
   wire n249427;
   wire n249428;
   wire n249429;
   wire n249430;
   wire n249431;
   wire n249432;
   wire n249433;
   wire n249434;
   wire n249435;
   wire n249436;
   wire n249437;
   wire n249438;
   wire n249439;
   wire n249440;
   wire n249441;
   wire n249442;
   wire n249443;
   wire n249444;
   wire n249445;
   wire n249446;
   wire n249447;
   wire n249448;
   wire n249449;
   wire n249450;
   wire n249451;
   wire n249452;
   wire n249453;
   wire n249454;
   wire n249455;
   wire n249456;
   wire n249457;
   wire n249458;
   wire n249459;
   wire n249460;
   wire n249461;
   wire n249462;
   wire n249463;
   wire n249464;
   wire n249465;
   wire n249466;
   wire n249467;
   wire n249468;
   wire n249469;
   wire n249470;
   wire n249471;
   wire n249472;
   wire n249473;
   wire n249474;
   wire n249475;
   wire n249476;
   wire n249477;
   wire n249478;
   wire n249479;
   wire n249480;
   wire n249481;
   wire n249482;
   wire n249483;
   wire n249484;
   wire n249485;
   wire n249486;
   wire n249487;
   wire n249488;
   wire n249489;
   wire n249490;
   wire n249491;
   wire n249492;
   wire n249493;
   wire n249494;
   wire n249495;
   wire n249496;
   wire n249497;
   wire n249498;
   wire n249499;
   wire n249500;
   wire n249501;
   wire n249502;
   wire n249503;
   wire n249504;
   wire n249505;
   wire n249506;
   wire n249507;
   wire n249508;
   wire n249509;
   wire n249510;
   wire n249511;
   wire n249512;
   wire n249513;
   wire n249514;
   wire n249515;
   wire n249516;
   wire n249517;
   wire n249518;
   wire n249519;
   wire n249520;
   wire n249521;
   wire n249522;
   wire n249523;
   wire n249524;
   wire n249525;
   wire n249526;
   wire n249527;
   wire n249528;
   wire n249529;
   wire n249530;
   wire n249531;
   wire n249532;
   wire n249533;
   wire n249534;
   wire n249535;
   wire n249536;
   wire n249537;
   wire n249538;
   wire n249539;
   wire n249540;
   wire n249541;
   wire n249542;
   wire n249543;
   wire n249544;
   wire n249545;
   wire n249546;
   wire n249547;
   wire n249548;
   wire n249549;
   wire n249550;
   wire n249551;
   wire n249552;
   wire n249553;
   wire n249554;
   wire n249555;
   wire n249556;
   wire n249557;
   wire n249558;
   wire n249559;
   wire n249560;
   wire n249561;
   wire n249562;
   wire n249563;
   wire n249564;
   wire n249565;
   wire n249566;
   wire n249567;
   wire n249568;
   wire n249569;
   wire n249570;
   wire n249571;
   wire n249572;
   wire n249573;
   wire n249574;
   wire n249575;
   wire n249576;
   wire n249577;
   wire n249578;
   wire n249579;
   wire n249580;
   wire n249581;
   wire n249582;
   wire n249583;
   wire n249584;
   wire n249585;
   wire n249586;
   wire n249587;
   wire n249588;
   wire n249589;
   wire n249590;
   wire n249591;
   wire n249592;
   wire n249593;
   wire n249594;
   wire n249595;
   wire n249596;
   wire n249597;
   wire n249598;
   wire n249599;
   wire n249600;
   wire n249601;
   wire n249602;
   wire n249603;
   wire n249604;
   wire n249605;
   wire n249606;
   wire n249607;
   wire n249608;
   wire n249609;
   wire n249610;
   wire n249611;
   wire n249612;
   wire n249613;
   wire n249614;
   wire n249615;
   wire n249616;
   wire n249617;
   wire n249618;
   wire n249619;
   wire n249620;
   wire n249621;
   wire n249622;
   wire n249623;
   wire n249624;
   wire n249625;
   wire n249626;
   wire n249627;
   wire n249628;
   wire n249629;
   wire n249630;
   wire n249631;
   wire n249632;
   wire n249633;
   wire n249634;
   wire n249635;
   wire n249636;
   wire n249637;
   wire n249638;
   wire n249639;
   wire n249640;
   wire n249641;
   wire n249642;
   wire n249643;
   wire n249644;
   wire n249645;
   wire n249646;
   wire n249647;
   wire n249648;
   wire n249649;
   wire n249651;
   wire n249652;
   wire n249653;
   wire n249654;
   wire n249655;
   wire n249656;
   wire n249657;
   wire n249658;
   wire n249659;
   wire n249660;
   wire n249661;
   wire n249662;
   wire n249663;
   wire n249664;
   wire n249665;
   wire n249666;
   wire n249667;
   wire n249668;
   wire n249669;
   wire n249670;
   wire n249671;
   wire n249672;
   wire n249673;
   wire n249674;
   wire n249675;
   wire n249676;
   wire n249677;
   wire n249678;
   wire n249679;
   wire n249680;
   wire n249681;
   wire n249682;
   wire n249683;
   wire n249684;
   wire n249685;
   wire n249686;
   wire n249687;
   wire n249688;
   wire n249689;
   wire n249690;
   wire n249691;
   wire n249692;
   wire n249693;
   wire n249694;
   wire n249695;
   wire n249696;
   wire n249697;
   wire n249698;
   wire n249699;
   wire n249700;
   wire n249701;
   wire n249702;
   wire n249703;
   wire n249704;
   wire n249705;
   wire n249706;
   wire n249707;
   wire n249708;
   wire n249709;
   wire n249710;
   wire n249711;
   wire n249712;
   wire n249713;
   wire n249714;
   wire n249715;
   wire n249716;
   wire n249717;
   wire n249718;
   wire n249719;
   wire n249720;
   wire n249721;
   wire n249722;
   wire n249723;
   wire n249724;
   wire n249725;
   wire n249726;
   wire n249727;
   wire n249728;
   wire n249729;
   wire n249730;
   wire n249731;
   wire n249732;
   wire n249733;
   wire n249734;
   wire n249735;
   wire n249736;
   wire n249737;
   wire n249738;
   wire n249739;
   wire n249740;
   wire n249741;
   wire n249742;
   wire n249743;
   wire n249744;
   wire n249745;
   wire n249746;
   wire n249747;
   wire n249748;
   wire n249749;
   wire n249750;
   wire n249751;
   wire n249752;
   wire n249753;
   wire n249754;
   wire n249755;
   wire n249756;
   wire n249757;
   wire n249758;
   wire n249759;
   wire n249760;
   wire n249761;
   wire n249762;
   wire n249763;
   wire n249764;
   wire n249765;
   wire n249766;
   wire n249767;
   wire n249768;
   wire n249769;
   wire n249770;
   wire n249771;
   wire n249772;
   wire n249773;
   wire n249774;
   wire n249775;
   wire n249776;
   wire n249777;
   wire n249778;
   wire n249779;
   wire n249780;
   wire n249781;
   wire n249782;
   wire n249783;
   wire n249784;
   wire n249785;
   wire n249786;
   wire n249787;
   wire n249788;
   wire n249789;
   wire n249791;
   wire n249792;
   wire n249793;
   wire n249794;
   wire n249795;
   wire n249796;
   wire n249797;
   wire n249798;
   wire n249799;
   wire n249800;
   wire n249801;
   wire n249802;
   wire n249803;
   wire n249804;
   wire n249805;
   wire n249806;
   wire n249807;
   wire n249808;
   wire n249809;
   wire n249810;
   wire n249811;
   wire n249812;
   wire n249813;
   wire n249815;
   wire n249816;
   wire n249817;
   wire n249818;
   wire n249819;
   wire n249820;
   wire n249821;
   wire n249822;
   wire n249823;
   wire n249824;
   wire n249825;
   wire n249826;
   wire n249827;
   wire n249828;
   wire n249829;
   wire n249830;
   wire n249831;
   wire n249832;
   wire n249833;
   wire n249834;
   wire n249835;
   wire n249836;
   wire n249838;
   wire n249841;
   wire n249842;
   wire n249843;
   wire n249844;
   wire n249845;
   wire n249846;
   wire n249847;
   wire n249848;
   wire n249849;
   wire n249850;
   wire n249851;
   wire n249852;
   wire n249853;
   wire n249854;
   wire n249855;
   wire n249856;
   wire n249857;
   wire n249858;
   wire n249859;
   wire n249860;
   wire n249861;
   wire n249862;
   wire n249863;
   wire n249864;
   wire n249865;
   wire n249866;
   wire n249867;
   wire n249868;
   wire n249869;
   wire n249870;
   wire n249871;
   wire n249872;
   wire n249873;
   wire n249874;
   wire n249875;
   wire n249876;
   wire n249877;
   wire n249878;
   wire n249879;
   wire n249880;
   wire n249881;
   wire n249882;
   wire n249883;
   wire n249884;
   wire n249885;
   wire n249886;
   wire n249887;
   wire n249888;
   wire n249889;
   wire n249890;
   wire n249891;
   wire n249892;
   wire n249893;
   wire n249894;
   wire n249895;
   wire n249896;
   wire n249897;
   wire n249898;
   wire n249899;
   wire n249900;
   wire n249901;
   wire n249902;
   wire n249903;
   wire n249904;
   wire n249905;
   wire n249906;
   wire n249907;
   wire n249908;
   wire n249909;
   wire n249910;
   wire n249911;
   wire n249912;
   wire n249913;
   wire n249914;
   wire n249915;
   wire n249916;
   wire n249917;
   wire n249918;
   wire n249919;
   wire n249920;
   wire n249921;
   wire n249922;
   wire n249923;
   wire n249924;
   wire n249925;
   wire n249926;
   wire n249927;
   wire n249928;
   wire n249929;
   wire n249930;
   wire n249931;
   wire n249932;
   wire n249933;
   wire n249934;
   wire n249935;
   wire n249936;
   wire n249937;
   wire n249938;
   wire n249939;
   wire n249940;
   wire n249941;
   wire n249942;
   wire n249943;
   wire n249944;
   wire n249945;
   wire n249946;
   wire n249947;
   wire n249948;
   wire n249949;
   wire n249950;
   wire n249951;
   wire n249952;
   wire n249953;
   wire n249954;
   wire n249955;
   wire n249956;
   wire n249957;
   wire n249958;
   wire n249959;
   wire n249960;
   wire n249961;
   wire n249962;
   wire n249963;
   wire n249964;
   wire n249965;
   wire n249966;
   wire n249967;
   wire n249968;
   wire n249969;
   wire n249970;
   wire n249971;
   wire n249972;
   wire n249973;
   wire n249974;
   wire n249976;
   wire n249977;
   wire n249978;
   wire n249979;
   wire n249980;
   wire n249981;
   wire n249982;
   wire n249983;
   wire n249984;
   wire n249985;
   wire n249986;
   wire n249987;
   wire n249988;
   wire n249989;
   wire n249990;
   wire n249991;
   wire n249992;
   wire n249993;
   wire n249994;
   wire n249995;
   wire n249996;
   wire n249997;
   wire n249998;
   wire n249999;
   wire n250000;
   wire n250001;
   wire n250002;
   wire n250003;
   wire n250004;
   wire n250005;
   wire n250006;
   wire n250007;
   wire n250008;
   wire n250009;
   wire n250011;
   wire n250012;
   wire n250013;
   wire n250014;
   wire n250015;
   wire n250016;
   wire n250018;
   wire n250019;
   wire n250020;
   wire n250021;
   wire n250022;
   wire n250023;
   wire n250024;
   wire n250025;
   wire n250026;
   wire n250027;
   wire n250028;
   wire n250029;
   wire n250030;
   wire n250031;
   wire n250032;
   wire n250033;
   wire n250034;
   wire n250035;
   wire n250036;
   wire n250037;
   wire n250038;
   wire n250039;
   wire n250040;
   wire n250041;
   wire n250042;
   wire n250043;
   wire n250044;
   wire n250045;
   wire n250047;
   wire n250048;
   wire n250049;
   wire n250050;
   wire n250051;
   wire n250052;
   wire n250053;
   wire n250054;
   wire n250055;
   wire n250056;
   wire n250057;
   wire n250058;
   wire n250059;
   wire n250060;
   wire n250061;
   wire n250062;
   wire n250063;
   wire n250064;
   wire n250065;
   wire n250066;
   wire n250067;
   wire n250068;
   wire n250069;
   wire n250070;
   wire n250071;
   wire n250072;
   wire n250073;
   wire n250074;
   wire n250075;
   wire n250076;
   wire n250077;
   wire n250078;
   wire n250079;
   wire n250080;
   wire n250081;
   wire n250083;
   wire n250084;
   wire n250085;
   wire n250086;
   wire n250087;
   wire n250088;
   wire n250089;
   wire n250090;
   wire n250092;
   wire n250093;
   wire n250094;
   wire n250095;
   wire n250096;
   wire n250097;
   wire n250098;
   wire n250099;
   wire n250100;
   wire n250101;
   wire n250102;
   wire n250103;
   wire n250104;
   wire n250105;
   wire n250106;
   wire n250107;
   wire n250108;
   wire n250109;
   wire n250110;
   wire n250111;
   wire n250112;
   wire n250113;
   wire n250114;
   wire n250115;
   wire n250116;
   wire n250117;
   wire n250119;
   wire n250120;
   wire n250121;
   wire n250122;
   wire n250123;
   wire n250124;
   wire n250126;
   wire n250127;
   wire n250128;
   wire n250129;
   wire n250130;
   wire n250131;
   wire n250132;
   wire n250133;
   wire n250134;
   wire n250135;
   wire n250136;
   wire n250137;
   wire n250138;
   wire n250139;
   wire n250140;
   wire n250141;
   wire n250142;
   wire n250143;
   wire n250144;
   wire n250145;
   wire n250146;
   wire n250147;
   wire n250148;
   wire n250149;
   wire n250150;
   wire n250151;
   wire n250152;
   wire n250153;
   wire n250154;
   wire n250156;
   wire n250157;
   wire n250158;
   wire n250159;
   wire n250160;
   wire n250161;
   wire n250162;
   wire n250163;
   wire n250164;
   wire n250165;
   wire n250166;
   wire n250167;
   wire n250168;
   wire n250169;
   wire n250170;
   wire n250171;
   wire n250172;
   wire n250173;
   wire n250174;
   wire n250175;
   wire n250176;
   wire n250177;
   wire n250178;
   wire n250179;
   wire n250180;
   wire n250181;
   wire n250182;
   wire n250183;
   wire n250184;
   wire n250185;
   wire n250186;
   wire n250187;
   wire n250188;
   wire n250189;
   wire n250190;
   wire n250192;
   wire n250193;
   wire n250194;
   wire n250195;
   wire n250196;
   wire n250197;
   wire n250198;
   wire n250199;
   wire n250200;
   wire n250201;
   wire n250202;
   wire n250203;
   wire n250204;
   wire n250205;
   wire n250206;
   wire n250207;
   wire n250208;
   wire n250209;
   wire n250210;
   wire n250211;
   wire n250212;
   wire n250213;
   wire n250214;
   wire n250215;
   wire n250216;
   wire n250217;
   wire n250218;
   wire n250219;
   wire n250220;
   wire n250221;
   wire n250222;
   wire n250223;
   wire n250224;
   wire n250225;
   wire n250226;
   wire n250227;
   wire n250228;
   wire n250230;
   wire n250231;
   wire n250232;
   wire n250233;
   wire n250234;
   wire n250235;
   wire n250237;
   wire n250238;
   wire n250239;
   wire n250240;
   wire n250241;
   wire n250242;
   wire n250243;
   wire n250244;
   wire n250245;
   wire n250246;
   wire n250247;
   wire n250248;
   wire n250249;
   wire n250250;
   wire n250251;
   wire n250252;
   wire n250253;
   wire n250254;
   wire n250255;
   wire n250256;
   wire n250257;
   wire n250258;
   wire n250259;
   wire n250260;
   wire n250261;
   wire n250262;
   wire n250263;
   wire n250264;
   wire n250266;
   wire n250267;
   wire n250268;
   wire n250269;
   wire n250270;
   wire n250271;
   wire n250272;
   wire n250273;
   wire n250274;
   wire n250275;
   wire n250276;
   wire n250277;
   wire n250278;
   wire n250279;
   wire n250280;
   wire n250281;
   wire n250282;
   wire n250283;
   wire n250284;
   wire n250285;
   wire n250286;
   wire n250287;
   wire n250288;
   wire n250289;
   wire n250290;
   wire n250291;
   wire n250292;
   wire n250293;
   wire n250294;
   wire n250295;
   wire n250296;
   wire n250297;
   wire n250298;
   wire n250299;
   wire n250301;
   wire n250302;
   wire n250303;
   wire n250304;
   wire n250305;
   wire n250306;
   wire n250307;
   wire n250308;
   wire n250309;
   wire n250310;
   wire n250311;
   wire n250312;
   wire n250313;
   wire n250314;
   wire n250315;
   wire n250316;
   wire n250317;
   wire n250318;
   wire n250319;
   wire n250320;
   wire n250321;
   wire n250322;
   wire n250323;
   wire n250324;
   wire n250325;
   wire n250326;
   wire n250327;
   wire n250328;
   wire n250329;
   wire n250330;
   wire n250331;
   wire n250332;
   wire n250333;
   wire n250334;
   wire n250336;
   wire n250337;
   wire n250338;
   wire n250339;
   wire n250340;
   wire n250341;
   wire n250343;
   wire n250344;
   wire n250345;
   wire n250346;
   wire n250347;
   wire n250348;
   wire n250349;
   wire n250350;
   wire n250351;
   wire n250352;
   wire n250353;
   wire n250354;
   wire n250355;
   wire n250356;
   wire n250357;
   wire n250358;
   wire n250359;
   wire n250360;
   wire n250361;
   wire n250362;
   wire n250363;
   wire n250364;
   wire n250365;
   wire n250366;
   wire n250367;
   wire n250368;
   wire n250369;
   wire n250370;
   wire n250372;
   wire n250373;
   wire n250374;
   wire n250375;
   wire n250376;
   wire n250377;
   wire n250378;
   wire n250379;
   wire n250380;
   wire n250381;
   wire n250382;
   wire n250383;
   wire n250384;
   wire n250385;
   wire n250386;
   wire n250387;
   wire n250388;
   wire n250389;
   wire n250390;
   wire n250391;
   wire n250392;
   wire n250393;
   wire n250394;
   wire n250395;
   wire n250396;
   wire n250397;
   wire n250398;
   wire n250399;
   wire n250400;
   wire n250401;
   wire n250402;
   wire n250403;
   wire n250404;
   wire n250405;
   wire n250407;
   wire n250408;
   wire n250409;
   wire n250410;
   wire n250411;
   wire n250412;
   wire n250413;
   wire n250414;
   wire n250415;
   wire n250416;
   wire n250417;
   wire n250418;
   wire n250419;
   wire n250420;
   wire n250421;
   wire n250422;
   wire n250423;
   wire n250424;
   wire n250425;
   wire n250426;
   wire n250427;
   wire n250428;
   wire n250429;
   wire n250430;
   wire n250431;
   wire n250432;
   wire n250433;
   wire n250434;
   wire n250435;
   wire n250436;
   wire n250437;
   wire n250438;
   wire n250439;
   wire n250440;
   wire n250442;
   wire n250443;
   wire n250444;
   wire n250445;
   wire n250446;
   wire n250447;
   wire n250449;
   wire n250450;
   wire n250451;
   wire n250452;
   wire n250453;
   wire n250454;
   wire n250455;
   wire n250456;
   wire n250457;
   wire n250458;
   wire n250459;
   wire n250460;
   wire n250461;
   wire n250462;
   wire n250463;
   wire n250464;
   wire n250465;
   wire n250466;
   wire n250467;
   wire n250468;
   wire n250469;
   wire n250470;
   wire n250471;
   wire n250472;
   wire n250473;
   wire n250474;
   wire n250475;
   wire n250476;
   wire n250478;
   wire n250479;
   wire n250480;
   wire n250481;
   wire n250482;
   wire n250483;
   wire n250484;
   wire n250485;
   wire n250486;
   wire n250487;
   wire n250488;
   wire n250489;
   wire n250490;
   wire n250491;
   wire n250492;
   wire n250493;
   wire n250494;
   wire n250495;
   wire n250496;
   wire n250497;
   wire n250498;
   wire n250499;
   wire n250500;
   wire n250501;
   wire n250502;
   wire n250503;
   wire n250504;
   wire n250505;
   wire n250506;
   wire n250507;
   wire n250508;
   wire n250509;
   wire n250510;
   wire n250511;
   wire n250512;
   wire n250514;
   wire n250515;
   wire n250516;
   wire n250517;
   wire n250518;
   wire n250519;
   wire n250520;
   wire n250521;
   wire n250522;
   wire n250523;
   wire n250524;
   wire n250525;
   wire n250526;
   wire n250527;
   wire n250528;
   wire n250529;
   wire n250530;
   wire n250531;
   wire n250532;
   wire n250533;
   wire n250534;
   wire n250535;
   wire n250536;
   wire n250537;
   wire n250538;
   wire n250539;
   wire n250540;
   wire n250541;
   wire n250542;
   wire n250543;
   wire n250544;
   wire n250545;
   wire n250546;
   wire n250547;
   wire n250549;
   wire n250550;
   wire n250551;
   wire n250552;
   wire n250553;
   wire n250554;
   wire n250556;
   wire n250557;
   wire n250558;
   wire n250559;
   wire n250560;
   wire n250561;
   wire n250562;
   wire n250563;
   wire n250564;
   wire n250565;
   wire n250566;
   wire n250567;
   wire n250568;
   wire n250569;
   wire n250570;
   wire n250571;
   wire n250572;
   wire n250573;
   wire n250574;
   wire n250575;
   wire n250576;
   wire n250577;
   wire n250578;
   wire n250579;
   wire n250580;
   wire n250581;
   wire n250582;
   wire n250583;
   wire n250585;
   wire n250586;
   wire n250587;
   wire n250588;
   wire n250589;
   wire n250590;
   wire n250591;
   wire n250592;
   wire n250593;
   wire n250594;
   wire n250595;
   wire n250596;
   wire n250597;
   wire n250598;
   wire n250599;
   wire n250600;
   wire n250601;
   wire n250602;
   wire n250603;
   wire n250604;
   wire n250605;
   wire n250606;
   wire n250607;
   wire n250608;
   wire n250609;
   wire n250610;
   wire n250611;
   wire n250612;
   wire n250613;
   wire n250614;
   wire n250615;
   wire n250616;
   wire n250617;
   wire n250618;
   wire n250620;
   wire n250621;
   wire n250622;
   wire n250623;
   wire n250624;
   wire n250625;
   wire n250626;
   wire n250627;
   wire n250628;
   wire n250629;
   wire n250630;
   wire n250631;
   wire n250632;
   wire n250633;
   wire n250634;
   wire n250635;
   wire n250636;
   wire n250637;
   wire n250638;
   wire n250639;
   wire n250640;
   wire n250641;
   wire n250642;
   wire n250643;
   wire n250644;
   wire n250645;
   wire n250646;
   wire n250647;
   wire n250648;
   wire n250649;
   wire n250650;
   wire n250651;
   wire n250652;
   wire n250653;
   wire n250655;
   wire n250656;
   wire n250657;
   wire n250658;
   wire n250659;
   wire n250660;
   wire n250662;
   wire n250663;
   wire n250664;
   wire n250665;
   wire n250666;
   wire n250667;
   wire n250668;
   wire n250669;
   wire n250670;
   wire n250671;
   wire n250672;
   wire n250673;
   wire n250674;
   wire n250675;
   wire n250676;
   wire n250677;
   wire n250678;
   wire n250679;
   wire n250680;
   wire n250681;
   wire n250682;
   wire n250683;
   wire n250684;
   wire n250685;
   wire n250686;
   wire n250687;
   wire n250688;
   wire n250689;
   wire n250691;
   wire n250692;
   wire n250693;
   wire n250694;
   wire n250695;
   wire n250696;
   wire n250697;
   wire n250698;
   wire n250699;
   wire n250700;
   wire n250701;
   wire n250702;
   wire n250703;
   wire n250704;
   wire n250705;
   wire n250706;
   wire n250707;
   wire n250708;
   wire n250709;
   wire n250710;
   wire n250711;
   wire n250712;
   wire n250713;
   wire n250714;
   wire n250715;
   wire n250716;
   wire n250717;
   wire n250718;
   wire n250719;
   wire n250720;
   wire n250721;
   wire n250722;
   wire n250723;
   wire n250724;
   wire n250726;
   wire n250727;
   wire n250728;
   wire n250729;
   wire n250730;
   wire n250731;
   wire n250732;
   wire n250733;
   wire n250734;
   wire n250735;
   wire n250736;
   wire n250737;
   wire n250738;
   wire n250739;
   wire n250740;
   wire n250741;
   wire n250742;
   wire n250743;
   wire n250744;
   wire n250745;
   wire n250746;
   wire n250747;
   wire n250748;
   wire n250749;
   wire n250750;
   wire n250751;
   wire n250752;
   wire n250753;
   wire n250754;
   wire n250755;
   wire n250756;
   wire n250757;
   wire n250758;
   wire n250759;
   wire n250761;
   wire n250762;
   wire n250763;
   wire n250764;
   wire n250765;
   wire n250766;
   wire n250768;
   wire n250769;
   wire n250770;
   wire n250771;
   wire n250772;
   wire n250773;
   wire n250774;
   wire n250775;
   wire n250776;
   wire n250777;
   wire n250778;
   wire n250779;
   wire n250780;
   wire n250781;
   wire n250782;
   wire n250783;
   wire n250784;
   wire n250785;
   wire n250786;
   wire n250787;
   wire n250788;
   wire n250789;
   wire n250790;
   wire n250791;
   wire n250792;
   wire n250793;
   wire n250794;
   wire n250795;
   wire n250796;
   wire n250798;
   wire n250799;
   wire n250800;
   wire n250801;
   wire n250802;
   wire n250803;
   wire n250804;
   wire n250805;
   wire n250806;
   wire n250807;
   wire n250808;
   wire n250809;
   wire n250810;
   wire n250811;
   wire n250812;
   wire n250813;
   wire n250814;
   wire n250815;
   wire n250816;
   wire n250817;
   wire n250818;
   wire n250819;
   wire n250820;
   wire n250821;
   wire n250822;
   wire n250823;
   wire n250824;
   wire n250825;
   wire n250826;
   wire n250827;
   wire n250828;
   wire n250829;
   wire n250830;
   wire n250831;
   wire n250833;
   wire n250834;
   wire n250835;
   wire n250836;
   wire n250837;
   wire n250838;
   wire n250839;
   wire n250840;
   wire n250841;
   wire n250842;
   wire n250843;
   wire n250844;
   wire n250845;
   wire n250846;
   wire n250847;
   wire n250848;
   wire n250849;
   wire n250850;
   wire n250851;
   wire n250852;
   wire n250853;
   wire n250854;
   wire n250855;
   wire n250856;
   wire n250857;
   wire n250858;
   wire n250859;
   wire n250860;
   wire n250861;
   wire n250862;
   wire n250863;
   wire n250864;
   wire n250865;
   wire n250866;
   wire n250868;
   wire n250869;
   wire n250870;
   wire n250871;
   wire n250872;
   wire n250873;
   wire n250875;
   wire n250876;
   wire n250877;
   wire n250878;
   wire n250879;
   wire n250880;
   wire n250881;
   wire n250882;
   wire n250883;
   wire n250884;
   wire n250885;
   wire n250886;
   wire n250887;
   wire n250888;
   wire n250889;
   wire n250890;
   wire n250891;
   wire n250892;
   wire n250893;
   wire n250894;
   wire n250895;
   wire n250896;
   wire n250897;
   wire n250898;
   wire n250899;
   wire n250900;
   wire n250901;
   wire n250902;
   wire n250904;
   wire n250905;
   wire n250906;
   wire n250907;
   wire n250908;
   wire n250909;
   wire n250910;
   wire n250911;
   wire n250912;
   wire n250913;
   wire n250914;
   wire n250915;
   wire n250916;
   wire n250917;
   wire n250918;
   wire n250919;
   wire n250920;
   wire n250921;
   wire n250922;
   wire n250923;
   wire n250924;
   wire n250925;
   wire n250926;
   wire n250927;
   wire n250928;
   wire n250929;
   wire n250930;
   wire n250931;
   wire n250932;
   wire n250933;
   wire n250934;
   wire n250935;
   wire n250936;
   wire n250937;
   wire n250939;
   wire n250940;
   wire n250941;
   wire n250942;
   wire n250943;
   wire n250944;
   wire n250945;
   wire n250946;
   wire n250947;
   wire n250948;
   wire n250949;
   wire n250950;
   wire n250951;
   wire n250952;
   wire n250953;
   wire n250954;
   wire n250955;
   wire n250956;
   wire n250957;
   wire n250958;
   wire n250959;
   wire n250960;
   wire n250961;
   wire n250962;
   wire n250963;
   wire n250964;
   wire n250965;
   wire n250966;
   wire n250967;
   wire n250968;
   wire n250969;
   wire n250970;
   wire n250971;
   wire n250972;
   wire n250974;
   wire n250975;
   wire n250976;
   wire n250977;
   wire n250978;
   wire n250979;
   wire n250981;
   wire n250982;
   wire n250983;
   wire n250984;
   wire n250985;
   wire n250986;
   wire n250987;
   wire n250988;
   wire n250989;
   wire n250990;
   wire n250991;
   wire n250992;
   wire n250993;
   wire n250994;
   wire n250995;
   wire n250996;
   wire n250997;
   wire n250998;
   wire n250999;
   wire n251000;
   wire n251001;
   wire n251002;
   wire n251003;
   wire n251004;
   wire n251005;
   wire n251006;
   wire n251007;
   wire n251008;
   wire n251010;
   wire n251011;
   wire n251012;
   wire n251013;
   wire n251014;
   wire n251015;
   wire n251016;
   wire n251017;
   wire n251018;
   wire n251019;
   wire n251020;
   wire n251021;
   wire n251022;
   wire n251023;
   wire n251024;
   wire n251025;
   wire n251026;
   wire n251027;
   wire n251028;
   wire n251029;
   wire n251030;
   wire n251031;
   wire n251032;
   wire n251033;
   wire n251034;
   wire n251035;
   wire n251036;
   wire n251037;
   wire n251038;
   wire n251039;
   wire n251040;
   wire n251041;
   wire n251042;
   wire n251043;
   wire n251045;
   wire n251046;
   wire n251047;
   wire n251048;
   wire n251049;
   wire n251050;
   wire n251051;
   wire n251052;
   wire n251053;
   wire n251054;
   wire n251055;
   wire n251056;
   wire n251057;
   wire n251058;
   wire n251059;
   wire n251060;
   wire n251061;
   wire n251062;
   wire n251063;
   wire n251064;
   wire n251065;
   wire n251066;
   wire n251067;
   wire n251068;
   wire n251069;
   wire n251070;
   wire n251071;
   wire n251072;
   wire n251073;
   wire n251074;
   wire n251075;
   wire n251076;
   wire n251077;
   wire n251078;
   wire n251079;
   wire n251081;
   wire n251082;
   wire n251083;
   wire n251084;
   wire n251085;
   wire n251086;
   wire n251088;
   wire n251089;
   wire n251090;
   wire n251091;
   wire n251092;
   wire n251093;
   wire n251094;
   wire n251095;
   wire n251096;
   wire n251097;
   wire n251098;
   wire n251099;
   wire n251100;
   wire n251101;
   wire n251102;
   wire n251103;
   wire n251104;
   wire n251105;
   wire n251106;
   wire n251107;
   wire n251108;
   wire n251109;
   wire n251110;
   wire n251111;
   wire n251112;
   wire n251113;
   wire n251114;
   wire n251115;
   wire n251117;
   wire n251118;
   wire n251119;
   wire n251120;
   wire n251121;
   wire n251122;
   wire n251123;
   wire n251124;
   wire n251125;
   wire n251126;
   wire n251127;
   wire n251128;
   wire n251129;
   wire n251130;
   wire n251131;
   wire n251132;
   wire n251133;
   wire n251134;
   wire n251135;
   wire n251136;
   wire n251137;
   wire n251138;
   wire n251139;
   wire n251140;
   wire n251141;
   wire n251142;
   wire n251143;
   wire n251144;
   wire n251145;
   wire n251146;
   wire n251147;
   wire n251148;
   wire n251149;
   wire n251150;
   wire n251152;
   wire n251153;
   wire n251154;
   wire n251155;
   wire n251156;
   wire n251157;
   wire n251158;
   wire n251159;
   wire n251160;
   wire n251161;
   wire n251162;
   wire n251163;
   wire n251164;
   wire n251165;
   wire n251166;
   wire n251167;
   wire n251168;
   wire n251169;
   wire n251170;
   wire n251171;
   wire n251172;
   wire n251173;
   wire n251174;
   wire n251175;
   wire n251176;
   wire n251177;
   wire n251178;
   wire n251179;
   wire n251180;
   wire n251181;
   wire n251182;
   wire n251183;
   wire n251184;
   wire n251185;
   wire n251187;
   wire n251188;
   wire n251189;
   wire n251190;
   wire n251191;
   wire n251192;
   wire n251194;
   wire n251195;
   wire n251196;
   wire n251197;
   wire n251198;
   wire n251199;
   wire n251200;
   wire n251201;
   wire n251202;
   wire n251203;
   wire n251204;
   wire n251205;
   wire n251206;
   wire n251207;
   wire n251208;
   wire n251209;
   wire n251210;
   wire n251211;
   wire n251212;
   wire n251213;
   wire n251214;
   wire n251215;
   wire n251216;
   wire n251217;
   wire n251218;
   wire n251219;
   wire n251220;
   wire n251221;
   wire n251223;
   wire n251224;
   wire n251225;
   wire n251226;
   wire n251227;
   wire n251228;
   wire n251229;
   wire n251230;
   wire n251231;
   wire n251232;
   wire n251233;
   wire n251234;
   wire n251235;
   wire n251236;
   wire n251237;
   wire n251238;
   wire n251239;
   wire n251240;
   wire n251241;
   wire n251242;
   wire n251243;
   wire n251244;
   wire n251245;
   wire n251246;
   wire n251247;
   wire n251248;
   wire n251249;
   wire n251250;
   wire n251251;
   wire n251252;
   wire n251253;
   wire n251254;
   wire n251255;
   wire n251256;
   wire n251258;
   wire n251259;
   wire n251260;
   wire n251261;
   wire n251262;
   wire n251263;
   wire n251264;
   wire n251265;
   wire n251266;
   wire n251267;
   wire n251268;
   wire n251269;
   wire n251270;
   wire n251271;
   wire n251272;
   wire n251273;
   wire n251274;
   wire n251275;
   wire n251276;
   wire n251277;
   wire n251278;
   wire n251279;
   wire n251280;
   wire n251281;
   wire n251282;
   wire n251283;
   wire n251284;
   wire n251285;
   wire n251286;
   wire n251287;
   wire n251288;
   wire n251289;
   wire n251290;
   wire n251291;
   wire n251293;
   wire n251294;
   wire n251295;
   wire n251296;
   wire n251297;
   wire n251298;
   wire n251300;
   wire n251301;
   wire n251302;
   wire n251303;
   wire n251304;
   wire n251305;
   wire n251306;
   wire n251307;
   wire n251308;
   wire n251309;
   wire n251310;
   wire n251311;
   wire n251312;
   wire n251313;
   wire n251314;
   wire n251315;
   wire n251316;
   wire n251317;
   wire n251318;
   wire n251319;
   wire n251320;
   wire n251321;
   wire n251322;
   wire n251323;
   wire n251324;
   wire n251325;
   wire n251326;
   wire n251327;
   wire n251329;
   wire n251330;
   wire n251331;
   wire n251332;
   wire n251333;
   wire n251334;
   wire n251335;
   wire n251336;
   wire n251337;
   wire n251338;
   wire n251339;
   wire n251340;
   wire n251341;
   wire n251342;
   wire n251343;
   wire n251344;
   wire n251345;
   wire n251346;
   wire n251347;
   wire n251348;
   wire n251349;
   wire n251350;
   wire n251351;
   wire n251352;
   wire n251353;
   wire n251354;
   wire n251355;
   wire n251356;
   wire n251357;
   wire n251358;
   wire n251359;
   wire n251360;
   wire n251361;
   wire n251362;
   wire n251363;
   wire n251365;
   wire n251366;
   wire n251367;
   wire n251368;
   wire n251369;
   wire n251370;
   wire n251371;
   wire n251372;
   wire n251373;
   wire n251374;
   wire n251375;
   wire n251376;
   wire n251377;
   wire n251378;
   wire n251379;
   wire n251380;
   wire n251381;
   wire n251382;
   wire n251383;
   wire n251384;
   wire n251385;
   wire n251386;
   wire n251387;
   wire n251388;
   wire n251389;
   wire n251390;
   wire n251391;
   wire n251392;
   wire n251393;
   wire n251394;
   wire n251395;
   wire n251396;
   wire n251397;
   wire n251398;
   wire n251400;
   wire n251401;
   wire n251402;
   wire n251403;
   wire n251404;
   wire n251405;
   wire n251407;
   wire n251408;
   wire n251409;
   wire n251410;
   wire n251411;
   wire n251412;
   wire n251413;
   wire n251414;
   wire n251415;
   wire n251416;
   wire n251417;
   wire n251418;
   wire n251419;
   wire n251420;
   wire n251421;
   wire n251422;
   wire n251423;
   wire n251424;
   wire n251425;
   wire n251426;
   wire n251427;
   wire n251428;
   wire n251429;
   wire n251430;
   wire n251431;
   wire n251432;
   wire n251433;
   wire n251434;
   wire n251436;
   wire n251437;
   wire n251438;
   wire n251439;
   wire n251440;
   wire n251441;
   wire n251442;
   wire n251443;
   wire n251444;
   wire n251445;
   wire n251446;
   wire n251447;
   wire n251448;
   wire n251449;
   wire n251450;
   wire n251451;
   wire n251452;
   wire n251453;
   wire n251454;
   wire n251455;
   wire n251456;
   wire n251457;
   wire n251458;
   wire n251459;
   wire n251460;
   wire n251461;
   wire n251462;
   wire n251463;
   wire n251464;
   wire n251465;
   wire n251466;
   wire n251467;
   wire n251468;
   wire n251469;
   wire n251471;
   wire n251472;
   wire n251473;
   wire n251474;
   wire n251475;
   wire n251476;
   wire n251477;
   wire n251478;
   wire n251479;
   wire n251480;
   wire n251481;
   wire n251482;
   wire n251483;
   wire n251484;
   wire n251485;
   wire n251486;
   wire n251487;
   wire n251488;
   wire n251489;
   wire n251490;
   wire n251491;
   wire n251492;
   wire n251493;
   wire n251494;
   wire n251495;
   wire n251496;
   wire n251497;
   wire n251498;
   wire n251499;
   wire n251500;
   wire n251501;
   wire n251502;
   wire n251503;
   wire n251504;
   wire n251506;
   wire n251507;
   wire n251508;
   wire n251509;
   wire n251510;
   wire n251511;
   wire n251513;
   wire n251514;
   wire n251515;
   wire n251516;
   wire n251517;
   wire n251518;
   wire n251519;
   wire n251520;
   wire n251521;
   wire n251522;
   wire n251523;
   wire n251524;
   wire n251525;
   wire n251526;
   wire n251527;
   wire n251528;
   wire n251529;
   wire n251530;
   wire n251531;
   wire n251532;
   wire n251533;
   wire n251534;
   wire n251535;
   wire n251536;
   wire n251537;
   wire n251538;
   wire n251539;
   wire n251540;
   wire n251542;
   wire n251543;
   wire n251544;
   wire n251545;
   wire n251546;
   wire n251547;
   wire n251548;
   wire n251549;
   wire n251550;
   wire n251551;
   wire n251552;
   wire n251553;
   wire n251554;
   wire n251555;
   wire n251556;
   wire n251557;
   wire n251558;
   wire n251559;
   wire n251560;
   wire n251561;
   wire n251562;
   wire n251563;
   wire n251564;
   wire n251565;
   wire n251566;
   wire n251567;
   wire n251568;
   wire n251569;
   wire n251570;
   wire n251571;
   wire n251572;
   wire n251573;
   wire n251574;
   wire n251575;
   wire n251577;
   wire n251578;
   wire n251579;
   wire n251580;
   wire n251581;
   wire n251582;
   wire n251583;
   wire n251584;
   wire n251585;
   wire n251586;
   wire n251587;
   wire n251588;
   wire n251589;
   wire n251590;
   wire n251591;
   wire n251592;
   wire n251593;
   wire n251594;
   wire n251595;
   wire n251596;
   wire n251597;
   wire n251598;
   wire n251599;
   wire n251600;
   wire n251601;
   wire n251602;
   wire n251603;
   wire n251604;
   wire n251605;
   wire n251606;
   wire n251607;
   wire n251608;
   wire n251609;
   wire n251610;
   wire n251612;
   wire n251613;
   wire n251614;
   wire n251615;
   wire n251616;
   wire n251617;
   wire n251619;
   wire n251620;
   wire n251621;
   wire n251622;
   wire n251623;
   wire n251624;
   wire n251625;
   wire n251626;
   wire n251627;
   wire n251628;
   wire n251629;
   wire n251630;
   wire n251631;
   wire n251632;
   wire n251633;
   wire n251634;
   wire n251635;
   wire n251636;
   wire n251637;
   wire n251638;
   wire n251639;
   wire n251640;
   wire n251641;
   wire n251642;
   wire n251643;
   wire n251644;
   wire n251645;
   wire n251646;
   wire n251647;
   wire n251649;
   wire n251650;
   wire n251651;
   wire n251652;
   wire n251653;
   wire n251654;
   wire n251655;
   wire n251656;
   wire n251657;
   wire n251658;
   wire n251659;
   wire n251660;
   wire n251661;
   wire n251662;
   wire n251663;
   wire n251664;
   wire n251665;
   wire n251666;
   wire n251667;
   wire n251668;
   wire n251669;
   wire n251670;
   wire n251671;
   wire n251672;
   wire n251673;
   wire n251674;
   wire n251675;
   wire n251676;
   wire n251677;
   wire n251678;
   wire n251679;
   wire n251680;
   wire n251681;
   wire n251682;
   wire n251684;
   wire n251685;
   wire n251686;
   wire n251687;
   wire n251688;
   wire n251689;
   wire n251690;
   wire n251691;
   wire n251692;
   wire n251693;
   wire n251694;
   wire n251695;
   wire n251696;
   wire n251697;
   wire n251698;
   wire n251699;
   wire n251700;
   wire n251701;
   wire n251702;
   wire n251703;
   wire n251704;
   wire n251705;
   wire n251706;
   wire n251707;
   wire n251708;
   wire n251709;
   wire n251710;
   wire n251711;
   wire n251712;
   wire n251713;
   wire n251714;
   wire n251715;
   wire n251716;
   wire n251717;
   wire n251719;
   wire n251720;
   wire n251721;
   wire n251722;
   wire n251723;
   wire n251724;
   wire n251726;
   wire n251727;
   wire n251728;
   wire n251729;
   wire n251730;
   wire n251731;
   wire n251732;
   wire n251733;
   wire n251734;
   wire n251735;
   wire n251736;
   wire n251737;
   wire n251738;
   wire n251739;
   wire n251740;
   wire n251741;
   wire n251742;
   wire n251743;
   wire n251744;
   wire n251745;
   wire n251746;
   wire n251747;
   wire n251748;
   wire n251749;
   wire n251750;
   wire n251751;
   wire n251752;
   wire n251753;
   wire n251755;
   wire n251756;
   wire n251757;
   wire n251758;
   wire n251759;
   wire n251760;
   wire n251761;
   wire n251762;
   wire n251763;
   wire n251764;
   wire n251765;
   wire n251766;
   wire n251767;
   wire n251768;
   wire n251769;
   wire n251770;
   wire n251771;
   wire n251772;
   wire n251773;
   wire n251774;
   wire n251775;
   wire n251776;
   wire n251777;
   wire n251778;
   wire n251779;
   wire n251780;
   wire n251781;
   wire n251782;
   wire n251783;
   wire n251784;
   wire n251785;
   wire n251786;
   wire n251787;
   wire n251788;
   wire n251790;
   wire n251791;
   wire n251792;
   wire n251793;
   wire n251794;
   wire n251795;
   wire n251796;
   wire n251797;
   wire n251798;
   wire n251799;
   wire n251800;
   wire n251801;
   wire n251802;
   wire n251803;
   wire n251804;
   wire n251805;
   wire n251806;
   wire n251807;
   wire n251808;
   wire n251809;
   wire n251810;
   wire n251811;
   wire n251812;
   wire n251813;
   wire n251814;
   wire n251815;
   wire n251816;
   wire n251817;
   wire n251818;
   wire n251819;
   wire n251820;
   wire n251821;
   wire n251822;
   wire n251823;
   wire n251825;
   wire n251826;
   wire n251827;
   wire n251828;
   wire n251829;
   wire n251830;
   wire n251832;
   wire n251833;
   wire n251834;
   wire n251835;
   wire n251836;
   wire n251837;
   wire n251838;
   wire n251839;
   wire n251840;
   wire n251841;
   wire n251842;
   wire n251843;
   wire n251844;
   wire n251845;
   wire n251846;
   wire n251847;
   wire n251848;
   wire n251849;
   wire n251850;
   wire n251851;
   wire n251852;
   wire n251853;
   wire n251854;
   wire n251855;
   wire n251856;
   wire n251857;
   wire n251858;
   wire n251859;
   wire n251861;
   wire n251862;
   wire n251863;
   wire n251864;
   wire n251865;
   wire n251866;
   wire n251867;
   wire n251868;
   wire n251869;
   wire n251870;
   wire n251871;
   wire n251872;
   wire n251873;
   wire n251874;
   wire n251875;
   wire n251876;
   wire n251877;
   wire n251878;
   wire n251879;
   wire n251880;
   wire n251881;
   wire n251882;
   wire n251883;
   wire n251884;
   wire n251885;
   wire n251886;
   wire n251887;
   wire n251888;
   wire n251889;
   wire n251890;
   wire n251891;
   wire n251892;
   wire n251893;
   wire n251894;
   wire n251896;
   wire n251897;
   wire n251898;
   wire n251899;
   wire n251900;
   wire n251901;
   wire n251902;
   wire n251903;
   wire n251904;
   wire n251905;
   wire n251906;
   wire n251907;
   wire n251908;
   wire n251909;
   wire n251910;
   wire n251911;
   wire n251912;
   wire n251913;
   wire n251914;
   wire n251915;
   wire n251916;
   wire n251917;
   wire n251918;
   wire n251919;
   wire n251920;
   wire n251921;
   wire n251922;
   wire n251923;
   wire n251924;
   wire n251925;
   wire n251926;
   wire n251927;
   wire n251928;
   wire n251929;
   wire n251930;
   wire n251932;
   wire n251933;
   wire n251934;
   wire n251935;
   wire n251936;
   wire n251937;
   wire n251939;
   wire n251940;
   wire n251941;
   wire n251942;
   wire n251943;
   wire n251944;
   wire n251945;
   wire n251946;
   wire n251947;
   wire n251948;
   wire n251949;
   wire n251950;
   wire n251951;
   wire n251952;
   wire n251953;
   wire n251954;
   wire n251955;
   wire n251956;
   wire n251957;
   wire n251958;
   wire n251959;
   wire n251960;
   wire n251961;
   wire n251962;
   wire n251963;
   wire n251964;
   wire n251965;
   wire n251966;
   wire n251967;
   wire n251969;
   wire n251970;
   wire n251971;
   wire n251972;
   wire n251973;
   wire n251974;
   wire n251975;
   wire n251976;
   wire n251977;
   wire n251978;
   wire n251979;
   wire n251980;
   wire n251981;
   wire n251982;
   wire n251983;
   wire n251984;
   wire n251985;
   wire n251986;
   wire n251987;
   wire n251988;
   wire n251989;
   wire n251990;
   wire n251991;
   wire n251992;
   wire n251993;
   wire n251994;
   wire n251995;
   wire n251996;
   wire n251997;
   wire n251998;
   wire n251999;
   wire n252000;
   wire n252001;
   wire n252002;
   wire n252003;
   wire n252005;
   wire n252006;
   wire n252007;
   wire n252008;
   wire n252009;
   wire n252010;
   wire n252011;
   wire n252012;
   wire n252013;
   wire n252014;
   wire n252015;
   wire n252016;
   wire n252017;
   wire n252018;
   wire n252019;
   wire n252020;
   wire n252021;
   wire n252022;
   wire n252023;
   wire n252024;
   wire n252025;
   wire n252026;
   wire n252027;
   wire n252028;
   wire n252029;
   wire n252030;
   wire n252031;
   wire n252032;
   wire n252033;
   wire n252034;
   wire n252035;
   wire n252036;
   wire n252037;
   wire n252038;
   wire n252039;
   wire n252041;
   wire n252042;
   wire n252043;
   wire n252044;
   wire n252045;
   wire n252046;
   wire n252048;
   wire n252049;
   wire n252050;
   wire n252051;
   wire n252052;
   wire n252053;
   wire n252054;
   wire n252055;
   wire n252056;
   wire n252057;
   wire n252058;
   wire n252059;
   wire n252060;
   wire n252061;
   wire n252062;
   wire n252063;
   wire n252064;
   wire n252065;
   wire n252066;
   wire n252067;
   wire n252068;
   wire n252069;
   wire n252070;
   wire n252071;
   wire n252072;
   wire n252073;
   wire n252074;
   wire n252075;
   wire n252076;
   wire n252078;
   wire n252079;
   wire n252080;
   wire n252081;
   wire n252082;
   wire n252083;
   wire n252084;
   wire n252085;
   wire n252086;
   wire n252087;
   wire n252088;
   wire n252089;
   wire n252090;
   wire n252091;
   wire n252092;
   wire n252093;
   wire n252094;
   wire n252095;
   wire n252096;
   wire n252097;
   wire n252098;
   wire n252099;
   wire n252100;
   wire n252101;
   wire n252102;
   wire n252103;
   wire n252104;
   wire n252105;
   wire n252106;
   wire n252107;
   wire n252108;
   wire n252109;
   wire n252110;
   wire n252111;
   wire n252112;
   wire n252114;
   wire n252115;
   wire n252116;
   wire n252117;
   wire n252118;
   wire n252119;
   wire n252120;
   wire n252121;
   wire n252122;
   wire n252123;
   wire n252124;
   wire n252125;
   wire n252126;
   wire n252127;
   wire n252128;
   wire n252129;
   wire n252130;
   wire n252131;
   wire n252132;
   wire n252133;
   wire n252134;
   wire n252135;
   wire n252136;
   wire n252137;
   wire n252138;
   wire n252139;
   wire n252140;
   wire n252141;
   wire n252142;
   wire n252143;
   wire n252144;
   wire n252145;
   wire n252146;
   wire n252147;
   wire n252148;
   wire n252150;
   wire n252151;
   wire n252152;
   wire n252153;
   wire n252154;
   wire n252155;
   wire n252157;
   wire n252158;
   wire n252159;
   wire n252160;
   wire n252161;
   wire n252162;
   wire n252163;
   wire n252164;
   wire n252165;
   wire n252166;
   wire n252167;
   wire n252168;
   wire n252169;
   wire n252170;
   wire n252171;
   wire n252172;
   wire n252173;
   wire n252174;
   wire n252175;
   wire n252176;
   wire n252177;
   wire n252178;
   wire n252179;
   wire n252180;
   wire n252181;
   wire n252182;
   wire n252183;
   wire n252184;
   wire n252185;
   wire n252187;
   wire n252188;
   wire n252189;
   wire n252190;
   wire n252191;
   wire n252192;
   wire n252193;
   wire n252194;
   wire n252195;
   wire n252196;
   wire n252197;
   wire n252198;
   wire n252199;
   wire n252200;
   wire n252201;
   wire n252202;
   wire n252203;
   wire n252204;
   wire n252205;
   wire n252206;
   wire n252207;
   wire n252208;
   wire n252209;
   wire n252210;
   wire n252211;
   wire n252212;
   wire n252213;
   wire n252214;
   wire n252215;
   wire n252216;
   wire n252217;
   wire n252218;
   wire n252219;
   wire n252220;
   wire n252221;
   wire n252222;
   wire n252224;
   wire n252225;
   wire n252226;
   wire n252227;
   wire n252228;
   wire n252229;
   wire n252230;
   wire n252231;
   wire n252232;
   wire n252233;
   wire n252234;
   wire n252235;
   wire n252236;
   wire n252238;
   wire n252239;
   wire n252240;
   wire n252241;
   wire n252242;
   wire n252243;
   wire n252244;
   wire n252245;
   wire n252246;
   wire n252247;
   wire n252248;
   wire n252249;
   wire n252250;
   wire n252251;
   wire n252252;
   wire n252253;
   wire n252254;
   wire n252255;
   wire n252256;
   wire n252257;
   wire n252258;
   wire n252259;
   wire n252260;
   wire n252261;
   wire n252262;
   wire n252263;
   wire n252264;
   wire n252265;
   wire n252266;
   wire n252267;
   wire n252268;
   wire n252269;
   wire n252270;
   wire n252271;
   wire n252272;
   wire n252273;
   wire n252274;
   wire n252275;
   wire n252276;
   wire n252277;
   wire n252278;
   wire n252279;
   wire n252280;
   wire n252281;
   wire n252282;
   wire n252283;
   wire n252284;
   wire n252285;
   wire n252286;
   wire n252287;
   wire n252288;
   wire n252289;
   wire n252290;
   wire n252291;
   wire n252292;
   wire n252293;
   wire n252294;
   wire n252295;
   wire n252296;
   wire n252297;
   wire n252298;
   wire n252299;
   wire n252300;
   wire n252301;
   wire n252302;
   wire n252303;
   wire n252304;
   wire n252305;
   wire n252306;
   wire n252307;
   wire n252308;
   wire n252309;
   wire n252310;
   wire n252311;
   wire n252312;
   wire n252313;
   wire n252314;
   wire n252315;
   wire n252316;
   wire n252317;
   wire n252318;
   wire n252319;
   wire n252320;
   wire n252321;
   wire n252322;
   wire n252323;
   wire n252324;
   wire n252325;
   wire n252326;
   wire n252327;
   wire n252328;
   wire n252329;
   wire n252330;
   wire n252331;
   wire n252332;
   wire n252333;
   wire n252334;
   wire n252335;
   wire n252336;
   wire n252337;
   wire n252338;
   wire n252339;
   wire n252340;
   wire n252341;
   wire n252342;
   wire n252343;
   wire n252344;
   wire n252345;
   wire n252346;
   wire n252347;
   wire n252348;
   wire n252349;
   wire n252350;
   wire n252351;
   wire n252352;
   wire n252353;
   wire n252354;
   wire n252355;
   wire n252356;
   wire n252357;
   wire n252358;
   wire n252359;
   wire n252360;
   wire n252361;
   wire n252362;
   wire n252363;
   wire n252364;
   wire n252365;
   wire n252366;
   wire n252367;
   wire n252368;
   wire n252369;
   wire n252370;
   wire n252371;
   wire n252372;
   wire n252373;
   wire n252374;
   wire n252375;
   wire n252376;
   wire n252377;
   wire n252378;
   wire n252379;
   wire n252380;
   wire n252381;
   wire n252382;
   wire n252383;
   wire n252384;
   wire n252385;
   wire n252386;
   wire n252387;
   wire n252388;
   wire n252389;
   wire n252390;
   wire n252391;
   wire n252392;
   wire n252393;
   wire n252394;
   wire n252395;
   wire n252396;
   wire n252397;
   wire n252398;
   wire n252399;
   wire n252400;
   wire n252401;
   wire n252402;
   wire n252403;
   wire n252404;
   wire n252405;
   wire n252406;
   wire n252407;
   wire n252408;
   wire n252409;
   wire n252410;
   wire n252411;
   wire n252412;
   wire n252413;
   wire n252414;
   wire n252415;
   wire n252416;
   wire n252417;
   wire n252418;
   wire n252419;
   wire n252420;
   wire n252421;
   wire n252422;
   wire n252423;
   wire n252424;
   wire n252425;
   wire n252426;
   wire n252427;
   wire n252428;
   wire n252429;
   wire n252430;
   wire n252431;
   wire n252432;
   wire n252433;
   wire n252434;
   wire n252435;
   wire n252436;
   wire n252437;
   wire n252438;
   wire n252439;
   wire n252440;
   wire n252441;
   wire n252442;
   wire n252443;
   wire n252444;
   wire n252445;
   wire n252446;
   wire n252447;
   wire n252448;
   wire n252449;
   wire n252450;
   wire n252451;
   wire n252452;
   wire n252453;
   wire n252454;
   wire n252455;
   wire n252456;
   wire n252457;
   wire n252458;
   wire n252459;
   wire n252460;
   wire n252461;
   wire n252462;
   wire n252463;
   wire n252464;
   wire n252465;
   wire n252466;
   wire n252467;
   wire n252468;
   wire n252469;
   wire n252470;
   wire n252471;
   wire n252472;
   wire n252473;
   wire n252474;
   wire n252475;
   wire n252476;
   wire n252477;
   wire n252478;
   wire n252479;
   wire n252480;
   wire n252481;
   wire n252482;
   wire n252483;
   wire n252484;
   wire n252485;
   wire n252486;
   wire n252487;
   wire n252488;
   wire n252489;
   wire n252490;
   wire n252491;
   wire n252492;
   wire n252493;
   wire n252494;
   wire n252495;
   wire n252496;
   wire n252497;
   wire n252498;
   wire n252499;
   wire n252500;
   wire n252501;
   wire n252502;
   wire n252503;
   wire n252504;
   wire n252505;
   wire n252506;
   wire n252507;
   wire n252508;
   wire n252509;
   wire n252510;
   wire n252511;
   wire n252512;
   wire n252513;
   wire n252514;
   wire n252515;
   wire n252516;
   wire n252517;
   wire n252518;
   wire n252519;
   wire n252520;
   wire n252521;
   wire n252522;
   wire n252523;
   wire n252524;
   wire n252525;
   wire n252526;
   wire n252527;
   wire n252528;
   wire n252529;
   wire n252530;
   wire n252531;
   wire n252532;
   wire n252533;
   wire n252534;
   wire n252535;
   wire n252536;
   wire n252537;
   wire n252538;
   wire n252540;
   wire n252541;
   wire n252542;
   wire n252543;
   wire n252544;
   wire n252545;
   wire n252546;
   wire n252547;
   wire n252548;
   wire n252549;
   wire n252550;
   wire n252551;
   wire n252552;
   wire n252553;
   wire n252554;
   wire n252555;
   wire n252556;
   wire n252557;
   wire n252558;
   wire n252559;
   wire n252560;
   wire n252561;
   wire n252562;
   wire n252563;
   wire n252564;
   wire n252565;
   wire n252566;
   wire n252567;
   wire n252568;
   wire n252569;
   wire n252570;
   wire n252571;
   wire n252572;
   wire n252573;
   wire n252574;
   wire n252575;
   wire n252576;
   wire n252577;
   wire n252578;
   wire n252579;
   wire n252580;
   wire n252581;
   wire n252582;
   wire n252583;
   wire n252584;
   wire n252585;
   wire n252586;
   wire n252587;
   wire n252588;
   wire n252589;
   wire n252590;
   wire n252591;
   wire n252592;
   wire n252593;
   wire n252594;
   wire n252595;
   wire n252596;
   wire n252597;
   wire n252598;
   wire n252599;
   wire n252600;
   wire n252601;
   wire n252602;
   wire n252603;
   wire n252604;
   wire n252605;
   wire n252606;
   wire n252607;
   wire n252608;
   wire n252609;
   wire n252610;
   wire n252611;
   wire n252612;
   wire n252613;
   wire n252614;
   wire n252615;
   wire n252616;
   wire n252617;
   wire n252618;
   wire n252619;
   wire n252620;
   wire n252621;
   wire n252622;
   wire n252623;
   wire n252624;
   wire n252625;
   wire n252626;
   wire n252627;
   wire n252628;
   wire n252629;
   wire n252630;
   wire n252631;
   wire n252632;
   wire n252633;
   wire n252634;
   wire n252635;
   wire n252636;
   wire n252637;
   wire n252638;
   wire n252639;
   wire n252640;
   wire n252641;
   wire n252642;
   wire n252643;
   wire n252644;
   wire n252645;
   wire n252646;
   wire n252647;
   wire n252648;
   wire n252649;
   wire n252650;
   wire n252651;
   wire n252652;
   wire n252653;
   wire n252654;
   wire n252655;
   wire n252656;
   wire n252657;
   wire n252658;
   wire n252659;
   wire n252660;
   wire n252661;
   wire n252662;
   wire n252663;
   wire n252664;
   wire n252665;
   wire n252666;
   wire n252667;
   wire n252668;
   wire n252669;
   wire n252670;
   wire n252671;
   wire n252672;
   wire n252673;
   wire n252674;
   wire n252675;
   wire n252676;
   wire n252677;
   wire n252678;
   wire n252679;
   wire n252680;
   wire n252681;
   wire n252682;
   wire n252683;
   wire n252684;
   wire n252685;
   wire n252686;
   wire n252687;
   wire n252688;
   wire n252689;
   wire n252690;
   wire n252691;
   wire n252692;
   wire n252693;
   wire n252694;
   wire n252695;
   wire n252696;
   wire n252697;
   wire n252698;
   wire n252699;
   wire n252700;
   wire n252701;
   wire n252702;
   wire n252703;
   wire n252704;
   wire n252705;
   wire n252706;
   wire n252707;
   wire n252708;
   wire n252709;
   wire n252710;
   wire n252711;
   wire n252712;
   wire n252713;
   wire n252714;
   wire n252715;
   wire n252716;
   wire n252717;
   wire n252718;
   wire n252719;
   wire n252720;
   wire n252721;
   wire n252722;
   wire n252723;
   wire n252724;
   wire n252725;
   wire n252726;
   wire n252727;
   wire n252728;
   wire n252729;
   wire n252730;
   wire n252731;
   wire n252732;
   wire n252733;
   wire n252734;
   wire n252735;
   wire n252736;
   wire n252737;
   wire n252738;
   wire n252739;
   wire n252740;
   wire n252741;
   wire n252742;
   wire n252743;
   wire n252744;
   wire n252745;
   wire n252746;
   wire n252747;
   wire n252748;
   wire n252749;
   wire n252750;
   wire n252751;
   wire n252752;
   wire n252753;
   wire n252754;
   wire n252755;
   wire n252756;
   wire n252757;
   wire n252758;
   wire n252759;
   wire n252760;
   wire n252761;
   wire n252762;
   wire n252763;
   wire n252764;
   wire n252765;
   wire n252766;
   wire n252767;
   wire n252768;
   wire n252769;
   wire n252770;
   wire n252771;
   wire n252772;
   wire n252773;
   wire n252774;
   wire n252775;
   wire n252776;
   wire n252777;
   wire n252778;
   wire n252779;
   wire n252780;
   wire n252781;
   wire n252782;
   wire n252783;
   wire n252784;
   wire n252785;
   wire n252786;
   wire n252787;
   wire n252788;
   wire n252789;
   wire n252790;
   wire n252791;
   wire n252792;
   wire n252793;
   wire n252794;
   wire n252795;
   wire n252796;
   wire n252797;
   wire n252798;
   wire n252799;
   wire n252800;
   wire n252801;
   wire n252802;
   wire n252803;
   wire n252804;
   wire n252805;
   wire n252806;
   wire n252807;
   wire n252808;
   wire n252809;
   wire n252810;
   wire n252811;
   wire n252812;
   wire n252813;
   wire n252814;
   wire n252815;
   wire n252816;
   wire n252817;
   wire n252818;
   wire n252819;
   wire n252820;
   wire n252821;
   wire n252822;
   wire n252823;
   wire n252824;
   wire n252825;
   wire n252826;
   wire n252827;
   wire n252828;
   wire n252829;
   wire n252831;
   wire n252832;
   wire n252834;
   wire n252835;
   wire n252836;
   wire n252837;
   wire n252838;
   wire n252839;
   wire n252840;
   wire n252841;
   wire n252842;
   wire n252843;
   wire n252844;
   wire n252845;
   wire n252846;
   wire n252847;
   wire n252848;
   wire n252849;
   wire n252850;
   wire n252851;
   wire n252852;
   wire n252853;
   wire n252854;
   wire n252855;
   wire n252856;
   wire n252857;
   wire n252858;
   wire n252859;
   wire n252860;
   wire n252861;
   wire n252862;
   wire n252863;
   wire n252865;
   wire n252866;
   wire n252867;
   wire n252868;
   wire n252869;
   wire n252871;
   wire n252872;
   wire n252873;
   wire n252874;
   wire n252875;
   wire n252876;
   wire n252877;
   wire n252878;
   wire n252879;
   wire n252880;
   wire n252881;
   wire n252882;
   wire n252883;
   wire n252884;
   wire n252885;
   wire n252886;
   wire n252887;
   wire n252888;
   wire n252889;
   wire n252890;
   wire n252891;
   wire n252892;
   wire n252893;
   wire n252894;
   wire n252895;
   wire n252896;
   wire n252897;
   wire n252898;
   wire n252899;
   wire n252900;
   wire n252901;
   wire n252902;
   wire n252903;
   wire n252904;
   wire n252905;
   wire n252906;
   wire n252907;
   wire n252908;
   wire n252909;
   wire n252911;
   wire n252912;
   wire n252913;
   wire n252914;
   wire n252915;
   wire n252916;
   wire n252917;
   wire n252918;
   wire n252919;
   wire n252920;
   wire n252921;
   wire n252922;
   wire n252923;
   wire n252924;
   wire n252925;
   wire n252926;
   wire n252927;
   wire n252928;
   wire n252929;
   wire n252930;
   wire n252931;
   wire n252932;
   wire n252933;
   wire n252934;
   wire n252935;
   wire n252936;
   wire n252937;
   wire n252938;
   wire n252939;
   wire n252940;
   wire n252941;
   wire n252942;
   wire n252943;
   wire n252944;
   wire n252945;
   wire n252946;
   wire n252947;
   wire n252948;
   wire n252949;
   wire n252950;
   wire n252951;
   wire n252952;
   wire n252953;
   wire n252954;
   wire n252955;
   wire n252956;
   wire n252957;
   wire n252958;
   wire n252960;
   wire n252961;
   wire n252962;
   wire n252963;
   wire n252964;
   wire n252965;
   wire n252966;
   wire n252967;
   wire n252968;
   wire n252969;
   wire n252970;
   wire n252971;
   wire n252972;
   wire n252973;
   wire n252974;
   wire n252975;
   wire n252976;
   wire n252977;
   wire n252978;
   wire n252979;
   wire n252980;
   wire n252981;
   wire n252982;
   wire n252983;
   wire n252984;
   wire n252985;
   wire n252986;
   wire n252987;
   wire n252988;
   wire n252989;
   wire n252990;
   wire n252991;
   wire n252992;
   wire n252993;
   wire n252994;
   wire n252995;
   wire n252996;
   wire n252997;
   wire n252998;
   wire n252999;
   wire n253000;
   wire n253001;
   wire n253002;
   wire n253003;
   wire n253004;
   wire n253005;
   wire n253006;
   wire n253007;
   wire n253008;
   wire n253009;
   wire n253010;
   wire n253011;
   wire n253012;
   wire n253013;
   wire n253014;
   wire n253015;
   wire n253016;
   wire n253017;
   wire n253018;
   wire n253019;
   wire n253020;
   wire n253021;
   wire n253022;
   wire n253023;
   wire n253024;
   wire n253025;
   wire n253026;
   wire n253027;
   wire n253028;
   wire n253029;
   wire n253030;
   wire n253037;
   wire n253038;
   wire n253039;
   wire n253040;
   wire n253041;
   wire n253042;
   wire n253043;
   wire n253044;
   wire n253045;
   wire n253046;
   wire n253047;
   wire n253048;
   wire n253049;
   wire n253050;
   wire n253051;
   wire n253052;
   wire n253053;
   wire n253054;
   wire n253055;
   wire n253056;
   wire n253057;
   wire n253058;
   wire n253059;
   wire n253060;
   wire n253061;
   wire n253062;
   wire n253063;
   wire n253064;
   wire n253065;
   wire n253066;
   wire n253067;
   wire n253068;
   wire n253069;
   wire n253070;
   wire n253071;
   wire n253072;
   wire n253073;
   wire n253074;
   wire n253075;
   wire n253076;
   wire n253077;
   wire n253078;
   wire n253079;
   wire n253080;
   wire n253081;
   wire n253082;
   wire n253083;
   wire n253084;
   wire n253085;
   wire n253086;
   wire n253087;
   wire n253088;
   wire n253089;
   wire n253090;
   wire n253091;
   wire n253092;
   wire n253093;
   wire n253094;
   wire n253095;
   wire n253096;
   wire n253097;
   wire n253098;
   wire n253099;
   wire n253100;
   wire n253101;
   wire n253102;
   wire n253103;
   wire n253104;
   wire n253105;
   wire n253106;
   wire n253107;
   wire n253108;
   wire n253109;
   wire n253110;
   wire n253111;
   wire n253112;
   wire n253113;
   wire n253114;
   wire n253115;
   wire n253116;
   wire n253117;
   wire n253118;
   wire n253119;
   wire n253120;
   wire n253121;
   wire n253122;
   wire n253123;
   wire n253124;
   wire n253125;
   wire [11:0] g_mbc_r;
   wire [11:0] g_pcut_r;
   wire [6:0] g_hs60p_r;
   wire [6:0] g_vs60p_r;
   wire [17:0] g_fcyc_r;
   wire [4:1] v_paramadr_r;
   wire [24:0] v_paramdata_r;
   wire [6:0] g_hsdc_r;
   wire [6:0] g_vsdc_r;
   wire [4:0] v_vldstatus_r;
   wire [1:0] g_vldmode_r;
   wire [31:0] y1_bs_data_r;
   wire [31:10] g_field_start_add_r;
   wire [11:0] g_field_offset_r;
   wire [11:0] g_cbcr_offset_r;
   wire [31:0] vh_1_ph_add;
   wire [4:1] vldtop_vld_syndec_ADP;
   wire [31:0] vldtop_vld_syndec_UREG;
   wire [4:1] vldtop_vld_syndec_vld_seqhed_pre_SHIFT;
   wire [1:0] vldtop_vld_syndec_vld_vscdet_v_prezerohld_r;
   wire [1:0] vldtop_vld_syndec_vld_vscdet_v_prezerotmp_r;
   wire [1:0] vldtop_vld_syndec_vld_vscdet_v_detvald_r;
   wire [31:0] vldtop_vld_syndec_vld_vlfeed_temporal;
   wire [31:0] vldtop_vld_syndec_vld_vlfeed_lower;
   wire [1:0] busrtop_b_rreq_vrh_cnt_16byte_r;
   wire [1:0] busrtop_b_rreq_vrh_cnt_18byte_r;
   wire [9:0] busrtop_b_rreq_vrh_add1_r;
   wire [31:13] busrtop_b_rreq_vrh_rrq_fldstatadd_r;
   wire [31:0] regtop_g_mem_rd2_r;
   wire [31:0] regtop_v1_hdi00_d;
   wire [5:0] regtop_v1_hdi00_a;
   wire [31:8] regtop_g_atscd_r;
   wire [31:8] regtop_g_usrd_r;
   wire [6:0] regtop_g_adb_cpu_r;
   wire [6:0] regtop_g_adb_r;
   wire [6:0] regtop_g_udb_cpu_r;
   wire [6:0] regtop_g_udb2_r;
   wire [6:0] regtop_g_udb1_r;
   wire [6:0] regtop_g_udb0_r;
   wire [15:0] regtop_g_fcvo2_r;
   wire [15:0] regtop_g_fcho2_r;
   wire [15:0] regtop_g_fcvo1_r;
   wire [15:0] regtop_g_fcho1_r;
   wire [15:0] regtop_g_fcvo0_r;
   wire [15:0] regtop_g_fcho0_r;
   wire [1:0] regtop_g_nfco_r;
   wire [7:0] regtop_g_scp_r;
   wire [6:0] regtop_g_ba_r;
   wire [2:0] regtop_g_fs_r;
   wire [1:0] regtop_g_pis_r;
   wire [15:0] regtop_g_vd_r;
   wire [2:0] regtop_g_pct_r;
   wire [9:0] regtop_g_tr_r;
   wire [23:0] regtop_g_tmc_r;
   wire [13:0] regtop_g_dvs_r;
   wire [13:0] regtop_g_dhs_r;
   wire [7:0] regtop_g_mc_r;
   wire [7:0] regtop_g_tc_r;
   wire [7:0] regtop_g_cp_r;
   wire [2:0] regtop_g_vf_r;
   wire [1:0] regtop_g_cf_r;
   wire [7:0] regtop_g_pali_r;
   wire [9:0] regtop_g_vbsv_r;
   wire [17:0] regtop_g_brv_r;
   wire [3:0] regtop_g_frc_r;
   wire [3:0] regtop_g_ari_r;
   wire [11:0] regtop_g_vsv_r;
   wire [11:0] regtop_g_hsv_r;
   wire [6:0] regtop_g_embv_adr_r;
   wire [6:0] regtop_g_embh_adr_r;
   wire [22:0] regtop_g_nfst_r;
   wire [9:0] regtop_g_fbst_r;
   wire [5:0] regtop_g_fpst_r;
   wire [2:0] regtop_g_init_cnt_r;
   wire [31:0] regtop_w1_hdi00_q;
   wire [3:0] regtop_g_dspfld_num2_r;
   wire [3:0] regtop_g_dspfld_num1_r;
   wire [4:0] regtop_g_vldstatus_r;
   wire [24:0] regtop_g_paramdata_r;
   wire [7:0] regtop_g_paramadr_r;
   wire [31:0] regtop_g_mem_rd_r;
   wire [31:0] regtop_g_wd_r;
   wire [8:2] regtop_g_a_r;
   wire [2047:0] regtop_dchdi_w1_hdi00;

   assign v1_dspfld_num1[3] = 1'b1 ;
   assign v1_dspfld_num1[2] = 1'b1 ;
   assign v1_dspfld_num1[1] = 1'b1 ;
   assign v1_dspfld_num1[0] = 1'b1 ;
   assign v1_dspfld_sc1 = 1'b0 ;
   assign v1_dspfld_num2[3] = 1'b1 ;
   assign v1_dspfld_num2[2] = 1'b1 ;
   assign v1_dspfld_num2[1] = 1'b1 ;
   assign v1_dspfld_num2[0] = 1'b1 ;
   assign v1_dspfld_sc2 = 1'b0 ;
   assign v1_dsp_ps = 1'b0 ;
   assign vmem_data_out[31] = 1'b0 ;
   assign vmem_data_out[30] = 1'b0 ;
   assign vmem_data_out[29] = 1'b0 ;
   assign vmem_data_out[28] = 1'b0 ;
   assign vmem_data_out[27] = 1'b0 ;
   assign vmem_data_out[26] = 1'b0 ;
   assign v1_sd_pichead_s = 1'b0 ;
   assign vmem_we_n[0] = vmem_we_n[1] ;
   assign vmem_we_n[2] = vmem_we_n[1] ;
   assign vmem_we_n[3] = vmem_we_n[1] ;

   na03f06 FE_RC_50_0 (.o(n245592),
	.a(n245591),
	.b(n245590),
	.c(n245589));
   ao22s02 FE_RC_49_0 (.o(n245485),
	.a(n245478),
	.b(FE_OFN4_n245443),
	.c(n249786),
	.d(g_vsdc_r[0]));
   na04f01 FE_RC_48_0 (.o(n245533),
	.a(n252564),
	.b(n252314),
	.c(n245569),
	.d(n245762));
   ao12f04 FE_RC_47_0 (.o(n245664),
	.a(n245331),
	.b(n245332),
	.c(n245734));
   oa12f02 FE_RC_46_0 (.o(n249213),
	.a(n249212),
	.b(n249242),
	.c(n252648));
   ao12f02 FE_RC_45_0 (.o(n246205),
	.a(n246203),
	.b(n246204),
	.c(FE_OFN4_n245443));
   na04f01 FE_RC_44_0 (.o(n248463),
	.a(n248455),
	.b(n248457),
	.c(n248456),
	.d(n248454));
   na04f02 FE_RC_43_0 (.o(n249819),
	.a(n249818),
	.b(n249815),
	.c(n249816),
	.d(n249817));
   ao12f04 FE_RC_42_0 (.o(n245697),
	.a(n245375),
	.b(n245675),
	.c(n245376));
   oa12f06 FE_RC_41_0 (.o(n245659),
	.a(n245695),
	.b(n245697),
	.c(n245694));
   ao22f04 FE_RC_40_0 (.o(n248991),
	.a(n249066),
	.b(n248984),
	.c(n249041),
	.d(regtop_g_adb_r[2]));
   ao12f06 FE_RC_39_0 (.o(n245652),
	.a(n245388),
	.b(n245659),
	.c(n245658));
   ao12f04 FE_RC_38_0 (.o(n245607),
	.a(n245424),
	.b(n245614),
	.c(n245613));
   oa12f02 FE_RC_37_0 (.o(n244990),
	.a(n249035),
	.b(n249077),
	.c(FE_OFN507_regtop_g_a_r_4_));
   oa12f06 FE_RC_36_0 (.o(n245644),
	.a(n245650),
	.b(n245652),
	.c(n245649));
   ao12f08 FE_RC_35_0 (.o(n245622),
	.a(n245412),
	.b(n245629),
	.c(n245628));
   oa12f08 FE_RC_34_0 (.o(n245614),
	.a(n245620),
	.b(n245622),
	.c(n245619));
   ao12f08 FE_RC_33_0 (.o(n245637),
	.a(n245400),
	.b(n245644),
	.c(n245643));
   no04f02 FE_RC_32_0 (.o(n248270),
	.a(n248247),
	.b(n248248),
	.c(n248246),
	.d(FE_OFN236_n248245));
   in01f04 FE_OCPC583_n247126 (.o(FE_OCPN583_n247126),
	.a(FE_OCPN582_n247126));
   in01f01 FE_OCPC582_n247126 (.o(FE_OCPN582_n247126),
	.a(n247126));
   no03f06 FE_RC_31_0 (.o(n246184),
	.a(n246181),
	.b(n246182),
	.c(n246183));
   oa12f04 FE_RC_29_0 (.o(n246109),
	.a(n246174),
	.b(n246173),
	.c(n246178));
   oa12f04 FE_RC_28_0 (.o(n245675),
	.a(n245355),
	.b(n245664),
	.c(n245356));
   oa12f02 FE_RC_26_0 (.o(n246108),
	.a(n246106),
	.b(n246152),
	.c(n246107));
   ao22f04 FE_RC_25_0 (.o(n248993),
	.a(n249066),
	.b(n248990),
	.c(n249041),
	.d(regtop_g_adb_r[3]));
   oa12f08 FE_RC_24_0 (.o(n245629),
	.a(n245635),
	.b(n245637),
	.c(n245634));
   ao12f04 FE_RC_23_0 (.o(n246146),
	.a(n246108),
	.b(n246110),
	.c(n246109));
   oa12f02 FE_RC_22_0 (.o(n244987),
	.a(n249075),
	.b(n249077),
	.c(FE_OFN509_regtop_g_a_r_7_));
   in01f02 FE_OFC581_n248442 (.o(FE_OFN581_n248442),
	.a(FE_OFN580_n248442));
   in01f01 FE_OFC580_n248442 (.o(FE_OFN580_n248442),
	.a(n248442));
   in01f02 FE_OFC579_n248820 (.o(FE_OFN579_n248820),
	.a(FE_OFN578_n248820));
   in01f01 FE_OFC578_n248820 (.o(FE_OFN578_n248820),
	.a(n248820));
   in01f08 FE_OFC577_n247126 (.o(FE_OFN577_n247126),
	.a(FE_OFN576_n247126));
   in01f02 FE_OFC576_n247126 (.o(FE_OFN576_n247126),
	.a(n247126));
   in01f02 FE_OFC575_n245444 (.o(FE_OFN575_n245444),
	.a(FE_OFN574_n245444));
   in01f01 FE_OFC574_n245444 (.o(FE_OFN574_n245444),
	.a(n245444));
   in01f01 FE_OFC573_n249242 (.o(FE_OFN573_n249242),
	.a(FE_OFN572_n249242));
   in01f01 FE_OFC572_n249242 (.o(FE_OFN572_n249242),
	.a(n249242));
   in01f01 FE_OFC571_n248074 (.o(FE_OFN571_n248074),
	.a(FE_OFN570_n248074));
   in01f01 FE_OFC570_n248074 (.o(FE_OFN570_n248074),
	.a(n248074));
   in01f02 FE_OFC569_n247780 (.o(FE_OFN569_n247780),
	.a(FE_OFN568_n247780));
   in01f02 FE_OFC568_n247780 (.o(FE_OFN568_n247780),
	.a(n247780));
   in01f02 FE_OFC567_n247541 (.o(FE_OFN567_n247541),
	.a(FE_OFN566_n247541));
   in01f01 FE_OFC566_n247541 (.o(FE_OFN566_n247541),
	.a(n247541));
   in01f02 FE_OFC565_n247738 (.o(FE_OFN565_n247738),
	.a(FE_OFN564_n247738));
   in01f01 FE_OFC564_n247738 (.o(FE_OFN564_n247738),
	.a(n247738));
   in01f04 FE_OFC563_n250717 (.o(FE_OFN563_n250717),
	.a(FE_OFN562_n250717));
   in01f01 FE_OFC562_n250717 (.o(FE_OFN562_n250717),
	.a(FE_OFN292_n250717));
   in01f03 FE_OFC561_n251852 (.o(FE_OFN561_n251852),
	.a(FE_OFN559_n251852));
   in01f01 FE_OFC560_n251852 (.o(FE_OFN560_n251852),
	.a(FE_OFN559_n251852));
   in01f01 FE_OFC559_n251852 (.o(FE_OFN559_n251852),
	.a(FE_OFN335_n251852));
   in01f04 FE_OFC558_n252630 (.o(FE_OFN558_n252630),
	.a(FE_OFN557_n252630));
   in01f01 FE_OFC557_n252630 (.o(FE_OFN557_n252630),
	.a(n252630));
   in01f04 FE_OFC556_n250770 (.o(FE_OFN556_n250770),
	.a(FE_OFN555_n250770));
   in01f02 FE_OFC555_n250770 (.o(FE_OFN555_n250770),
	.a(n250770));
   in01f02 FE_OFC554_n247778 (.o(FE_OFN554_n247778),
	.a(FE_OFN553_n247778));
   in01f01 FE_OFC553_n247778 (.o(FE_OFN553_n247778),
	.a(n247778));
   in01f01 FE_RC_20_0 (.o(n246636),
	.a(FE_RN_9_0));
   ao12f01 FE_RC_19_0 (.o(FE_RN_9_0),
	.a(n246633),
	.b(FE_OFN6_n246618),
	.c(n249079));
   in01f01 FE_RC_18_0 (.o(n245920),
	.a(FE_RN_8_0));
   ao12f01 FE_RC_17_0 (.o(FE_RN_8_0),
	.a(n245918),
	.b(FE_OFN218_n246238),
	.c(n249078));
   in01f01 FE_RC_16_0 (.o(n246632),
	.a(FE_RN_7_0));
   ao12f01 FE_RC_15_0 (.o(FE_RN_7_0),
	.a(n246629),
	.b(FE_OFN6_n246618),
	.c(n249079));
   in01f01 FE_RC_14_0 (.o(n245917),
	.a(FE_RN_6_0));
   ao12f01 FE_RC_13_0 (.o(FE_RN_6_0),
	.a(n245915),
	.b(FE_OFN218_n246238),
	.c(n249078));
   in01f01 FE_RC_12_0 (.o(n246628),
	.a(FE_RN_5_0));
   ao12f01 FE_RC_11_0 (.o(FE_RN_5_0),
	.a(n246625),
	.b(FE_OFN6_n246618),
	.c(n249079));
   in01f01 FE_RC_10_0 (.o(n245914),
	.a(FE_RN_4_0));
   ao12f01 FE_RC_9_0 (.o(FE_RN_4_0),
	.a(n245912),
	.b(FE_OFN218_n246238),
	.c(n249078));
   in01f01 FE_RC_8_0 (.o(n246624),
	.a(FE_RN_3_0));
   ao12f01 FE_RC_7_0 (.o(FE_RN_3_0),
	.a(n246621),
	.b(FE_OFN6_n246618),
	.c(n249079));
   in01f01 FE_RC_6_0 (.o(n245908),
	.a(FE_RN_2_0));
   ao12f01 FE_RC_5_0 (.o(FE_RN_2_0),
	.a(n245906),
	.b(FE_OFN218_n246238),
	.c(n249078));
   in01f01 FE_RC_4_0 (.o(n246620),
	.a(FE_RN_1_0));
   ao12f01 FE_RC_3_0 (.o(FE_RN_1_0),
	.a(n246615),
	.b(FE_OFN6_n246618),
	.c(n249079));
   in01f01 FE_RC_2_0 (.o(n245911),
	.a(FE_RN_0_0));
   ao12f01 FE_RC_1_0 (.o(FE_RN_0_0),
	.a(n245909),
	.b(FE_OFN218_n246238),
	.c(n249078));
   ao12f01 FE_RC_0_0 (.o(n249462),
	.a(n249548),
	.b(n252972),
	.c(g_field_start_add_r[14]));
   in01f04 FE_OFC552_n245462 (.o(FE_OFN552_n245462),
	.a(n245462));
   in01f03 FE_OFC551_n249140 (.o(FE_OFN551_n249140),
	.a(n249140));
   in01f03 FE_OFC550_n249113 (.o(FE_OFN550_n249113),
	.a(n249113));
   in01f01 FE_OFC549_regtop_g_a_r_2_ (.o(FE_OFN549_regtop_g_a_r_2_),
	.a(regtop_g_a_r[2]));
   in01f02 FE_OFC548_regtop_g_a_r_2_ (.o(FE_OFN548_regtop_g_a_r_2_),
	.a(regtop_g_a_r[2]));
   in01f01 FE_OFC547_n245460 (.o(FE_OFN547_n245460),
	.a(n245460));
   in01f02 FE_OFC546_n245460 (.o(FE_OFN546_n245460),
	.a(n245460));
   in01f02 FE_OFC545_n245460 (.o(FE_OFN545_n245460),
	.a(n245460));
   in01f02 FE_OFC544_n252912 (.o(FE_OFN544_n252912),
	.a(n252912));
   in01f01 FE_OFC543_vldtop_vld_syndec_vld_vlfeed_lower_26_ (.o(FE_OFN543_vldtop_vld_syndec_vld_vlfeed_lower_26_),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[26]));
   in01f01 FE_OFC542_n248424 (.o(FE_OFN542_n248424),
	.a(FE_OFN541_n248424));
   in01f02 FE_OFC541_n248424 (.o(FE_OFN541_n248424),
	.a(n248424));
   in01f01 FE_OFC540_vldtop_vld_syndec_vld_vlfeed_lower_12_ (.o(FE_OFN540_vldtop_vld_syndec_vld_vlfeed_lower_12_),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[12]));
   in01f01 FE_OFC537_vldtop_vld_syndec_vld_vlfeed_lower_18_ (.o(FE_OFN537_vldtop_vld_syndec_vld_vlfeed_lower_18_),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[18]));
   in01f02 FE_OFC534_regtop_g_a_r_5_ (.o(FE_OFN534_regtop_g_a_r_5_),
	.a(regtop_g_a_r[5]));
   in01f02 FE_OFC532_regtop_g_a_r_5_ (.o(FE_OFN532_regtop_g_a_r_5_),
	.a(regtop_g_a_r[5]));
   in01f01 FE_OFC530_vldtop_vld_syndec_vld_vlfeed_lower_14_ (.o(FE_OFN530_vldtop_vld_syndec_vld_vlfeed_lower_14_),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[14]));
   in01f06 FE_OFC527_n249828 (.o(FE_OFN527_n249828),
	.a(n249828));
   in01f01 FE_OFC526_n249548 (.o(FE_OFN526_n249548),
	.a(n249548));
   in01f01 FE_OFC525_vldtop_vld_syndec_vld_vlfeed_lower_16_ (.o(FE_OFN525_vldtop_vld_syndec_vld_vlfeed_lower_16_),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[16]));
   in01f02 FE_OFC524_n247696 (.o(FE_OFN524_n247696),
	.a(FE_OFN523_n247696));
   in01f01 FE_OFC523_n247696 (.o(FE_OFN523_n247696),
	.a(n247696));
   in01f02 FE_OFC522_n248508 (.o(FE_OFN522_n248508),
	.a(FE_OFN521_n248508));
   in01f01 FE_OFC521_n248508 (.o(FE_OFN521_n248508),
	.a(n248508));
   in01f04 FE_OFC520_regtop_g_a_r_6_ (.o(FE_OFN520_regtop_g_a_r_6_),
	.a(regtop_g_a_r[6]));
   in01f01 FE_OFC519_regtop_g_a_r_6_ (.o(FE_OFN519_regtop_g_a_r_6_),
	.a(regtop_g_a_r[6]));
   in01f01 FE_OFC517_regtop_g_a_r_6_ (.o(FE_OFN517_regtop_g_a_r_6_),
	.a(regtop_g_a_r[6]));
   in01f02 FE_OFC516_regtop_v1_hdi00_a_0_ (.o(FE_OFN516_regtop_v1_hdi00_a_0_),
	.a(regtop_v1_hdi00_a[0]));
   in01f03 FE_OFC514_n247538 (.o(FE_OFN514_n247538),
	.a(FE_OFN513_n247538));
   in01f01 FE_OFC513_n247538 (.o(FE_OFN513_n247538),
	.a(n247538));
   in01f01 FE_OFC512_n248634 (.o(FE_OFN512_n248634),
	.a(FE_OFN511_n248634));
   in01f01 FE_OFC511_n248634 (.o(FE_OFN511_n248634),
	.a(n248634));
   in01f01 FE_OFC510_regtop_g_a_r_7_ (.o(FE_OFN510_regtop_g_a_r_7_),
	.a(regtop_g_a_r[7]));
   in01f02 FE_OFC509_regtop_g_a_r_7_ (.o(FE_OFN509_regtop_g_a_r_7_),
	.a(regtop_g_a_r[7]));
   in01f04 FE_OFC508_n252540 (.o(FE_OFN508_n252540),
	.a(n252540));
   in01f02 FE_OFC507_regtop_g_a_r_4_ (.o(FE_OFN507_regtop_g_a_r_4_),
	.a(regtop_g_a_r[4]));
   in01f01 FE_OFC506_regtop_g_a_r_4_ (.o(FE_OFN506_regtop_g_a_r_4_),
	.a(regtop_g_a_r[4]));
   in01f01 FE_OFC505_regtop_g_a_r_4_ (.o(FE_OFN505_regtop_g_a_r_4_),
	.a(regtop_g_a_r[4]));
   in01f01 FE_OFC504_regtop_g_a_r_4_ (.o(FE_OFN504_regtop_g_a_r_4_),
	.a(regtop_g_a_r[4]));
   in01f01 FE_OFC503_n246205 (.o(FE_OFN503_n246205),
	.a(FE_OFN502_n246205));
   in01f06 FE_OFC502_n246205 (.o(FE_OFN502_n246205),
	.a(FE_OFN500_n246205));
   in01f02 FE_OFC501_n246205 (.o(FE_OFN501_n246205),
	.a(FE_OFN500_n246205));
   in01f02 FE_OFC500_n246205 (.o(FE_OFN500_n246205),
	.a(n246205));
   in01f01 FE_OFC499_n253015 (.o(FE_OFN499_n253015),
	.a(FE_OFN498_n253015));
   in01f02 FE_OFC498_n253015 (.o(FE_OFN498_n253015),
	.a(n253015));
   in01f02 FE_OFC497_n249947 (.o(FE_OFN497_n249947),
	.a(n249947));
   in01f01 FE_OFC496_n249242 (.o(FE_OFN496_n249242),
	.a(n249242));
   in01f03 FE_OFC494_n252377 (.o(FE_OFN494_n252377),
	.a(n252377));
   in01f01 FE_OFC493_n252377 (.o(FE_OFN493_n252377),
	.a(n252377));
   in01f01 FE_OFC492_n252377 (.o(FE_OFN492_n252377),
	.a(n252377));
   in01f04 FE_OFC491_regtop_g_a_r_3_ (.o(FE_OFN491_regtop_g_a_r_3_),
	.a(regtop_g_a_r[3]));
   in01f01 FE_OFC490_regtop_g_a_r_3_ (.o(FE_OFN490_regtop_g_a_r_3_),
	.a(regtop_g_a_r[3]));
   in01f06 FE_OFC489_n249763 (.o(FE_OFN489_n249763),
	.a(n249763));
   in01f01 FE_OFC488_n245940 (.o(FE_OFN488_n245940),
	.a(FE_OFN485_n245940));
   in01f04 FE_OFC486_n245940 (.o(FE_OFN486_n245940),
	.a(FE_OFN484_n245940));
   in01f01 FE_OFC485_n245940 (.o(FE_OFN485_n245940),
	.a(FE_OFN484_n245940));
   in01f01 FE_OFC484_n245940 (.o(FE_OFN484_n245940),
	.a(n245940));
   in01f02 FE_OFC483_n249211 (.o(FE_OFN483_n249211),
	.a(n249211));
   in01f01 FE_OFC478_n249800 (.o(FE_OFN478_n249800),
	.a(FE_OFN477_n249800));
   in01f01 FE_OFC477_n249800 (.o(FE_OFN477_n249800),
	.a(n249800));
   in01f01 FE_OFC472_n244982 (.o(FE_OFN472_n244982),
	.a(FE_OFN471_n244982));
   in01f01 FE_OFC471_n244982 (.o(FE_OFN471_n244982),
	.a(n244982));
   in01f01 FE_OFC470_n244978 (.o(FE_OFN470_n244978),
	.a(FE_OFN469_n244978));
   in01f01 FE_OFC469_n244978 (.o(FE_OFN469_n244978),
	.a(n244978));
   in01f01 FE_OFC468_n244218 (.o(FE_OFN468_n244218),
	.a(FE_OFN467_n244218));
   in01f01 FE_OFC467_n244218 (.o(FE_OFN467_n244218),
	.a(n244218));
   in01f01 FE_OFC466_n249845 (.o(FE_OFN466_n249845),
	.a(FE_OFN465_n249845));
   in01f01 FE_OFC465_n249845 (.o(FE_OFN465_n249845),
	.a(n249845));
   in01f02 FE_OFC464_n249821 (.o(FE_OFN464_n249821),
	.a(FE_OFN463_n249821));
   in01f01 FE_OFC463_n249821 (.o(FE_OFN463_n249821),
	.a(n249821));
   in01f01 FE_OFC462_n249378 (.o(FE_OFN462_n249378),
	.a(FE_OFN461_n249378));
   in01f01 FE_OFC461_n249378 (.o(FE_OFN461_n249378),
	.a(n249378));
   in01f04 FE_OFC458_n252996 (.o(FE_OFN458_n252996),
	.a(FE_OFN457_n252996));
   in01f01 FE_OFC457_n252996 (.o(FE_OFN457_n252996),
	.a(n252996));
   in01f04 FE_OFC456_n252942 (.o(FE_OFN456_n252942),
	.a(FE_OFN455_n252942));
   in01f01 FE_OFC455_n252942 (.o(FE_OFN455_n252942),
	.a(n252942));
   in01f06 FE_OFC454_n252863 (.o(FE_OFN454_n252863),
	.a(FE_OFN453_n252863));
   in01f01 FE_OFC453_n252863 (.o(FE_OFN453_n252863),
	.a(n252863));
   in01f01 FE_OFC449_n249831 (.o(FE_OFN449_n249831),
	.a(FE_OFN448_n249831));
   in01f01 FE_OFC448_n249831 (.o(FE_OFN448_n249831),
	.a(n249831));
   in01f01 FE_OFC445_n249391 (.o(FE_OFN445_n249391),
	.a(FE_OFN444_n249391));
   in01f01 FE_OFC444_n249391 (.o(FE_OFN444_n249391),
	.a(n249391));
   in01f06 FE_OFC441_n252905 (.o(FE_OFN441_n252905),
	.a(FE_OFN440_n252905));
   in01f01 FE_OFC440_n252905 (.o(FE_OFN440_n252905),
	.a(n252905));
   in01f02 FE_OFC439_n252264 (.o(FE_OFN439_n252264),
	.a(n252270));
   in01f04 FE_OFC437_n252069 (.o(FE_OFN437_n252069),
	.a(FE_OFN435_n252069));
   in01f03 FE_OFC436_n252069 (.o(FE_OFN436_n252069),
	.a(FE_OFN435_n252069));
   in01f01 FE_OFC435_n252069 (.o(FE_OFN435_n252069),
	.a(n252069));
   in01f08 FE_OFC434_n251996 (.o(FE_OFN434_n251996),
	.a(FE_OFN433_n251996));
   in01f01 FE_OFC433_n251996 (.o(FE_OFN433_n251996),
	.a(n251996));
   in01f08 FE_OFC432_n251781 (.o(FE_OFN432_n251781),
	.a(FE_OFN431_n251781));
   in01f01 FE_OFC431_n251781 (.o(FE_OFN431_n251781),
	.a(n251781));
   in01f06 FE_OFC430_n251710 (.o(FE_OFN430_n251710),
	.a(FE_OFN429_n251710));
   in01f01 FE_OFC429_n251710 (.o(FE_OFN429_n251710),
	.a(n251710));
   in01f08 FE_OFC428_n251494 (.o(FE_OFN428_n251494),
	.a(FE_OFN427_n251494));
   in01f01 FE_OFC427_n251494 (.o(FE_OFN427_n251494),
	.a(n251494));
   in01f08 FE_OFC426_n251424 (.o(FE_OFN426_n251424),
	.a(FE_OFN425_n251424));
   in01f01 FE_OFC425_n251424 (.o(FE_OFN425_n251424),
	.a(n251424));
   in01f06 FE_OFC424_n251300 (.o(FE_OFN424_n251300),
	.a(FE_OFN423_n251300));
   in01f01 FE_OFC423_n251300 (.o(FE_OFN423_n251300),
	.a(n251300));
   in01f06 FE_OFC422_n251211 (.o(FE_OFN422_n251211),
	.a(FE_OFN421_n251211));
   in01f01 FE_OFC421_n251211 (.o(FE_OFN421_n251211),
	.a(n251211));
   in01f08 FE_OFC420_n251140 (.o(FE_OFN420_n251140),
	.a(FE_OFN419_n251140));
   in01f01 FE_OFC419_n251140 (.o(FE_OFN419_n251140),
	.a(n251140));
   in01f08 FE_OFC418_n250930 (.o(FE_OFN418_n250930),
	.a(FE_OFN417_n250930));
   in01f01 FE_OFC417_n250930 (.o(FE_OFN417_n250930),
	.a(n250930));
   in01f08 FE_OFC416_n250859 (.o(FE_OFN416_n250859),
	.a(FE_OFN415_n250859));
   in01f01 FE_OFC415_n250859 (.o(FE_OFN415_n250859),
	.a(n250859));
   in01f08 FE_OFC414_n250646 (.o(FE_OFN414_n250646),
	.a(FE_OFN413_n250646));
   in01f01 FE_OFC413_n250646 (.o(FE_OFN413_n250646),
	.a(n250646));
   in01f08 FE_OFC412_n250576 (.o(FE_OFN412_n250576),
	.a(FE_OFN411_n250576));
   in01f01 FE_OFC411_n250576 (.o(FE_OFN411_n250576),
	.a(n250576));
   in01f08 FE_OFC410_n250360 (.o(FE_OFN410_n250360),
	.a(FE_OFN409_n250360));
   in01f01 FE_OFC409_n250360 (.o(FE_OFN409_n250360),
	.a(n250360));
   in01f08 FE_OFC408_n250289 (.o(FE_OFN408_n250289),
	.a(FE_OFN407_n250289));
   in01f01 FE_OFC407_n250289 (.o(FE_OFN407_n250289),
	.a(n250289));
   in01f03 FE_OFC406_n250162 (.o(FE_OFN406_n250162),
	.a(FE_OFN405_n250162));
   in01f01 FE_OFC405_n250162 (.o(FE_OFN405_n250162),
	.a(n250162));
   in01f06 FE_OFC404_n250071 (.o(FE_OFN404_n250071),
	.a(FE_OFN403_n250071));
   in01f01 FE_OFC403_n250071 (.o(FE_OFN403_n250071),
	.a(n250071));
   in01f06 FE_OFC402_n249999 (.o(FE_OFN402_n249999),
	.a(FE_OFN401_n249999));
   in01f01 FE_OFC401_n249999 (.o(FE_OFN401_n249999),
	.a(n249999));
   in01f02 FE_OFC400_n249836 (.o(FE_OFN400_n249836),
	.a(FE_OFN399_n249836));
   in01f01 FE_OFC399_n249836 (.o(FE_OFN399_n249836),
	.a(n249836));
   in01f04 FE_OFC398_n249646 (.o(FE_OFN398_n249646),
	.a(FE_OFN397_n249646));
   in01f01 FE_OFC397_n249646 (.o(FE_OFN397_n249646),
	.a(n249646));
   in01f03 FE_OFC396_n249640 (.o(FE_OFN396_n249640),
	.a(FE_OFN395_n249640));
   in01f01 FE_OFC395_n249640 (.o(FE_OFN395_n249640),
	.a(n249640));
   in01f02 FE_OFC392_n249635 (.o(FE_OFN392_n249635),
	.a(FE_OFN391_n249635));
   in01f01 FE_OFC391_n249635 (.o(FE_OFN391_n249635),
	.a(n249635));
   in01f01 FE_OFC390_n249480 (.o(FE_OFN390_n249480),
	.a(FE_OFN389_n249480));
   in01f01 FE_OFC389_n249480 (.o(FE_OFN389_n249480),
	.a(n249480));
   in01f01 FE_OFC388_n249468 (.o(FE_OFN388_n249468),
	.a(FE_OFN387_n249468));
   in01f01 FE_OFC387_n249468 (.o(FE_OFN387_n249468),
	.a(n249468));
   in01f02 FE_OFC386_n248760 (.o(FE_OFN386_n248760),
	.a(FE_OFN385_n248760));
   in01f01 FE_OFC385_n248760 (.o(FE_OFN385_n248760),
	.a(n248760));
   in01f01 FE_OFC384_n248677 (.o(FE_OFN384_n248677),
	.a(FE_OFN383_n248677));
   in01f01 FE_OFC383_n248677 (.o(FE_OFN383_n248677),
	.a(n248677));
   in01f01 FE_OFC382_n248549 (.o(FE_OFN382_n248549),
	.a(FE_OFN381_n248549));
   in01f01 FE_OFC381_n248549 (.o(FE_OFN381_n248549),
	.a(n248549));
   in01f02 FE_OFC376_n248352 (.o(FE_OFN376_n248352),
	.a(FE_OFN375_n248352));
   in01f01 FE_OFC375_n248352 (.o(FE_OFN375_n248352),
	.a(n248352));
   in01f02 FE_OFC374_n248311 (.o(FE_OFN374_n248311),
	.a(FE_OFN373_n248311));
   in01f01 FE_OFC373_n248311 (.o(FE_OFN373_n248311),
	.a(n248311));
   in01f01 FE_OFC372_n247737 (.o(FE_OFN372_n247737),
	.a(FE_OFN371_n247737));
   in01f01 FE_OFC371_n247737 (.o(FE_OFN371_n247737),
	.a(n247737));
   in01f02 FE_OFC368_n247123 (.o(FE_OFN368_n247123),
	.a(FE_OFN367_n247123));
   in01f01 FE_OFC367_n247123 (.o(FE_OFN367_n247123),
	.a(n247123));
   in01f06 FE_OFC366_n246266 (.o(FE_OFN366_n246266),
	.a(FE_OFN365_n246266));
   in01f01 FE_OFC365_n246266 (.o(FE_OFN365_n246266),
	.a(n246266));
   in01f08 FE_OFC362_n252748 (.o(FE_OFN362_n252748),
	.a(FE_OFN361_n252748));
   in01f01 FE_OFC361_n252748 (.o(FE_OFN361_n252748),
	.a(n252748));
   in01f04 FE_OFC360_n252728 (.o(FE_OFN360_n252728),
	.a(FE_OFN359_n252728));
   in01f01 FE_OFC359_n252728 (.o(FE_OFN359_n252728),
	.a(n252728));
   in01f04 FE_OFC356_n252508 (.o(FE_OFN356_n252508),
	.a(FE_OFN355_n252508));
   in01f01 FE_OFC355_n252508 (.o(FE_OFN355_n252508),
	.a(n252508));
   in01f06 FE_OFC354_n252338 (.o(FE_OFN354_n252338),
	.a(FE_OFN353_n252338));
   in01f01 FE_OFC353_n252338 (.o(FE_OFN353_n252338),
	.a(n252338));
   in01f01 FE_OFC352_n252242 (.o(FE_OFN352_n252242),
	.a(FE_OFN351_n252242));
   in01f01 FE_OFC351_n252242 (.o(FE_OFN351_n252242),
	.a(n252242));
   in01f08 FE_OFC350_n252215 (.o(FE_OFN350_n252215),
	.a(FE_OFN349_n252215));
   in01f01 FE_OFC349_n252215 (.o(FE_OFN349_n252215),
	.a(n252215));
   in01f08 FE_OFC348_n252178 (.o(FE_OFN348_n252178),
	.a(FE_OFN347_n252178));
   in01f01 FE_OFC347_n252178 (.o(FE_OFN347_n252178),
	.a(n252178));
   in01f06 FE_OFC346_n252141 (.o(FE_OFN346_n252141),
	.a(FE_OFN344_n252141));
   in01f03 FE_OFC345_n252141 (.o(FE_OFN345_n252141),
	.a(FE_OFN344_n252141));
   in01f02 FE_OFC344_n252141 (.o(FE_OFN344_n252141),
	.a(n252141));
   in01f06 FE_OFC343_n252032 (.o(FE_OFN343_n252032),
	.a(FE_OFN342_n252032));
   in01f01 FE_OFC342_n252032 (.o(FE_OFN342_n252032),
	.a(n252032));
   in01f06 FE_OFC341_n251960 (.o(FE_OFN341_n251960),
	.a(FE_OFN340_n251960));
   in01f01 FE_OFC340_n251960 (.o(FE_OFN340_n251960),
	.a(n251960));
   in01f08 FE_OFC339_n251923 (.o(FE_OFN339_n251923),
	.a(FE_OFN338_n251923));
   in01f01 FE_OFC338_n251923 (.o(FE_OFN338_n251923),
	.a(n251923));
   in01f06 FE_OFC337_n251887 (.o(FE_OFN337_n251887),
	.a(FE_OFN336_n251887));
   in01f01 FE_OFC336_n251887 (.o(FE_OFN336_n251887),
	.a(n251887));
   in01f06 FE_OFC335_n251852 (.o(FE_OFN335_n251852),
	.a(FE_OFN334_n251852));
   in01f01 FE_OFC334_n251852 (.o(FE_OFN334_n251852),
	.a(n251852));
   in01f06 FE_OFC333_n251746 (.o(FE_OFN333_n251746),
	.a(FE_OFN332_n251746));
   in01f01 FE_OFC332_n251746 (.o(FE_OFN332_n251746),
	.a(n251746));
   in01f08 FE_OFC331_n251675 (.o(FE_OFN331_n251675),
	.a(FE_OFN330_n251675));
   in01f01 FE_OFC330_n251675 (.o(FE_OFN330_n251675),
	.a(n251675));
   in01f08 FE_OFC329_n251637 (.o(FE_OFN329_n251637),
	.a(FE_OFN328_n251637));
   in01f01 FE_OFC328_n251637 (.o(FE_OFN328_n251637),
	.a(n251637));
   in01f08 FE_OFC327_n251600 (.o(FE_OFN327_n251600),
	.a(FE_OFN326_n251600));
   in01f01 FE_OFC326_n251600 (.o(FE_OFN326_n251600),
	.a(n251600));
   in01f06 FE_OFC325_n251565 (.o(FE_OFN325_n251565),
	.a(FE_OFN323_n251565));
   in01f03 FE_OFC324_n251565 (.o(FE_OFN324_n251565),
	.a(FE_OFN323_n251565));
   in01f02 FE_OFC323_n251565 (.o(FE_OFN323_n251565),
	.a(n251565));
   in01f08 FE_OFC322_n251459 (.o(FE_OFN322_n251459),
	.a(FE_OFN321_n251459));
   in01f01 FE_OFC321_n251459 (.o(FE_OFN321_n251459),
	.a(n251459));
   in01f06 FE_OFC320_n251388 (.o(FE_OFN320_n251388),
	.a(FE_OFN319_n251388));
   in01f01 FE_OFC319_n251388 (.o(FE_OFN319_n251388),
	.a(n251388));
   in01f08 FE_OFC318_n251353 (.o(FE_OFN318_n251353),
	.a(FE_OFN317_n251353));
   in01f01 FE_OFC317_n251353 (.o(FE_OFN317_n251353),
	.a(n251353));
   in01f08 FE_OFC316_n251317 (.o(FE_OFN316_n251317),
	.a(FE_OFN315_n251317));
   in01f01 FE_OFC315_n251317 (.o(FE_OFN315_n251317),
	.a(n251317));
   in01f06 FE_OFC314_n251281 (.o(FE_OFN314_n251281),
	.a(FE_OFN312_n251281));
   in01f03 FE_OFC313_n251281 (.o(FE_OFN313_n251281),
	.a(FE_OFN312_n251281));
   in01f02 FE_OFC312_n251281 (.o(FE_OFN312_n251281),
	.a(n251281));
   in01f08 FE_OFC311_n251175 (.o(FE_OFN311_n251175),
	.a(FE_OFN310_n251175));
   in01f01 FE_OFC310_n251175 (.o(FE_OFN310_n251175),
	.a(n251175));
   in01f06 FE_OFC309_n251105 (.o(FE_OFN309_n251105),
	.a(FE_OFN308_n251105));
   in01f01 FE_OFC308_n251105 (.o(FE_OFN308_n251105),
	.a(n251105));
   in01f06 FE_OFC307_n251072 (.o(FE_OFN307_n251072),
	.a(FE_OFN305_n251072));
   in01f03 FE_OFC306_n251072 (.o(FE_OFN306_n251072),
	.a(FE_OFN305_n251072));
   in01f02 FE_OFC305_n251072 (.o(FE_OFN305_n251072),
	.a(n251072));
   in01f08 FE_OFC304_n251036 (.o(FE_OFN304_n251036),
	.a(FE_OFN303_n251036));
   in01f01 FE_OFC303_n251036 (.o(FE_OFN303_n251036),
	.a(n251036));
   in01f08 FE_OFC302_n251001 (.o(FE_OFN302_n251001),
	.a(FE_OFN301_n251001));
   in01f01 FE_OFC301_n251001 (.o(FE_OFN301_n251001),
	.a(n251001));
   in01f08 FE_OFC300_n250895 (.o(FE_OFN300_n250895),
	.a(FE_OFN299_n250895));
   in01f01 FE_OFC299_n250895 (.o(FE_OFN299_n250895),
	.a(n250895));
   in01f06 FE_OFC298_n250824 (.o(FE_OFN298_n250824),
	.a(FE_OFN297_n250824));
   in01f01 FE_OFC297_n250824 (.o(FE_OFN297_n250824),
	.a(n250824));
   in01f08 FE_OFC296_n250789 (.o(FE_OFN296_n250789),
	.a(FE_OFN295_n250789));
   in01f01 FE_OFC295_n250789 (.o(FE_OFN295_n250789),
	.a(n250789));
   in01f08 FE_OFC294_n250752 (.o(FE_OFN294_n250752),
	.a(FE_OFN293_n250752));
   in01f01 FE_OFC293_n250752 (.o(FE_OFN293_n250752),
	.a(n250752));
   in01f06 FE_OFC292_n250717 (.o(FE_OFN292_n250717),
	.a(FE_OFN291_n250717));
   in01f01 FE_OFC291_n250717 (.o(FE_OFN291_n250717),
	.a(n250717));
   in01f08 FE_OFC290_n250611 (.o(FE_OFN290_n250611),
	.a(FE_OFN289_n250611));
   in01f01 FE_OFC289_n250611 (.o(FE_OFN289_n250611),
	.a(n250611));
   in01f06 FE_OFC288_n250540 (.o(FE_OFN288_n250540),
	.a(FE_OFN287_n250540));
   in01f01 FE_OFC287_n250540 (.o(FE_OFN287_n250540),
	.a(n250540));
   in01f04 FE_OFC286_n250502 (.o(FE_OFN286_n250502),
	.a(FE_OFN285_n250502));
   in01f01 FE_OFC285_n250502 (.o(FE_OFN285_n250502),
	.a(n250502));
   in01f06 FE_OFC284_n250466 (.o(FE_OFN284_n250466),
	.a(FE_OFN283_n250466));
   in01f01 FE_OFC283_n250466 (.o(FE_OFN283_n250466),
	.a(n250466));
   in01f08 FE_OFC282_n250430 (.o(FE_OFN282_n250430),
	.a(FE_OFN281_n250430));
   in01f01 FE_OFC281_n250430 (.o(FE_OFN281_n250430),
	.a(n250430));
   in01f08 FE_OFC280_n250324 (.o(FE_OFN280_n250324),
	.a(FE_OFN279_n250324));
   in01f01 FE_OFC279_n250324 (.o(FE_OFN279_n250324),
	.a(n250324));
   in01f06 FE_OFC278_n250254 (.o(FE_OFN278_n250254),
	.a(FE_OFN277_n250254));
   in01f01 FE_OFC277_n250254 (.o(FE_OFN277_n250254),
	.a(n250254));
   in01f08 FE_OFC276_n250218 (.o(FE_OFN276_n250218),
	.a(FE_OFN275_n250218));
   in01f01 FE_OFC275_n250218 (.o(FE_OFN275_n250218),
	.a(n250218));
   in01f08 FE_OFC274_n250180 (.o(FE_OFN274_n250180),
	.a(FE_OFN273_n250180));
   in01f01 FE_OFC273_n250180 (.o(FE_OFN273_n250180),
	.a(n250180));
   in01f08 FE_OFC272_n250144 (.o(FE_OFN272_n250144),
	.a(FE_OFN271_n250144));
   in01f01 FE_OFC271_n250144 (.o(FE_OFN271_n250144),
	.a(n250144));
   in01f06 FE_OFC270_n250035 (.o(FE_OFN270_n250035),
	.a(FE_OFN269_n250035));
   in01f01 FE_OFC269_n250035 (.o(FE_OFN269_n250035),
	.a(n250035));
   in01f06 FE_OFC268_n249964 (.o(FE_OFN268_n249964),
	.a(FE_OFN267_n249964));
   in01f01 FE_OFC267_n249964 (.o(FE_OFN267_n249964),
	.a(n249964));
   in01f02 FE_OFC266_n249787 (.o(FE_OFN266_n249787),
	.a(FE_OFN265_n249787));
   in01f01 FE_OFC265_n249787 (.o(FE_OFN265_n249787),
	.a(n249787));
   in01f04 FE_OFC264_n249636 (.o(FE_OFN264_n249636),
	.a(FE_OFN263_n249636));
   in01f01 FE_OFC263_n249636 (.o(FE_OFN263_n249636),
	.a(n249636));
   in01f02 FE_OFC256_n248843 (.o(FE_OFN256_n248843),
	.a(FE_OFN255_n248843));
   in01f01 FE_OFC255_n248843 (.o(FE_OFN255_n248843),
	.a(n248843));
   in01f01 FE_OFC252_n248799 (.o(FE_OFN252_n248799),
	.a(FE_OFN251_n248799));
   in01f01 FE_OFC251_n248799 (.o(FE_OFN251_n248799),
	.a(n248799));
   in01f01 FE_OFC248_n248527 (.o(FE_OFN248_n248527),
	.a(FE_OFN247_n248527));
   in01f01 FE_OFC247_n248527 (.o(FE_OFN247_n248527),
	.a(n248527));
   in01f01 FE_OFC246_n248465 (.o(FE_OFN246_n248465),
	.a(FE_OFN245_n248465));
   in01f01 FE_OFC245_n248465 (.o(FE_OFN245_n248465),
	.a(n248465));
   in01f01 FE_OFC244_n248463 (.o(FE_OFN244_n248463),
	.a(FE_OFN243_n248463));
   in01f01 FE_OFC243_n248463 (.o(FE_OFN243_n248463),
	.a(n248463));
   in01f01 FE_OFC240_n248389 (.o(FE_OFN240_n248389),
	.a(FE_OFN239_n248389));
   in01f01 FE_OFC239_n248389 (.o(FE_OFN239_n248389),
	.a(n248389));
   in01f01 FE_OFC236_n248245 (.o(FE_OFN236_n248245),
	.a(FE_OFN235_n248245));
   in01f01 FE_OFC235_n248245 (.o(FE_OFN235_n248245),
	.a(n248245));
   in01f02 FE_OFC234_n248115 (.o(FE_OFN234_n248115),
	.a(FE_OFN233_n248115));
   in01f01 FE_OFC233_n248115 (.o(FE_OFN233_n248115),
	.a(n248115));
   in01f01 FE_OFC230_n247987 (.o(FE_OFN230_n247987),
	.a(FE_OFN229_n247987));
   in01f01 FE_OFC229_n247987 (.o(FE_OFN229_n247987),
	.a(n247987));
   in01f01 FE_OFC228_n247903 (.o(FE_OFN228_n247903),
	.a(FE_OFN227_n247903));
   in01f01 FE_OFC227_n247903 (.o(FE_OFN227_n247903),
	.a(n247903));
   in01f02 FE_OFC220_n246261 (.o(FE_OFN220_n246261),
	.a(FE_OFN219_n246261));
   in01f01 FE_OFC219_n246261 (.o(FE_OFN219_n246261),
	.a(n246261));
   in01f04 FE_OFC218_n246238 (.o(FE_OFN218_n246238),
	.a(FE_OFN217_n246238));
   in01f01 FE_OFC217_n246238 (.o(FE_OFN217_n246238),
	.a(n246238));
   in01f08 FE_OFC214_n252483 (.o(FE_OFN214_n252483),
	.a(FE_OFN213_n252483));
   in01f01 FE_OFC213_n252483 (.o(FE_OFN213_n252483),
	.a(n252483));
   in01f04 FE_OFC212_n252422 (.o(FE_OFN212_n252422),
	.a(FE_OFN211_n252422));
   in01f01 FE_OFC211_n252422 (.o(FE_OFN211_n252422),
	.a(n252422));
   in01f02 FE_OFC210_n252159 (.o(FE_OFN210_n252159),
	.a(FE_OFN209_n252159));
   in01f01 FE_OFC209_n252159 (.o(FE_OFN209_n252159),
	.a(n252159));
   in01f08 FE_OFC208_n252105 (.o(FE_OFN208_n252105),
	.a(FE_OFN207_n252105));
   in01f01 FE_OFC207_n252105 (.o(FE_OFN207_n252105),
	.a(n252105));
   in01f08 FE_OFC206_n251816 (.o(FE_OFN206_n251816),
	.a(FE_OFN205_n251816));
   in01f01 FE_OFC205_n251816 (.o(FE_OFN205_n251816),
	.a(n251816));
   in01f08 FE_OFC204_n251530 (.o(FE_OFN204_n251530),
	.a(FE_OFN203_n251530));
   in01f01 FE_OFC203_n251530 (.o(FE_OFN203_n251530),
	.a(n251530));
   in01f06 FE_OFC202_n251246 (.o(FE_OFN202_n251246),
	.a(FE_OFN201_n251246));
   in01f01 FE_OFC201_n251246 (.o(FE_OFN201_n251246),
	.a(n251246));
   in01f08 FE_OFC200_n250965 (.o(FE_OFN200_n250965),
	.a(FE_OFN199_n250965));
   in01f01 FE_OFC199_n250965 (.o(FE_OFN199_n250965),
	.a(n250965));
   in01f04 FE_OFC198_n250682 (.o(FE_OFN198_n250682),
	.a(FE_OFN196_n250682));
   in01f02 FE_OFC197_n250682 (.o(FE_OFN197_n250682),
	.a(FE_OFN196_n250682));
   in01f01 FE_OFC196_n250682 (.o(FE_OFN196_n250682),
	.a(n250682));
   in01f08 FE_OFC195_n250395 (.o(FE_OFN195_n250395),
	.a(FE_OFN194_n250395));
   in01f01 FE_OFC194_n250395 (.o(FE_OFN194_n250395),
	.a(n250395));
   in01f04 FE_OFC193_n250107 (.o(FE_OFN193_n250107),
	.a(FE_OFN191_n250107));
   in01f03 FE_OFC192_n250107 (.o(FE_OFN192_n250107),
	.a(FE_OFN191_n250107));
   in01f01 FE_OFC191_n250107 (.o(FE_OFN191_n250107),
	.a(n250107));
   in01f08 FE_OFC185_n248415 (.o(FE_OFN185_n248415),
	.a(FE_OFN184_n248415));
   in01f01 FE_OFC184_n248415 (.o(FE_OFN184_n248415),
	.a(n248415));
   in01f08 FE_OFC183_n248414 (.o(FE_OFN183_n248414),
	.a(FE_OFN182_n248414));
   in01f01 FE_OFC182_n248414 (.o(FE_OFN182_n248414),
	.a(n248414));
   in01f08 FE_OFC181_n248413 (.o(FE_OFN181_n248413),
	.a(FE_OFN180_n248413));
   in01f01 FE_OFC180_n248413 (.o(FE_OFN180_n248413),
	.a(n248413));
   in01f08 FE_OFC179_n248408 (.o(FE_OFN179_n248408),
	.a(FE_OFN178_n248408));
   in01f01 FE_OFC178_n248408 (.o(FE_OFN178_n248408),
	.a(n248408));
   in01f08 FE_OFC177_n248407 (.o(FE_OFN177_n248407),
	.a(FE_OFN176_n248407));
   in01f01 FE_OFC176_n248407 (.o(FE_OFN176_n248407),
	.a(n248407));
   in01f08 FE_OFC175_n248406 (.o(FE_OFN175_n248406),
	.a(FE_OFN174_n248406));
   in01f01 FE_OFC174_n248406 (.o(FE_OFN174_n248406),
	.a(n248406));
   in01f08 FE_OFC173_n248405 (.o(FE_OFN173_n248405),
	.a(FE_OFN172_n248405));
   in01f01 FE_OFC172_n248405 (.o(FE_OFN172_n248405),
	.a(n248405));
   in01f08 FE_OFC171_n248404 (.o(FE_OFN171_n248404),
	.a(FE_OFN170_n248404));
   in01f01 FE_OFC170_n248404 (.o(FE_OFN170_n248404),
	.a(n248404));
   in01f06 FE_OFC169_n248399 (.o(FE_OFN169_n248399),
	.a(FE_OFN168_n248399));
   in01f01 FE_OFC168_n248399 (.o(FE_OFN168_n248399),
	.a(n248399));
   in01f06 FE_OFC167_n248398 (.o(FE_OFN167_n248398),
	.a(FE_OFN166_n248398));
   in01f01 FE_OFC166_n248398 (.o(FE_OFN166_n248398),
	.a(n248398));
   in01f08 FE_OFC165_n248393 (.o(FE_OFN165_n248393),
	.a(FE_OFN164_n248393));
   in01f01 FE_OFC164_n248393 (.o(FE_OFN164_n248393),
	.a(n248393));
   in01f08 FE_OFC163_n248392 (.o(FE_OFN163_n248392),
	.a(FE_OFN162_n248392));
   in01f01 FE_OFC162_n248392 (.o(FE_OFN162_n248392),
	.a(n248392));
   in01f08 FE_OFC161_n248391 (.o(FE_OFN161_n248391),
	.a(FE_OFN160_n248391));
   in01f01 FE_OFC160_n248391 (.o(FE_OFN160_n248391),
	.a(n248391));
   in01f06 FE_OFC159_n248382 (.o(FE_OFN159_n248382),
	.a(FE_OFN158_n248382));
   in01f01 FE_OFC158_n248382 (.o(FE_OFN158_n248382),
	.a(n248382));
   in01f08 FE_OFC157_n248381 (.o(FE_OFN157_n248381),
	.a(FE_OFN156_n248381));
   in01f01 FE_OFC156_n248381 (.o(FE_OFN156_n248381),
	.a(n248381));
   in01f08 FE_OFC155_n248380 (.o(FE_OFN155_n248380),
	.a(FE_OFN154_n248380));
   in01f01 FE_OFC154_n248380 (.o(FE_OFN154_n248380),
	.a(n248380));
   in01f06 FE_OFC153_n248375 (.o(FE_OFN153_n248375),
	.a(FE_OFN152_n248375));
   in01f01 FE_OFC152_n248375 (.o(FE_OFN152_n248375),
	.a(n248375));
   in01f06 FE_OFC151_n248374 (.o(FE_OFN151_n248374),
	.a(FE_OFN150_n248374));
   in01f01 FE_OFC150_n248374 (.o(FE_OFN150_n248374),
	.a(n248374));
   in01f06 FE_OFC149_n248373 (.o(FE_OFN149_n248373),
	.a(FE_OFN148_n248373));
   in01f01 FE_OFC148_n248373 (.o(FE_OFN148_n248373),
	.a(n248373));
   in01f06 FE_OFC147_n248372 (.o(FE_OFN147_n248372),
	.a(FE_OFN145_n248372));
   in01f01 FE_OFC146_n248372 (.o(FE_OFN146_n248372),
	.a(FE_OFN145_n248372));
   in01f01 FE_OFC145_n248372 (.o(FE_OFN145_n248372),
	.a(n248372));
   in01f06 FE_OFC144_n248371 (.o(FE_OFN144_n248371),
	.a(FE_OFN143_n248371));
   in01f01 FE_OFC143_n248371 (.o(FE_OFN143_n248371),
	.a(n248371));
   in01f06 FE_OFC142_n248370 (.o(FE_OFN142_n248370),
	.a(FE_OFN141_n248370));
   in01f01 FE_OFC141_n248370 (.o(FE_OFN141_n248370),
	.a(n248370));
   in01f06 FE_OFC140_n248369 (.o(FE_OFN140_n248369),
	.a(FE_OFN139_n248369));
   in01f01 FE_OFC139_n248369 (.o(FE_OFN139_n248369),
	.a(n248369));
   in01f06 FE_OFC138_n248364 (.o(FE_OFN138_n248364),
	.a(FE_OFN137_n248364));
   in01f01 FE_OFC137_n248364 (.o(FE_OFN137_n248364),
	.a(n248364));
   in01f08 FE_OFC136_n248363 (.o(FE_OFN136_n248363),
	.a(FE_OFN135_n248363));
   in01f01 FE_OFC135_n248363 (.o(FE_OFN135_n248363),
	.a(n248363));
   in01f08 FE_OFC134_n248362 (.o(FE_OFN134_n248362),
	.a(FE_OFN133_n248362));
   in01f01 FE_OFC133_n248362 (.o(FE_OFN133_n248362),
	.a(n248362));
   in01f08 FE_OFC132_n248357 (.o(FE_OFN132_n248357),
	.a(FE_OFN131_n248357));
   in01f01 FE_OFC131_n248357 (.o(FE_OFN131_n248357),
	.a(n248357));
   in01f08 FE_OFC130_n248356 (.o(FE_OFN130_n248356),
	.a(FE_OFN129_n248356));
   in01f01 FE_OFC129_n248356 (.o(FE_OFN129_n248356),
	.a(n248356));
   in01f08 FE_OFC128_n248355 (.o(FE_OFN128_n248355),
	.a(FE_OFN127_n248355));
   in01f01 FE_OFC127_n248355 (.o(FE_OFN127_n248355),
	.a(n248355));
   in01f08 FE_OFC126_n248176 (.o(FE_OFN126_n248176),
	.a(FE_OFN125_n248176));
   in01f01 FE_OFC125_n248176 (.o(FE_OFN125_n248176),
	.a(n248176));
   in01f08 FE_OFC124_n248175 (.o(FE_OFN124_n248175),
	.a(FE_OFN123_n248175));
   in01f01 FE_OFC123_n248175 (.o(FE_OFN123_n248175),
	.a(n248175));
   in01f08 FE_OFC122_n248174 (.o(FE_OFN122_n248174),
	.a(FE_OFN121_n248174));
   in01f01 FE_OFC121_n248174 (.o(FE_OFN121_n248174),
	.a(n248174));
   in01f08 FE_OFC120_n248173 (.o(FE_OFN120_n248173),
	.a(FE_OFN119_n248173));
   in01f01 FE_OFC119_n248173 (.o(FE_OFN119_n248173),
	.a(n248173));
   in01f08 FE_OFC116_n248167 (.o(FE_OFN116_n248167),
	.a(FE_OFN115_n248167));
   in01f01 FE_OFC115_n248167 (.o(FE_OFN115_n248167),
	.a(n248167));
   in01f06 FE_OFC114_n248162 (.o(FE_OFN114_n248162),
	.a(FE_OFN112_n248162));
   in01f01 FE_OFC113_n248162 (.o(FE_OFN113_n248162),
	.a(FE_OFN112_n248162));
   in01f01 FE_OFC112_n248162 (.o(FE_OFN112_n248162),
	.a(n248162));
   in01f06 FE_OFC109_n248160 (.o(FE_OFN109_n248160),
	.a(FE_OFN107_n248160));
   in01f01 FE_OFC108_n248160 (.o(FE_OFN108_n248160),
	.a(FE_OFN107_n248160));
   in01f01 FE_OFC107_n248160 (.o(FE_OFN107_n248160),
	.a(n248160));
   in01f08 FE_OFC106_n248159 (.o(FE_OFN106_n248159),
	.a(FE_OFN105_n248159));
   in01f01 FE_OFC105_n248159 (.o(FE_OFN105_n248159),
	.a(n248159));
   in01f08 FE_OFC104_n248158 (.o(FE_OFN104_n248158),
	.a(FE_OFN103_n248158));
   in01f01 FE_OFC103_n248158 (.o(FE_OFN103_n248158),
	.a(n248158));
   in01f08 FE_OFC102_n248153 (.o(FE_OFN102_n248153),
	.a(FE_OFN101_n248153));
   in01f01 FE_OFC101_n248153 (.o(FE_OFN101_n248153),
	.a(n248153));
   in01f08 FE_OFC100_n248152 (.o(FE_OFN100_n248152),
	.a(FE_OFN99_n248152));
   in01f01 FE_OFC99_n248152 (.o(FE_OFN99_n248152),
	.a(n248152));
   in01f08 FE_OFC98_n248151 (.o(FE_OFN98_n248151),
	.a(FE_OFN97_n248151));
   in01f01 FE_OFC97_n248151 (.o(FE_OFN97_n248151),
	.a(n248151));
   in01f08 FE_OFC96_n248150 (.o(FE_OFN96_n248150),
	.a(FE_OFN95_n248150));
   in01f01 FE_OFC95_n248150 (.o(FE_OFN95_n248150),
	.a(n248150));
   in01f06 FE_OFC94_n248141 (.o(FE_OFN94_n248141),
	.a(FE_OFN93_n248141));
   in01f01 FE_OFC93_n248141 (.o(FE_OFN93_n248141),
	.a(n248141));
   in01f06 FE_OFC90_n248139 (.o(FE_OFN90_n248139),
	.a(FE_OFN89_n248139));
   in01f01 FE_OFC89_n248139 (.o(FE_OFN89_n248139),
	.a(n248139));
   in01f08 FE_OFC88_n248138 (.o(FE_OFN88_n248138),
	.a(FE_OFN87_n248138));
   in01f01 FE_OFC87_n248138 (.o(FE_OFN87_n248138),
	.a(n248138));
   in01f06 FE_OFC86_n248129 (.o(FE_OFN86_n248129),
	.a(FE_OFN85_n248129));
   in01f01 FE_OFC85_n248129 (.o(FE_OFN85_n248129),
	.a(n248129));
   in01f08 FE_OFC84_n248128 (.o(FE_OFN84_n248128),
	.a(FE_OFN83_n248128));
   in01f01 FE_OFC83_n248128 (.o(FE_OFN83_n248128),
	.a(n248128));
   in01f06 FE_OFC82_n248127 (.o(FE_OFN82_n248127),
	.a(FE_OFN80_n248127));
   in01f01 FE_OFC81_n248127 (.o(FE_OFN81_n248127),
	.a(FE_OFN80_n248127));
   in01f01 FE_OFC80_n248127 (.o(FE_OFN80_n248127),
	.a(n248127));
   in01f08 FE_OFC79_n248126 (.o(FE_OFN79_n248126),
	.a(FE_OFN78_n248126));
   in01f01 FE_OFC78_n248126 (.o(FE_OFN78_n248126),
	.a(n248126));
   in01f08 FE_OFC77_n248121 (.o(FE_OFN77_n248121),
	.a(FE_OFN76_n248121));
   in01f01 FE_OFC76_n248121 (.o(FE_OFN76_n248121),
	.a(n248121));
   in01f08 FE_OFC75_n248120 (.o(FE_OFN75_n248120),
	.a(FE_OFN74_n248120));
   in01f01 FE_OFC74_n248120 (.o(FE_OFN74_n248120),
	.a(n248120));
   in01f06 FE_OFC73_n248119 (.o(FE_OFN73_n248119),
	.a(FE_OFN71_n248119));
   in01f03 FE_OFC72_n248119 (.o(FE_OFN72_n248119),
	.a(FE_OFN71_n248119));
   in01f01 FE_OFC71_n248119 (.o(FE_OFN71_n248119),
	.a(n248119));
   in01f08 FE_OFC70_n248118 (.o(FE_OFN70_n248118),
	.a(FE_OFN69_n248118));
   in01f01 FE_OFC69_n248118 (.o(FE_OFN69_n248118),
	.a(n248118));
   in01f08 FE_OFC68_n247591 (.o(FE_OFN68_n247591),
	.a(FE_OFN67_n247591));
   in01f01 FE_OFC67_n247591 (.o(FE_OFN67_n247591),
	.a(n247591));
   in01f08 FE_OFC66_n247531 (.o(FE_OFN66_n247531),
	.a(FE_OFN65_n247531));
   in01f01 FE_OFC65_n247531 (.o(FE_OFN65_n247531),
	.a(n247531));
   in01f06 FE_OFC64_n247509 (.o(FE_OFN64_n247509),
	.a(FE_OFN63_n247509));
   in01f01 FE_OFC63_n247509 (.o(FE_OFN63_n247509),
	.a(n247509));
   in01f08 FE_OFC62_n247107 (.o(FE_OFN62_n247107),
	.a(FE_OFN61_n247107));
   in01f01 FE_OFC61_n247107 (.o(FE_OFN61_n247107),
	.a(n247107));
   in01f06 FE_OFC60_n247099 (.o(FE_OFN60_n247099),
	.a(FE_OFN59_n247099));
   in01f01 FE_OFC59_n247099 (.o(FE_OFN59_n247099),
	.a(n247099));
   in01f08 FE_OFC58_n247092 (.o(FE_OFN58_n247092),
	.a(FE_OFN57_n247092));
   in01f01 FE_OFC57_n247092 (.o(FE_OFN57_n247092),
	.a(n247092));
   in01f06 FE_OFC56_n247074 (.o(FE_OFN56_n247074),
	.a(FE_OFN55_n247074));
   in01f01 FE_OFC55_n247074 (.o(FE_OFN55_n247074),
	.a(n247074));
   in01f03 FE_OFC54_n247067 (.o(FE_OFN54_n247067),
	.a(FE_OFN52_n247067));
   in01f04 FE_OFC53_n247067 (.o(FE_OFN53_n247067),
	.a(FE_OFN52_n247067));
   in01f01 FE_OFC52_n247067 (.o(FE_OFN52_n247067),
	.a(n247067));
   in01f06 FE_OFC51_n247057 (.o(FE_OFN51_n247057),
	.a(FE_OFN50_n247057));
   in01f01 FE_OFC50_n247057 (.o(FE_OFN50_n247057),
	.a(n247057));
   in01f02 FE_OFC45_n252700 (.o(FE_OFN45_n252700),
	.a(FE_OFN44_n252700));
   in01f01 FE_OFC44_n252700 (.o(FE_OFN44_n252700),
	.a(n252700));
   in01f03 FE_OFC43_n252668 (.o(FE_OFN43_n252668),
	.a(FE_OFN42_n252668));
   in01f01 FE_OFC42_n252668 (.o(FE_OFN42_n252668),
	.a(n252668));
   in01f03 FE_OFC41_n252640 (.o(FE_OFN41_n252640),
	.a(FE_OFN40_n252640));
   in01f01 FE_OFC40_n252640 (.o(FE_OFN40_n252640),
	.a(n252640));
   in01f01 FE_OFC39_n252462 (.o(FE_OFN39_n252462),
	.a(FE_OFN38_n252462));
   in01f01 FE_OFC38_n252462 (.o(FE_OFN38_n252462),
	.a(n252462));
   in01f03 FE_OFC37_n252446 (.o(FE_OFN37_n252446),
	.a(FE_OFN36_n252446));
   in01f01 FE_OFC36_n252446 (.o(FE_OFN36_n252446),
	.a(n252446));
   in01f02 FE_OFC33_n251904 (.o(FE_OFN33_n251904),
	.a(FE_OFN31_n251904));
   in01f03 FE_OFC32_n251904 (.o(FE_OFN32_n251904),
	.a(FE_OFN31_n251904));
   in01f01 FE_OFC31_n251904 (.o(FE_OFN31_n251904),
	.a(n251904));
   in01f06 FE_OFC28_n251337 (.o(FE_OFN28_n251337),
	.a(FE_OFN27_n251337));
   in01f01 FE_OFC27_n251337 (.o(FE_OFN27_n251337),
	.a(n251337));
   in01f06 FE_OFC24_n250486 (.o(FE_OFN24_n250486),
	.a(FE_OFN23_n250486));
   in01f01 FE_OFC23_n250486 (.o(FE_OFN23_n250486),
	.a(n250486));
   in01f06 FE_OFC22_n250202 (.o(FE_OFN22_n250202),
	.a(FE_OFN21_n250202));
   in01f01 FE_OFC21_n250202 (.o(FE_OFN21_n250202),
	.a(n250202));
   in01f01 FE_OFC20_n249394 (.o(FE_OFN20_n249394),
	.a(FE_OFN19_n249394));
   in01f01 FE_OFC19_n249394 (.o(FE_OFN19_n249394),
	.a(n249394));
   in01f10 FE_OFC18_n247494 (.o(FE_OFN18_n247494),
	.a(FE_OFN17_n247494));
   in01f04 FE_OFC17_n247494 (.o(FE_OFN17_n247494),
	.a(n247494));
   in01f08 FE_OFC16_n247350 (.o(FE_OFN16_n247350),
	.a(FE_OFN15_n247350));
   in01f02 FE_OFC15_n247350 (.o(FE_OFN15_n247350),
	.a(n247350));
   in01f06 FE_OFC14_n247150 (.o(FE_OFN14_n247150),
	.a(FE_OFN13_n247150));
   in01f02 FE_OFC13_n247150 (.o(FE_OFN13_n247150),
	.a(n247150));
   in01f01 FE_OFC8_n247076 (.o(FE_OFN8_n247076),
	.a(FE_OFN7_n247076));
   in01f01 FE_OFC7_n247076 (.o(FE_OFN7_n247076),
	.a(n247076));
   in01f06 FE_OFC6_n246618 (.o(FE_OFN6_n246618),
	.a(FE_OFN5_n246618));
   in01f01 FE_OFC5_n246618 (.o(FE_OFN5_n246618),
	.a(n246618));
   in01f08 FE_OFC4_n245443 (.o(FE_OFN4_n245443),
	.a(FE_OFN3_n245443));
   in01f01 FE_OFC3_n245443 (.o(FE_OFN3_n245443),
	.a(n245443));
   in01f06 FE_OFC2_g_swrst_r_n (.o(FE_OFN2_g_swrst_r_n),
	.a(FE_OFN1_g_swrst_r_n));
   in01f01 FE_OFC1_g_swrst_r_n (.o(FE_OFN1_g_swrst_r_n),
	.a(g_swrst_r_n));
   in01f02 FE_DBTC0_vmem_we_1_ (.o(vmem_we_n[1]),
	.a(vmem_we[1]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_0_ (.o(y1_bs_data_r[0]),
	.ck(clk),
	.d(y1_bs_data[0]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_1_ (.o(y1_bs_data_r[1]),
	.ck(clk),
	.d(y1_bs_data[1]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_2_ (.o(y1_bs_data_r[2]),
	.ck(clk),
	.d(y1_bs_data[2]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_3_ (.o(y1_bs_data_r[3]),
	.ck(clk),
	.d(y1_bs_data[3]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_4_ (.o(y1_bs_data_r[4]),
	.ck(clk),
	.d(y1_bs_data[4]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_5_ (.o(y1_bs_data_r[5]),
	.ck(clk),
	.d(y1_bs_data[5]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_6_ (.o(y1_bs_data_r[6]),
	.ck(clk),
	.d(y1_bs_data[6]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_7_ (.o(y1_bs_data_r[7]),
	.ck(clk),
	.d(y1_bs_data[7]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_8_ (.o(y1_bs_data_r[8]),
	.ck(clk),
	.d(y1_bs_data[8]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_9_ (.o(y1_bs_data_r[9]),
	.ck(clk),
	.d(y1_bs_data[9]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_10_ (.o(y1_bs_data_r[10]),
	.ck(clk),
	.d(y1_bs_data[10]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_11_ (.o(y1_bs_data_r[11]),
	.ck(clk),
	.d(y1_bs_data[11]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_12_ (.o(y1_bs_data_r[12]),
	.ck(clk),
	.d(y1_bs_data[12]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_13_ (.o(y1_bs_data_r[13]),
	.ck(clk),
	.d(y1_bs_data[13]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_14_ (.o(y1_bs_data_r[14]),
	.ck(clk),
	.d(y1_bs_data[14]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_15_ (.o(y1_bs_data_r[15]),
	.ck(clk),
	.d(y1_bs_data[15]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_16_ (.o(y1_bs_data_r[16]),
	.ck(clk),
	.d(y1_bs_data[16]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_17_ (.o(y1_bs_data_r[17]),
	.ck(clk),
	.d(y1_bs_data[17]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_18_ (.o(y1_bs_data_r[18]),
	.ck(clk),
	.d(y1_bs_data[18]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_19_ (.o(y1_bs_data_r[19]),
	.ck(clk),
	.d(y1_bs_data[19]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_20_ (.o(y1_bs_data_r[20]),
	.ck(clk),
	.d(y1_bs_data[20]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_21_ (.o(y1_bs_data_r[21]),
	.ck(clk),
	.d(y1_bs_data[21]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_22_ (.o(y1_bs_data_r[22]),
	.ck(clk),
	.d(y1_bs_data[22]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_23_ (.o(y1_bs_data_r[23]),
	.ck(clk),
	.d(y1_bs_data[23]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_24_ (.o(y1_bs_data_r[24]),
	.ck(clk),
	.d(y1_bs_data[24]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_25_ (.o(y1_bs_data_r[25]),
	.ck(clk),
	.d(y1_bs_data[25]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_26_ (.o(y1_bs_data_r[26]),
	.ck(clk),
	.d(y1_bs_data[26]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_27_ (.o(y1_bs_data_r[27]),
	.ck(clk),
	.d(y1_bs_data[27]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_28_ (.o(y1_bs_data_r[28]),
	.ck(clk),
	.d(y1_bs_data[28]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_29_ (.o(y1_bs_data_r[29]),
	.ck(clk),
	.d(y1_bs_data[29]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_30_ (.o(y1_bs_data_r[30]),
	.ck(clk),
	.d(y1_bs_data[30]));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_y1_bs_data_r_reg_31_ (.o(y1_bs_data_r[31]),
	.ck(clk),
	.d(y1_bs_data[31]));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_10_ (.o(busrtop_b_rreq_N295),
	.ck(clk),
	.d(busrtop_b_rreq_N85));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_11_ (.o(busrtop_b_rreq_N296),
	.ck(clk),
	.d(busrtop_b_rreq_N86));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_12_ (.o(busrtop_b_rreq_N229),
	.ck(clk),
	.d(busrtop_b_rreq_N87));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_13_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[13]),
	.ck(clk),
	.d(busrtop_b_rreq_N88));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_14_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[14]),
	.ck(clk),
	.d(busrtop_b_rreq_N89));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_15_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[15]),
	.ck(clk),
	.d(busrtop_b_rreq_N90));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_16_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[16]),
	.ck(clk),
	.d(busrtop_b_rreq_N91));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_17_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[17]),
	.ck(clk),
	.d(busrtop_b_rreq_N92));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_18_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[18]),
	.ck(clk),
	.d(busrtop_b_rreq_N93));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_19_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[19]),
	.ck(clk),
	.d(busrtop_b_rreq_N94));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_20_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[20]),
	.ck(clk),
	.d(busrtop_b_rreq_N95));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_21_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[21]),
	.ck(clk),
	.d(busrtop_b_rreq_N96));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_22_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[22]),
	.ck(clk),
	.d(busrtop_b_rreq_N97));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_23_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[23]),
	.ck(clk),
	.d(busrtop_b_rreq_N98));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_24_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[24]),
	.ck(clk),
	.d(busrtop_b_rreq_N99));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_25_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[25]),
	.ck(clk),
	.d(busrtop_b_rreq_N100));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_26_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[26]),
	.ck(clk),
	.d(busrtop_b_rreq_N101));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_27_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[27]),
	.ck(clk),
	.d(busrtop_b_rreq_N102));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_28_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[28]),
	.ck(clk),
	.d(busrtop_b_rreq_N103));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_29_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[29]),
	.ck(clk),
	.d(busrtop_b_rreq_N104));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_30_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[30]),
	.ck(clk),
	.d(busrtop_b_rreq_N105));
   ms00f80 busrtop_b_rreq_vrh_rrq_fldstatadd_r_reg_31_ (.o(busrtop_b_rreq_vrh_rrq_fldstatadd_r[31]),
	.ck(clk),
	.d(busrtop_b_rreq_N106));
   ms00f80 regtop_g_mem_rd_r_reg_0_ (.o(regtop_g_mem_rd_r[0]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[0]));
   ms00f80 regtop_g_mem_rd_r_reg_1_ (.o(regtop_g_mem_rd_r[1]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[1]));
   ms00f80 regtop_g_mem_rd_r_reg_2_ (.o(regtop_g_mem_rd_r[2]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[2]));
   ms00f80 regtop_g_mem_rd_r_reg_3_ (.o(regtop_g_mem_rd_r[3]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[3]));
   ms00f80 regtop_g_mem_rd_r_reg_4_ (.o(regtop_g_mem_rd_r[4]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[4]));
   ms00f80 regtop_g_mem_rd_r_reg_5_ (.o(regtop_g_mem_rd_r[5]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[5]));
   ms00f80 regtop_g_mem_rd_r_reg_6_ (.o(regtop_g_mem_rd_r[6]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[6]));
   ms00f80 regtop_g_mem_rd_r_reg_7_ (.o(regtop_g_mem_rd_r[7]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[7]));
   ms00f80 regtop_g_mem_rd_r_reg_8_ (.o(regtop_g_mem_rd_r[8]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[8]));
   ms00f80 regtop_g_mem_rd_r_reg_9_ (.o(regtop_g_mem_rd_r[9]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[9]));
   ms00f80 regtop_g_mem_rd_r_reg_10_ (.o(regtop_g_mem_rd_r[10]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[10]));
   ms00f80 regtop_g_mem_rd_r_reg_11_ (.o(regtop_g_mem_rd_r[11]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[11]));
   ms00f80 regtop_g_mem_rd_r_reg_12_ (.o(regtop_g_mem_rd_r[12]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[12]));
   ms00f80 regtop_g_mem_rd_r_reg_13_ (.o(regtop_g_mem_rd_r[13]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[13]));
   ms00f80 regtop_g_mem_rd_r_reg_14_ (.o(regtop_g_mem_rd_r[14]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[14]));
   ms00f80 regtop_g_mem_rd_r_reg_15_ (.o(regtop_g_mem_rd_r[15]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[15]));
   ms00f80 regtop_g_mem_rd_r_reg_16_ (.o(regtop_g_mem_rd_r[16]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[16]));
   ms00f80 regtop_g_mem_rd_r_reg_17_ (.o(regtop_g_mem_rd_r[17]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[17]));
   ms00f80 regtop_g_mem_rd_r_reg_18_ (.o(regtop_g_mem_rd_r[18]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[18]));
   ms00f80 regtop_g_mem_rd_r_reg_19_ (.o(regtop_g_mem_rd_r[19]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[19]));
   ms00f80 regtop_g_mem_rd_r_reg_20_ (.o(regtop_g_mem_rd_r[20]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[20]));
   ms00f80 regtop_g_mem_rd_r_reg_21_ (.o(regtop_g_mem_rd_r[21]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[21]));
   ms00f80 regtop_g_mem_rd_r_reg_22_ (.o(regtop_g_mem_rd_r[22]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[22]));
   ms00f80 regtop_g_mem_rd_r_reg_23_ (.o(regtop_g_mem_rd_r[23]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[23]));
   ms00f80 regtop_g_mem_rd_r_reg_24_ (.o(regtop_g_mem_rd_r[24]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[24]));
   ms00f80 regtop_g_mem_rd_r_reg_25_ (.o(regtop_g_mem_rd_r[25]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[25]));
   ms00f80 regtop_g_mem_rd_r_reg_26_ (.o(regtop_g_mem_rd_r[26]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[26]));
   ms00f80 regtop_g_mem_rd_r_reg_27_ (.o(regtop_g_mem_rd_r[27]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[27]));
   ms00f80 regtop_g_mem_rd_r_reg_28_ (.o(regtop_g_mem_rd_r[28]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[28]));
   ms00f80 regtop_g_mem_rd_r_reg_29_ (.o(regtop_g_mem_rd_r[29]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[29]));
   ms00f80 regtop_g_mem_rd_r_reg_30_ (.o(regtop_g_mem_rd_r[30]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[30]));
   ms00f80 regtop_g_mem_rd_r_reg_31_ (.o(regtop_g_mem_rd_r[31]),
	.ck(clk),
	.d(regtop_w1_hdi00_q[31]));
   ms00f80 regtop_g_dacksh_r_n_reg (.o(regtop_g_dacksh_r_n),
	.ck(clk),
	.d(sc_dmaack8_n));
   ms00f80 regtop_g_dack32_r_n_reg (.o(regtop_g_dack32_r_n),
	.ck(clk),
	.d(mr_dmaack8_n));
   ms00f80 regtop_g_wd_r_reg_0_ (.o(regtop_g_wd_r[0]),
	.ck(clk),
	.d(wbb_dat_i[0]));
   ms00f80 regtop_g_wd_r_reg_1_ (.o(regtop_g_wd_r[1]),
	.ck(clk),
	.d(wbb_dat_i[1]));
   ms00f80 regtop_g_wd_r_reg_2_ (.o(regtop_g_wd_r[2]),
	.ck(clk),
	.d(wbb_dat_i[2]));
   ms00f80 regtop_g_wd_r_reg_3_ (.o(regtop_g_wd_r[3]),
	.ck(clk),
	.d(wbb_dat_i[3]));
   ms00f80 regtop_g_wd_r_reg_4_ (.o(regtop_g_wd_r[4]),
	.ck(clk),
	.d(wbb_dat_i[4]));
   ms00f80 regtop_g_wd_r_reg_5_ (.o(regtop_g_wd_r[5]),
	.ck(clk),
	.d(wbb_dat_i[5]));
   ms00f80 regtop_g_wd_r_reg_6_ (.o(regtop_g_wd_r[6]),
	.ck(clk),
	.d(wbb_dat_i[6]));
   ms00f80 regtop_g_wd_r_reg_7_ (.o(regtop_g_wd_r[7]),
	.ck(clk),
	.d(wbb_dat_i[7]));
   ms00f80 regtop_g_wd_r_reg_8_ (.o(regtop_g_wd_r[8]),
	.ck(clk),
	.d(wbb_dat_i[8]));
   ms00f80 regtop_g_wd_r_reg_9_ (.o(regtop_g_wd_r[9]),
	.ck(clk),
	.d(wbb_dat_i[9]));
   ms00f80 regtop_g_wd_r_reg_10_ (.o(regtop_g_wd_r[10]),
	.ck(clk),
	.d(wbb_dat_i[10]));
   ms00f80 regtop_g_wd_r_reg_11_ (.o(regtop_g_wd_r[11]),
	.ck(clk),
	.d(wbb_dat_i[11]));
   ms00f80 regtop_g_wd_r_reg_12_ (.o(regtop_g_wd_r[12]),
	.ck(clk),
	.d(wbb_dat_i[12]));
   ms00f80 regtop_g_wd_r_reg_13_ (.o(regtop_g_wd_r[13]),
	.ck(clk),
	.d(wbb_dat_i[13]));
   ms00f80 regtop_g_wd_r_reg_14_ (.o(regtop_g_wd_r[14]),
	.ck(clk),
	.d(wbb_dat_i[14]));
   ms00f80 regtop_g_wd_r_reg_15_ (.o(regtop_g_wd_r[15]),
	.ck(clk),
	.d(wbb_dat_i[15]));
   ms00f80 regtop_g_wd_r_reg_16_ (.o(regtop_g_wd_r[16]),
	.ck(clk),
	.d(wbb_dat_i[16]));
   ms00f80 regtop_g_wd_r_reg_17_ (.o(regtop_g_wd_r[17]),
	.ck(clk),
	.d(wbb_dat_i[17]));
   ms00f80 regtop_g_wd_r_reg_18_ (.o(regtop_g_wd_r[18]),
	.ck(clk),
	.d(wbb_dat_i[18]));
   ms00f80 regtop_g_wd_r_reg_19_ (.o(regtop_g_wd_r[19]),
	.ck(clk),
	.d(wbb_dat_i[19]));
   ms00f80 regtop_g_wd_r_reg_20_ (.o(regtop_g_wd_r[20]),
	.ck(clk),
	.d(wbb_dat_i[20]));
   ms00f80 regtop_g_wd_r_reg_21_ (.o(regtop_g_wd_r[21]),
	.ck(clk),
	.d(wbb_dat_i[21]));
   ms00f80 regtop_g_wd_r_reg_22_ (.o(regtop_g_wd_r[22]),
	.ck(clk),
	.d(wbb_dat_i[22]));
   ms00f80 regtop_g_wd_r_reg_23_ (.o(regtop_g_wd_r[23]),
	.ck(clk),
	.d(wbb_dat_i[23]));
   ms00f80 regtop_g_wd_r_reg_24_ (.o(regtop_g_wd_r[24]),
	.ck(clk),
	.d(wbb_dat_i[24]));
   ms00f80 regtop_g_wd_r_reg_25_ (.o(regtop_g_wd_r[25]),
	.ck(clk),
	.d(wbb_dat_i[25]));
   ms00f80 regtop_g_wd_r_reg_26_ (.o(regtop_g_wd_r[26]),
	.ck(clk),
	.d(wbb_dat_i[26]));
   ms00f80 regtop_g_wd_r_reg_27_ (.o(regtop_g_wd_r[27]),
	.ck(clk),
	.d(wbb_dat_i[27]));
   ms00f80 regtop_g_wd_r_reg_28_ (.o(regtop_g_wd_r[28]),
	.ck(clk),
	.d(wbb_dat_i[28]));
   ms00f80 regtop_g_wd_r_reg_29_ (.o(regtop_g_wd_r[29]),
	.ck(clk),
	.d(wbb_dat_i[29]));
   ms00f80 regtop_g_wd_r_reg_30_ (.o(regtop_g_wd_r[30]),
	.ck(clk),
	.d(wbb_dat_i[30]));
   ms00f80 regtop_g_wd_r_reg_31_ (.o(regtop_g_wd_r[31]),
	.ck(clk),
	.d(wbb_dat_i[31]));
   ms00f80 regtop_g_a_r_reg_2_ (.o(regtop_g_a_r[2]),
	.ck(clk),
	.d(wbb_adr_i[2]));
   ms00f80 regtop_g_a_r_reg_3_ (.o(regtop_g_a_r[3]),
	.ck(clk),
	.d(wbb_adr_i[3]));
   ms00f80 regtop_g_a_r_reg_4_ (.o(regtop_g_a_r[4]),
	.ck(clk),
	.d(wbb_adr_i[4]));
   ms00f80 regtop_g_a_r_reg_5_ (.o(regtop_g_a_r[5]),
	.ck(clk),
	.d(wbb_adr_i[5]));
   ms00f80 regtop_g_a_r_reg_6_ (.o(regtop_g_a_r[6]),
	.ck(clk),
	.d(wbb_adr_i[6]));
   ms00f80 regtop_g_a_r_reg_7_ (.o(regtop_g_a_r[7]),
	.ck(clk),
	.d(wbb_adr_i[7]));
   ms00f80 regtop_g_a_r_reg_8_ (.o(regtop_g_a_r[8]),
	.ck(clk),
	.d(wbb_adr_i[8]));
   ms00f80 regtop_g_write_r_n_reg (.o(regtop_g_write_r_n),
	.ck(clk),
	.d(n243097));
   ms00f80 regtop_g_read_r_n_reg (.o(regtop_g_read_r_n),
	.ck(clk),
	.d(wbb_we_i));
   ms00f80 regtop_g_ms_r_n_reg (.o(regtop_g_ms_r_n),
	.ck(clk),
	.d(n243096));
   ms00f80 regtop_g_line_offset_r_reg (.o(g_line_offset_r),
	.ck(clk),
	.d(n212788));
   ms00f80 regtop_g_cbcr_offset_r_reg_0_ (.o(g_cbcr_offset_r[0]),
	.ck(clk),
	.d(n212787));
   ms00f80 regtop_g_cbcr_offset_r_reg_11_ (.o(g_cbcr_offset_r[11]),
	.ck(clk),
	.d(n212786));
   ms00f80 regtop_g_cbcr_offset_r_reg_10_ (.o(g_cbcr_offset_r[10]),
	.ck(clk),
	.d(n212785));
   ms00f80 regtop_g_cbcr_offset_r_reg_9_ (.o(g_cbcr_offset_r[9]),
	.ck(clk),
	.d(n212784));
   ms00f80 regtop_g_cbcr_offset_r_reg_8_ (.o(g_cbcr_offset_r[8]),
	.ck(clk),
	.d(n212783));
   ms00f80 regtop_g_cbcr_offset_r_reg_7_ (.o(g_cbcr_offset_r[7]),
	.ck(clk),
	.d(n212782));
   ms00f80 regtop_g_cbcr_offset_r_reg_6_ (.o(g_cbcr_offset_r[6]),
	.ck(clk),
	.d(n212781));
   ms00f80 regtop_g_cbcr_offset_r_reg_5_ (.o(g_cbcr_offset_r[5]),
	.ck(clk),
	.d(n212780));
   ms00f80 regtop_g_cbcr_offset_r_reg_4_ (.o(g_cbcr_offset_r[4]),
	.ck(clk),
	.d(n212779));
   ms00f80 regtop_g_cbcr_offset_r_reg_3_ (.o(g_cbcr_offset_r[3]),
	.ck(clk),
	.d(n212778));
   ms00f80 regtop_g_cbcr_offset_r_reg_2_ (.o(g_cbcr_offset_r[2]),
	.ck(clk),
	.d(n212777));
   ms00f80 regtop_g_cbcr_offset_r_reg_1_ (.o(g_cbcr_offset_r[1]),
	.ck(clk),
	.d(n212776));
   ms00f80 regtop_g_field_offset_r_reg_0_ (.o(g_field_offset_r[0]),
	.ck(clk),
	.d(n212775));
   ms00f80 regtop_g_field_offset_r_reg_11_ (.o(g_field_offset_r[11]),
	.ck(clk),
	.d(n212774));
   ms00f80 regtop_g_field_offset_r_reg_10_ (.o(g_field_offset_r[10]),
	.ck(clk),
	.d(n212773));
   ms00f80 regtop_g_field_offset_r_reg_9_ (.o(g_field_offset_r[9]),
	.ck(clk),
	.d(n212772));
   ms00f80 regtop_g_field_offset_r_reg_8_ (.o(g_field_offset_r[8]),
	.ck(clk),
	.d(n212771));
   ms00f80 regtop_g_field_offset_r_reg_7_ (.o(g_field_offset_r[7]),
	.ck(clk),
	.d(n212770));
   ms00f80 regtop_g_field_offset_r_reg_6_ (.o(g_field_offset_r[6]),
	.ck(clk),
	.d(n212769));
   ms00f80 regtop_g_field_offset_r_reg_5_ (.o(g_field_offset_r[5]),
	.ck(clk),
	.d(n212768));
   ms00f80 regtop_g_field_offset_r_reg_4_ (.o(g_field_offset_r[4]),
	.ck(clk),
	.d(n212767));
   ms00f80 regtop_g_field_offset_r_reg_3_ (.o(g_field_offset_r[3]),
	.ck(clk),
	.d(n212766));
   ms00f80 regtop_g_field_offset_r_reg_2_ (.o(g_field_offset_r[2]),
	.ck(clk),
	.d(n212765));
   ms00f80 regtop_g_field_offset_r_reg_1_ (.o(g_field_offset_r[1]),
	.ck(clk),
	.d(n212764));
   ms00f80 regtop_g_field_start_add_r_reg_10_ (.o(g_field_start_add_r[10]),
	.ck(clk),
	.d(n212763));
   ms00f80 regtop_g_field_start_add_r_reg_31_ (.o(g_field_start_add_r[31]),
	.ck(clk),
	.d(n212762));
   ms00f80 regtop_g_field_start_add_r_reg_30_ (.o(g_field_start_add_r[30]),
	.ck(clk),
	.d(n212761));
   ms00f80 regtop_g_field_start_add_r_reg_29_ (.o(g_field_start_add_r[29]),
	.ck(clk),
	.d(n212760));
   ms00f80 regtop_g_field_start_add_r_reg_28_ (.o(g_field_start_add_r[28]),
	.ck(clk),
	.d(n212759));
   ms00f80 regtop_g_field_start_add_r_reg_27_ (.o(g_field_start_add_r[27]),
	.ck(clk),
	.d(n212758));
   ms00f80 regtop_g_field_start_add_r_reg_26_ (.o(g_field_start_add_r[26]),
	.ck(clk),
	.d(n212757));
   ms00f80 regtop_g_field_start_add_r_reg_25_ (.o(g_field_start_add_r[25]),
	.ck(clk),
	.d(n212756));
   ms00f80 regtop_g_field_start_add_r_reg_24_ (.o(g_field_start_add_r[24]),
	.ck(clk),
	.d(n212755));
   ms00f80 regtop_g_field_start_add_r_reg_23_ (.o(g_field_start_add_r[23]),
	.ck(clk),
	.d(n212754));
   ms00f80 regtop_g_field_start_add_r_reg_22_ (.o(g_field_start_add_r[22]),
	.ck(clk),
	.d(n212753));
   ms00f80 regtop_g_field_start_add_r_reg_21_ (.o(g_field_start_add_r[21]),
	.ck(clk),
	.d(n212752));
   ms00f80 regtop_g_field_start_add_r_reg_20_ (.o(g_field_start_add_r[20]),
	.ck(clk),
	.d(n212751));
   ms00f80 regtop_g_field_start_add_r_reg_19_ (.o(g_field_start_add_r[19]),
	.ck(clk),
	.d(n212750));
   ms00f80 regtop_g_field_start_add_r_reg_18_ (.o(g_field_start_add_r[18]),
	.ck(clk),
	.d(n212749));
   ms00f80 regtop_g_field_start_add_r_reg_17_ (.o(g_field_start_add_r[17]),
	.ck(clk),
	.d(n212748));
   ms00f80 regtop_g_field_start_add_r_reg_16_ (.o(g_field_start_add_r[16]),
	.ck(clk),
	.d(n212747));
   ms00f80 regtop_g_field_start_add_r_reg_15_ (.o(g_field_start_add_r[15]),
	.ck(clk),
	.d(n212746));
   ms00f80 regtop_g_field_start_add_r_reg_14_ (.o(g_field_start_add_r[14]),
	.ck(clk),
	.d(n212745));
   ms00f80 regtop_g_field_start_add_r_reg_13_ (.o(g_field_start_add_r[13]),
	.ck(clk),
	.d(n212744));
   ms00f80 regtop_g_field_start_add_r_reg_12_ (.o(g_field_start_add_r[12]),
	.ck(clk),
	.d(n212743));
   ms00f80 regtop_g_field_start_add_r_reg_11_ (.o(g_field_start_add_r[11]),
	.ck(clk),
	.d(n212742));
   ms00f80 regtop_g_icdc_r_reg (.o(regtop_g_icdc_r),
	.ck(clk),
	.d(n212741));
   ms00f80 regtop_g_icsh_r_reg (.o(regtop_g_icsh_r),
	.ck(clk),
	.d(n212740));
   ms00f80 regtop_g_icph_r_reg (.o(regtop_g_icph_r),
	.ck(clk),
	.d(n212739));
   ms00f80 regtop_g_icpi_r_reg (.o(regtop_g_icpi_r),
	.ck(clk),
	.d(n212738));
   ms00f80 regtop_g_icnf_r_reg (.o(regtop_g_icnf_r),
	.ck(clk),
	.d(n212737));
   ms00f80 regtop_g_icfb_r_reg (.o(regtop_g_icfb_r),
	.ck(clk),
	.d(n212736));
   ms00f80 regtop_g_icfp_r_reg (.o(regtop_g_icfp_r),
	.ck(clk),
	.d(n212735));
   ms00f80 regtop_g_icsr_r_reg (.o(regtop_g_icsr_r),
	.ck(clk),
	.d(n212734));
   ms00f80 regtop_g_icsw_r_reg (.o(regtop_g_icsw_r),
	.ck(clk),
	.d(n212733));
   ms00f80 regtop_g_icuc_r_reg (.o(regtop_g_icuc_r),
	.ck(clk),
	.d(n212732));
   ms00f80 regtop_g_amod_r_reg (.o(g_vldmode_r[0]),
	.ck(clk),
	.d(n212731));
   ms00f80 regtop_g_imod_r_reg (.o(regtop_g_imod_r),
	.ck(clk),
	.d(n212730));
   ms00f80 regtop_g_bmod_r_reg (.o(g_bmod_r),
	.ck(clk),
	.d(n212729));
   ms00f80 regtop_g_dmod_r_reg (.o(regtop_g_dmod_r),
	.ck(clk),
	.d(n212728));
   ms00f80 regtop_g_pmod_r_reg (.o(g_pmod_r),
	.ck(clk),
	.d(n212727));
   ms00f80 regtop_g_mmod_r_reg (.o(g_vldmode_r[1]),
	.ck(clk),
	.d(n212726));
   ms00f80 regtop_g_fcyc_en_r_reg (.o(g_fcyc_en_r),
	.ck(clk),
	.d(n212725));
   ms00f80 regtop_g_fcyc_r_reg_1_ (.o(g_fcyc_r[1]),
	.ck(clk),
	.d(n212724));
   ms00f80 regtop_g_fcyc_r_reg_2_ (.o(g_fcyc_r[2]),
	.ck(clk),
	.d(n212723));
   ms00f80 regtop_g_fcyc_r_reg_3_ (.o(g_fcyc_r[3]),
	.ck(clk),
	.d(n212722));
   ms00f80 regtop_g_fcyc_r_reg_4_ (.o(g_fcyc_r[4]),
	.ck(clk),
	.d(n212721));
   ms00f80 regtop_g_fcyc_r_reg_5_ (.o(g_fcyc_r[5]),
	.ck(clk),
	.d(n212720));
   ms00f80 regtop_g_fcyc_r_reg_6_ (.o(g_fcyc_r[6]),
	.ck(clk),
	.d(n212719));
   ms00f80 regtop_g_fcyc_r_reg_7_ (.o(g_fcyc_r[7]),
	.ck(clk),
	.d(n212718));
   ms00f80 regtop_g_fcyc_r_reg_8_ (.o(g_fcyc_r[8]),
	.ck(clk),
	.d(n212717));
   ms00f80 regtop_g_fcyc_r_reg_9_ (.o(g_fcyc_r[9]),
	.ck(clk),
	.d(n212716));
   ms00f80 regtop_g_fcyc_r_reg_10_ (.o(g_fcyc_r[10]),
	.ck(clk),
	.d(n212715));
   ms00f80 regtop_g_fcyc_r_reg_11_ (.o(g_fcyc_r[11]),
	.ck(clk),
	.d(n212714));
   ms00f80 regtop_g_fcyc_r_reg_12_ (.o(g_fcyc_r[12]),
	.ck(clk),
	.d(n212713));
   ms00f80 regtop_g_fcyc_r_reg_13_ (.o(g_fcyc_r[13]),
	.ck(clk),
	.d(n212712));
   ms00f80 regtop_g_fcyc_r_reg_14_ (.o(g_fcyc_r[14]),
	.ck(clk),
	.d(n212711));
   ms00f80 regtop_g_fcyc_r_reg_15_ (.o(g_fcyc_r[15]),
	.ck(clk),
	.d(n212710));
   ms00f80 regtop_g_fcyc_r_reg_16_ (.o(g_fcyc_r[16]),
	.ck(clk),
	.d(n212709));
   ms00f80 regtop_g_fcyc_r_reg_17_ (.o(g_fcyc_r[17]),
	.ck(clk),
	.d(n212708));
   ms00f80 regtop_g_fcyc_r_reg_0_ (.o(g_fcyc_r[0]),
	.ck(clk),
	.d(n212707));
   ms00f80 regtop_g_pcut_r_reg_0_ (.o(g_pcut_r[0]),
	.ck(clk),
	.d(n212706));
   ms00f80 regtop_g_pcut_r_reg_11_ (.o(g_pcut_r[11]),
	.ck(clk),
	.d(n212705));
   ms00f80 regtop_g_pcut_r_reg_10_ (.o(g_pcut_r[10]),
	.ck(clk),
	.d(n212704));
   ms00f80 regtop_g_pcut_r_reg_9_ (.o(g_pcut_r[9]),
	.ck(clk),
	.d(n212703));
   ms00f80 regtop_g_pcut_r_reg_8_ (.o(g_pcut_r[8]),
	.ck(clk),
	.d(n212702));
   ms00f80 regtop_g_pcut_r_reg_7_ (.o(g_pcut_r[7]),
	.ck(clk),
	.d(n212701));
   ms00f80 regtop_g_pcut_r_reg_6_ (.o(g_pcut_r[6]),
	.ck(clk),
	.d(n212700));
   ms00f80 regtop_g_pcut_r_reg_5_ (.o(g_pcut_r[5]),
	.ck(clk),
	.d(n212699));
   ms00f80 regtop_g_pcut_r_reg_4_ (.o(g_pcut_r[4]),
	.ck(clk),
	.d(n212698));
   ms00f80 regtop_g_pcut_r_reg_3_ (.o(g_pcut_r[3]),
	.ck(clk),
	.d(n212697));
   ms00f80 regtop_g_pcut_r_reg_2_ (.o(g_pcut_r[2]),
	.ck(clk),
	.d(n212696));
   ms00f80 regtop_g_pcut_r_reg_1_ (.o(g_pcut_r[1]),
	.ck(clk),
	.d(n212695));
   ms00f80 regtop_g_mbc_en_r_reg (.o(g_mbc_en_r),
	.ck(clk),
	.d(n212694));
   ms00f80 regtop_g_mbc_r_reg_1_ (.o(g_mbc_r[1]),
	.ck(clk),
	.d(n212693));
   ms00f80 regtop_g_mbc_r_reg_2_ (.o(g_mbc_r[2]),
	.ck(clk),
	.d(n212692));
   ms00f80 regtop_g_mbc_r_reg_3_ (.o(g_mbc_r[3]),
	.ck(clk),
	.d(n212691));
   ms00f80 regtop_g_mbc_r_reg_4_ (.o(g_mbc_r[4]),
	.ck(clk),
	.d(n212690));
   ms00f80 regtop_g_mbc_r_reg_5_ (.o(g_mbc_r[5]),
	.ck(clk),
	.d(n212689));
   ms00f80 regtop_g_mbc_r_reg_6_ (.o(g_mbc_r[6]),
	.ck(clk),
	.d(n212688));
   ms00f80 regtop_g_mbc_r_reg_7_ (.o(g_mbc_r[7]),
	.ck(clk),
	.d(n212687));
   ms00f80 regtop_g_mbc_r_reg_8_ (.o(g_mbc_r[8]),
	.ck(clk),
	.d(n212686));
   ms00f80 regtop_g_mbc_r_reg_9_ (.o(g_mbc_r[9]),
	.ck(clk),
	.d(n212685));
   ms00f80 regtop_g_mbc_r_reg_10_ (.o(g_mbc_r[10]),
	.ck(clk),
	.d(n212684));
   ms00f80 regtop_g_mbc_r_reg_11_ (.o(g_mbc_r[11]),
	.ck(clk),
	.d(n212683));
   ms00f80 regtop_g_mbc_r_reg_0_ (.o(g_mbc_r[0]),
	.ck(clk),
	.d(n212682));
   ms00f80 regtop_g_init_cnt_r_reg_1_ (.o(regtop_g_init_cnt_r[1]),
	.ck(clk),
	.d(n245109));
   ms00f80 regtop_g_init_cnt_r_reg_2_ (.o(regtop_g_init_cnt_r[2]),
	.ck(clk),
	.d(n245110));
   ms00f80 regtop_g_init_vld_r_s_reg (.o(g_init_vld_r_s),
	.ck(clk),
	.d(n212681));
   ms00f80 regtop_g_init_cnt_r_reg_0_ (.o(regtop_g_init_cnt_r[0]),
	.ck(clk),
	.d(n245111));
   ms00f80 regtop_g_swrst_r_n_reg (.o(g_swrst_r_n),
	.ck(clk),
	.d(n212680));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_feed_on_reg (.o(vldtop_vld_syndec_vld_vlfeed_feed_on),
	.ck(clk),
	.d(n212679));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_v1_bs_req_n_reg (.o(v1_bs_req_n),
	.ck(clk),
	.d(n212678));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_dselect_r_reg (.o(vldtop_vld_syndec_vld_vlfeed_dselect_r),
	.ck(clk),
	.d(n212677));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_0_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[0]),
	.ck(clk),
	.d(n253070));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_1_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[1]),
	.ck(clk),
	.d(n253069));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_2_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[2]),
	.ck(clk),
	.d(n253068));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_3_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[3]),
	.ck(clk),
	.d(n253067));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_4_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[4]),
	.ck(clk),
	.d(n253066));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_5_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[5]),
	.ck(clk),
	.d(n253065));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_6_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[6]),
	.ck(clk),
	.d(n253064));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_7_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[7]),
	.ck(clk),
	.d(n253063));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_8_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[8]),
	.ck(clk),
	.d(n253062));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_9_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[9]),
	.ck(clk),
	.d(n253061));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_10_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[10]),
	.ck(clk),
	.d(n253060));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_11_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[11]),
	.ck(clk),
	.d(n253059));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_12_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[12]),
	.ck(clk),
	.d(n253058));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_13_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[13]),
	.ck(clk),
	.d(n253057));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_14_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[14]),
	.ck(clk),
	.d(n253056));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_15_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[15]),
	.ck(clk),
	.d(n253055));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_16_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[16]),
	.ck(clk),
	.d(n253054));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_17_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[17]),
	.ck(clk),
	.d(n253053));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_18_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[18]),
	.ck(clk),
	.d(n253052));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_19_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[19]),
	.ck(clk),
	.d(n253051));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_20_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[20]),
	.ck(clk),
	.d(n253050));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_21_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[21]),
	.ck(clk),
	.d(n253049));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_22_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[22]),
	.ck(clk),
	.d(n253048));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_23_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[23]),
	.ck(clk),
	.d(n253047));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_24_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[24]),
	.ck(clk),
	.d(n253046));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_25_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[25]),
	.ck(clk),
	.d(n253045));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_26_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[26]),
	.ck(clk),
	.d(n253044));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_27_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[27]),
	.ck(clk),
	.d(n253043));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_28_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[28]),
	.ck(clk),
	.d(n253042));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_29_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[29]),
	.ck(clk),
	.d(n253041));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_30_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[30]),
	.ck(clk),
	.d(n253040));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_temporal_reg_31_ (.o(vldtop_vld_syndec_vld_vlfeed_temporal[31]),
	.ck(clk),
	.d(n253039));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_0_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[0]),
	.ck(clk),
	.d(n212644));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_0_ (.o(vldtop_vld_syndec_UREG[0]),
	.ck(clk),
	.d(n253102));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_1_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[1]),
	.ck(clk),
	.d(n212642));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_1_ (.o(vldtop_vld_syndec_UREG[1]),
	.ck(clk),
	.d(n253101));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_2_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[2]),
	.ck(clk),
	.d(n212640));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_2_ (.o(vldtop_vld_syndec_UREG[2]),
	.ck(clk),
	.d(n253100));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_3_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[3]),
	.ck(clk),
	.d(n212638));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_3_ (.o(vldtop_vld_syndec_UREG[3]),
	.ck(clk),
	.d(n253099));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_4_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[4]),
	.ck(clk),
	.d(n212636));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_4_ (.o(vldtop_vld_syndec_UREG[4]),
	.ck(clk),
	.d(n253098));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_5_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[5]),
	.ck(clk),
	.d(n212634));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_5_ (.o(vldtop_vld_syndec_UREG[5]),
	.ck(clk),
	.d(n253097));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_6_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[6]),
	.ck(clk),
	.d(n212632));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_6_ (.o(vldtop_vld_syndec_UREG[6]),
	.ck(clk),
	.d(n253096));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_7_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[7]),
	.ck(clk),
	.d(n212630));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_7_ (.o(vldtop_vld_syndec_UREG[7]),
	.ck(clk),
	.d(n253095));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_8_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[8]),
	.ck(clk),
	.d(n212628));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_8_ (.o(vldtop_vld_syndec_UREG[8]),
	.ck(clk),
	.d(n253094));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_9_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[9]),
	.ck(clk),
	.d(n212626));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_9_ (.o(vldtop_vld_syndec_UREG[9]),
	.ck(clk),
	.d(n253093));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_10_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[10]),
	.ck(clk),
	.d(n212624));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_10_ (.o(vldtop_vld_syndec_UREG[10]),
	.ck(clk),
	.d(n253092));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_11_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[11]),
	.ck(clk),
	.d(n212622));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_11_ (.o(vldtop_vld_syndec_UREG[11]),
	.ck(clk),
	.d(n253091));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_12_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[12]),
	.ck(clk),
	.d(n212620));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_12_ (.o(vldtop_vld_syndec_UREG[12]),
	.ck(clk),
	.d(n253090));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_13_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[13]),
	.ck(clk),
	.d(n212618));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_13_ (.o(vldtop_vld_syndec_UREG[13]),
	.ck(clk),
	.d(n253089));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_14_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[14]),
	.ck(clk),
	.d(n212616));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_14_ (.o(vldtop_vld_syndec_UREG[14]),
	.ck(clk),
	.d(n253088));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_15_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[15]),
	.ck(clk),
	.d(n212614));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_15_ (.o(vldtop_vld_syndec_UREG[15]),
	.ck(clk),
	.d(n253087));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_16_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[16]),
	.ck(clk),
	.d(n212612));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_16_ (.o(vldtop_vld_syndec_UREG[16]),
	.ck(clk),
	.d(n253086));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_17_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[17]),
	.ck(clk),
	.d(n212610));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_17_ (.o(vldtop_vld_syndec_UREG[17]),
	.ck(clk),
	.d(n253085));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_18_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[18]),
	.ck(clk),
	.d(n212608));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_18_ (.o(vldtop_vld_syndec_UREG[18]),
	.ck(clk),
	.d(n253084));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_19_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[19]),
	.ck(clk),
	.d(n212606));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_19_ (.o(vldtop_vld_syndec_UREG[19]),
	.ck(clk),
	.d(n253083));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_20_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[20]),
	.ck(clk),
	.d(n212604));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_20_ (.o(vldtop_vld_syndec_UREG[20]),
	.ck(clk),
	.d(n253082));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_21_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[21]),
	.ck(clk),
	.d(n212602));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_21_ (.o(vldtop_vld_syndec_UREG[21]),
	.ck(clk),
	.d(n253081));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_22_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[22]),
	.ck(clk),
	.d(n212600));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_22_ (.o(vldtop_vld_syndec_UREG[22]),
	.ck(clk),
	.d(n253080));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_23_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[23]),
	.ck(clk),
	.d(n212598));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_23_ (.o(vldtop_vld_syndec_UREG[23]),
	.ck(clk),
	.d(n253079));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_24_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[24]),
	.ck(clk),
	.d(n212596));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_24_ (.o(vldtop_vld_syndec_UREG[24]),
	.ck(clk),
	.d(n253078));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_25_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[25]),
	.ck(clk),
	.d(n212594));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_25_ (.o(vldtop_vld_syndec_UREG[25]),
	.ck(clk),
	.d(n253077));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_26_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[26]),
	.ck(clk),
	.d(n212592));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_26_ (.o(vldtop_vld_syndec_UREG[26]),
	.ck(clk),
	.d(n253076));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_27_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[27]),
	.ck(clk),
	.d(n212590));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_27_ (.o(vldtop_vld_syndec_UREG[27]),
	.ck(clk),
	.d(n253075));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_28_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[28]),
	.ck(clk),
	.d(n212588));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_28_ (.o(vldtop_vld_syndec_UREG[28]),
	.ck(clk),
	.d(n253074));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_29_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[29]),
	.ck(clk),
	.d(n212586));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_29_ (.o(vldtop_vld_syndec_UREG[29]),
	.ck(clk),
	.d(n253073));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_30_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[30]),
	.ck(clk),
	.d(n212584));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_30_ (.o(vldtop_vld_syndec_UREG[30]),
	.ck(clk),
	.d(n253072));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_lower_reg_31_ (.o(vldtop_vld_syndec_vld_vlfeed_lower[31]),
	.ck(clk),
	.d(n212582));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_UREG_reg_31_ (.o(vldtop_vld_syndec_UREG[31]),
	.ck(clk),
	.d(n253071));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_ADP_reg_1_ (.o(vldtop_vld_syndec_ADP[1]),
	.ck(clk),
	.d(n212579));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_ADP_reg_2_ (.o(vldtop_vld_syndec_ADP[2]),
	.ck(clk),
	.d(n212578));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_ADP_reg_3_ (.o(vldtop_vld_syndec_ADP[3]),
	.ck(clk),
	.d(n212577));
   ms00f80 vldtop_vld_syndec_vld_vlfeed_ADP_reg_4_ (.o(vldtop_vld_syndec_ADP[4]),
	.ck(clk),
	.d(n212576));
   ms00f80 vldtop_vld_syndec_vld_vscdet_v_prezerotmp_r_reg_1_ (.o(vldtop_vld_syndec_vld_vscdet_v_prezerotmp_r[1]),
	.ck(clk),
	.d(n212574));
   ms00f80 vldtop_vld_syndec_vld_vscdet_v_prezerohld_r_reg_1_ (.o(vldtop_vld_syndec_vld_vscdet_v_prezerohld_r[1]),
	.ck(clk),
	.d(n212573));
   ms00f80 vldtop_vld_syndec_vld_vscdet_v_prezerotmp_r_reg_0_ (.o(vldtop_vld_syndec_vld_vscdet_v_prezerotmp_r[0]),
	.ck(clk),
	.d(n212572));
   ms00f80 vldtop_vld_syndec_vld_vscdet_v_prezerohld_r_reg_0_ (.o(vldtop_vld_syndec_vld_vscdet_v_prezerohld_r[0]),
	.ck(clk),
	.d(n212571));
   ms00f80 regtop_g_dcnt_r_reg (.o(regtop_g_dcnt_r),
	.ck(clk),
	.d(n212562));
   ms00f80 regtop_g_hsdc_r_reg_0_ (.o(g_hsdc_r[0]),
	.ck(clk),
	.d(n212561));
   ms00f80 regtop_g_hsdc_r_reg_6_ (.o(g_hsdc_r[6]),
	.ck(clk),
	.d(n212560));
   ms00f80 regtop_g_hsdc_r_reg_5_ (.o(g_hsdc_r[5]),
	.ck(clk),
	.d(n212559));
   ms00f80 regtop_g_hsdc_r_reg_4_ (.o(g_hsdc_r[4]),
	.ck(clk),
	.d(n212558));
   ms00f80 regtop_g_hsdc_r_reg_3_ (.o(g_hsdc_r[3]),
	.ck(clk),
	.d(n212557));
   ms00f80 regtop_g_hsdc_r_reg_2_ (.o(g_hsdc_r[2]),
	.ck(clk),
	.d(n212556));
   ms00f80 regtop_g_hsdc_r_reg_1_ (.o(g_hsdc_r[1]),
	.ck(clk),
	.d(n212555));
   ms00f80 regtop_g_vsdc_r_reg_1_ (.o(g_vsdc_r[1]),
	.ck(clk),
	.d(n212554));
   ms00f80 regtop_g_vsdc_r_reg_2_ (.o(g_vsdc_r[2]),
	.ck(clk),
	.d(n212553));
   ms00f80 regtop_g_vsdc_r_reg_3_ (.o(g_vsdc_r[3]),
	.ck(clk),
	.d(n212552));
   ms00f80 regtop_g_vsdc_r_reg_4_ (.o(g_vsdc_r[4]),
	.ck(clk),
	.d(n212551));
   ms00f80 regtop_g_vsdc_r_reg_5_ (.o(g_vsdc_r[5]),
	.ck(clk),
	.d(n212550));
   ms00f80 regtop_g_vsdc_r_reg_6_ (.o(g_vsdc_r[6]),
	.ck(clk),
	.d(n212549));
   ms00f80 regtop_g_vsdc_r_reg_0_ (.o(g_vsdc_r[0]),
	.ck(clk),
	.d(n212548));
   ms00f80 regtop_g_hs60p_r_reg_1_ (.o(g_hs60p_r[1]),
	.ck(clk),
	.d(n212547));
   ms00f80 regtop_g_hs60p_r_reg_2_ (.o(g_hs60p_r[2]),
	.ck(clk),
	.d(n212546));
   ms00f80 regtop_g_hs60p_r_reg_3_ (.o(g_hs60p_r[3]),
	.ck(clk),
	.d(n212545));
   ms00f80 regtop_g_hs60p_r_reg_4_ (.o(g_hs60p_r[4]),
	.ck(clk),
	.d(n212544));
   ms00f80 regtop_g_hs60p_r_reg_5_ (.o(g_hs60p_r[5]),
	.ck(clk),
	.d(n212543));
   ms00f80 regtop_g_hs60p_r_reg_6_ (.o(g_hs60p_r[6]),
	.ck(clk),
	.d(n212542));
   ms00f80 regtop_g_hs60p_r_reg_0_ (.o(g_hs60p_r[0]),
	.ck(clk),
	.d(n212541));
   ms00f80 regtop_g_vs60p_r_reg_1_ (.o(g_vs60p_r[1]),
	.ck(clk),
	.d(n212540));
   ms00f80 regtop_g_vs60p_r_reg_2_ (.o(g_vs60p_r[2]),
	.ck(clk),
	.d(n212539));
   ms00f80 regtop_g_vs60p_r_reg_3_ (.o(g_vs60p_r[3]),
	.ck(clk),
	.d(n212538));
   ms00f80 regtop_g_vs60p_r_reg_4_ (.o(g_vs60p_r[4]),
	.ck(clk),
	.d(n212537));
   ms00f80 regtop_g_vs60p_r_reg_5_ (.o(g_vs60p_r[5]),
	.ck(clk),
	.d(n212536));
   ms00f80 regtop_g_vs60p_r_reg_6_ (.o(g_vs60p_r[6]),
	.ck(clk),
	.d(n212535));
   ms00f80 regtop_g_vs60p_r_reg_0_ (.o(g_vs60p_r[0]),
	.ck(clk),
	.d(n212534));
   ms00f80 regtop_g_vden_r_reg (.o(g_vden_r),
	.ck(clk),
	.d(n212533));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_ferror_r_reg (.o(v_ferror_r),
	.ck(clk),
	.d(n253037));
   ms00f80 regtop_g_ferror_r_reg (.o(regtop_g_ferror_r),
	.ck(clk),
	.d(v_ferror_r));
   ms00f80 vldtop_vld_syndec_vld_vscdet_v_search_1st_r_reg (.o(vldtop_vld_syndec_vld_vscdet_v_search_1st_r),
	.ck(clk),
	.d(n212488));
   ms00f80 vldtop_vld_syndec_vld_vscdet_v_detvald_r_reg_0_ (.o(vldtop_vld_syndec_vld_vscdet_v_detvald_r[0]),
	.ck(clk),
	.d(n212487));
   ms00f80 vldtop_vld_syndec_vld_vscdet_v_detvald_r_reg_1_ (.o(vldtop_vld_syndec_vld_vscdet_v_detvald_r[1]),
	.ck(clk),
	.d(n212486));
   ms00f80 vldtop_vld_syndec_vld_vscdet_v_seqstrt_r_reg (.o(v_seqstrt_r),
	.ck(clk),
	.d(n212465));
   ms00f80 regtop_g_seqstrt_r_reg (.o(regtop_g_seqstrt_r),
	.ck(clk),
	.d(v_seqstrt_r));
   ms00f80 vldtop_vld_syndec_vld_vscdet_v_seqerr_r_reg (.o(vldtop_vld_syndec_vld_vscdet_v_seqerr_r),
	.ck(clk),
	.d(n212463));
   ms00f80 vldtop_vld_syndec_vld_vscdet_v_vld_state_r_reg_4_ (.o(v_vldstatus_r[4]),
	.ck(clk),
	.d(n243163));
   ms00f80 regtop_g_vldstatus_r_reg_4_ (.o(regtop_g_vldstatus_r[4]),
	.ck(clk),
	.d(v_vldstatus_r[4]));
   ms00f80 vldtop_vld_syndec_vld_vscdet_v_vld_state_r_reg_0_ (.o(v_vldstatus_r[0]),
	.ck(clk),
	.d(n243167));
   ms00f80 regtop_g_vldstatus_r_reg_0_ (.o(regtop_g_vldstatus_r[0]),
	.ck(clk),
	.d(v_vldstatus_r[0]));
   ms00f80 vldtop_vld_syndec_vld_vscdet_v_vld_state_r_reg_1_ (.o(v_vldstatus_r[1]),
	.ck(clk),
	.d(n243166));
   ms00f80 regtop_g_vldstatus_r_reg_1_ (.o(regtop_g_vldstatus_r[1]),
	.ck(clk),
	.d(v_vldstatus_r[1]));
   ms00f80 vldtop_vld_syndec_vld_seqhed_state_reg_0_ (.o(vldtop_vld_syndec_vld_seqhed_state_0_),
	.ck(clk),
	.d(n212425));
   ms00f80 vldtop_vld_syndec_vld_seqhed_pre_SHIFT_reg_3_ (.o(vldtop_vld_syndec_vld_seqhed_pre_SHIFT[3]),
	.ck(clk),
	.d(n212423));
   ms00f80 vldtop_vld_syndec_vld_seqhed_pre_SHIFT_reg_4_ (.o(vldtop_vld_syndec_vld_seqhed_pre_SHIFT[4]),
	.ck(clk),
	.d(n212416));
   ms00f80 vldtop_vld_syndec_vld_seqhed_pre_SHIFT_reg_1_ (.o(vldtop_vld_syndec_vld_seqhed_pre_SHIFT[1]),
	.ck(clk),
	.d(n212415));
   ms00f80 regtop_g_paramadr_r_reg_3_ (.o(regtop_g_paramadr_r[3]),
	.ck(clk),
	.d(v_paramadr_r[4]));
   ms00f80 regtop_g_paramadr_r_reg_2_ (.o(regtop_g_paramadr_r[2]),
	.ck(clk),
	.d(v_paramadr_r[4]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_nferror_r_reg (.o(v_nferror_r),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N44));
   ms00f80 regtop_g_nferror_r_reg (.o(regtop_g_nferror_r),
	.ck(clk),
	.d(v_nferror_r));
   ms00f80 regtop_g_paramadr_r_reg_6_ (.o(regtop_g_paramadr_r[6]),
	.ck(clk),
	.d(v_paramadr_r[4]));
   ms00f80 regtop_g_paramadr_r_reg_7_ (.o(regtop_g_paramadr_r[7]),
	.ck(clk),
	.d(v_paramadr_r[4]));
   ms00f80 regtop_g_paramadr_r_reg_0_ (.o(regtop_g_paramadr_r[0]),
	.ck(clk),
	.d(v_paramadr_r[4]));
   ms00f80 regtop_g_paramadr_r_reg_5_ (.o(regtop_g_paramadr_r[5]),
	.ck(clk),
	.d(v_paramadr_r[4]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramadr_r_reg_4_ (.o(v_paramadr_r[4]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N52));
   ms00f80 regtop_g_paramadr_r_reg_4_ (.o(regtop_g_paramadr_r[4]),
	.ck(clk),
	.d(v_paramadr_r[4]));
   ms00f80 regtop_g_nfst15_r_reg (.o(regtop_g_nfst_r[14]),
	.ck(clk),
	.d(n212292));
   ms00f80 regtop_g_fpst04_r_reg (.o(regtop_g_fpst_r[3]),
	.ck(clk),
	.d(n212291));
   ms00f80 regtop_g_nfst14_r_reg (.o(regtop_g_nfst_r[13]),
	.ck(clk),
	.d(n212290));
   ms00f80 regtop_g_fpst03_r_reg (.o(regtop_g_fpst_r[2]),
	.ck(clk),
	.d(n212289));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_0_ (.o(v_paramdata_r[0]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N463));
   ms00f80 regtop_g_paramdata_r_reg_0_ (.o(regtop_g_paramdata_r[0]),
	.ck(clk),
	.d(v_paramdata_r[0]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_1_ (.o(v_paramdata_r[1]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N464));
   ms00f80 regtop_g_paramdata_r_reg_1_ (.o(regtop_g_paramdata_r[1]),
	.ck(clk),
	.d(v_paramdata_r[1]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_2_ (.o(v_paramdata_r[2]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N465));
   ms00f80 regtop_g_paramdata_r_reg_2_ (.o(regtop_g_paramdata_r[2]),
	.ck(clk),
	.d(v_paramdata_r[2]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_3_ (.o(v_paramdata_r[3]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N466));
   ms00f80 regtop_g_paramdata_r_reg_3_ (.o(regtop_g_paramdata_r[3]),
	.ck(clk),
	.d(v_paramdata_r[3]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_4_ (.o(v_paramdata_r[4]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N467));
   ms00f80 regtop_g_paramdata_r_reg_4_ (.o(regtop_g_paramdata_r[4]),
	.ck(clk),
	.d(v_paramdata_r[4]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_5_ (.o(v_paramdata_r[5]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N468));
   ms00f80 regtop_g_paramdata_r_reg_5_ (.o(regtop_g_paramdata_r[5]),
	.ck(clk),
	.d(v_paramdata_r[5]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_6_ (.o(v_paramdata_r[6]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N469));
   ms00f80 regtop_g_paramdata_r_reg_6_ (.o(regtop_g_paramdata_r[6]),
	.ck(clk),
	.d(v_paramdata_r[6]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_16_ (.o(v_paramdata_r[16]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N479));
   ms00f80 regtop_g_paramdata_r_reg_16_ (.o(regtop_g_paramdata_r[16]),
	.ck(clk),
	.d(v_paramdata_r[16]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_7_ (.o(v_paramdata_r[7]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N470));
   ms00f80 regtop_g_paramdata_r_reg_7_ (.o(regtop_g_paramdata_r[7]),
	.ck(clk),
	.d(v_paramdata_r[7]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_8_ (.o(v_paramdata_r[8]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N471));
   ms00f80 regtop_g_paramdata_r_reg_8_ (.o(regtop_g_paramdata_r[8]),
	.ck(clk),
	.d(v_paramdata_r[8]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_9_ (.o(v_paramdata_r[9]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N472));
   ms00f80 regtop_g_paramdata_r_reg_9_ (.o(regtop_g_paramdata_r[9]),
	.ck(clk),
	.d(v_paramdata_r[9]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_10_ (.o(v_paramdata_r[10]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N473));
   ms00f80 regtop_g_paramdata_r_reg_10_ (.o(regtop_g_paramdata_r[10]),
	.ck(clk),
	.d(v_paramdata_r[10]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_11_ (.o(v_paramdata_r[11]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N474));
   ms00f80 regtop_g_paramdata_r_reg_11_ (.o(regtop_g_paramdata_r[11]),
	.ck(clk),
	.d(v_paramdata_r[11]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_12_ (.o(v_paramdata_r[12]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N475));
   ms00f80 regtop_g_paramdata_r_reg_12_ (.o(regtop_g_paramdata_r[12]),
	.ck(clk),
	.d(v_paramdata_r[12]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_13_ (.o(v_paramdata_r[13]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N476));
   ms00f80 regtop_g_paramdata_r_reg_13_ (.o(regtop_g_paramdata_r[13]),
	.ck(clk),
	.d(v_paramdata_r[13]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_14_ (.o(v_paramdata_r[14]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N477));
   ms00f80 regtop_g_paramdata_r_reg_14_ (.o(regtop_g_paramdata_r[14]),
	.ck(clk),
	.d(v_paramdata_r[14]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_15_ (.o(v_paramdata_r[15]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N478));
   ms00f80 regtop_g_paramdata_r_reg_15_ (.o(regtop_g_paramdata_r[15]),
	.ck(clk),
	.d(v_paramdata_r[15]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_17_ (.o(v_paramdata_r[17]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N480));
   ms00f80 regtop_g_paramdata_r_reg_17_ (.o(regtop_g_paramdata_r[17]),
	.ck(clk),
	.d(v_paramdata_r[17]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_18_ (.o(v_paramdata_r[18]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N481));
   ms00f80 regtop_g_paramdata_r_reg_18_ (.o(regtop_g_paramdata_r[18]),
	.ck(clk),
	.d(v_paramdata_r[18]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_19_ (.o(v_paramdata_r[19]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N482));
   ms00f80 regtop_g_paramdata_r_reg_19_ (.o(regtop_g_paramdata_r[19]),
	.ck(clk),
	.d(v_paramdata_r[19]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_20_ (.o(v_paramdata_r[20]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N483));
   ms00f80 regtop_g_paramdata_r_reg_20_ (.o(regtop_g_paramdata_r[20]),
	.ck(clk),
	.d(v_paramdata_r[20]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_21_ (.o(v_paramdata_r[21]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N484));
   ms00f80 regtop_g_paramdata_r_reg_21_ (.o(regtop_g_paramdata_r[21]),
	.ck(clk),
	.d(v_paramdata_r[21]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_22_ (.o(v_paramdata_r[22]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N485));
   ms00f80 regtop_g_paramdata_r_reg_22_ (.o(regtop_g_paramdata_r[22]),
	.ck(clk),
	.d(v_paramdata_r[22]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_23_ (.o(v_paramdata_r[23]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N486));
   ms00f80 regtop_g_paramdata_r_reg_23_ (.o(regtop_g_paramdata_r[23]),
	.ck(clk),
	.d(v_paramdata_r[23]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramdata_r_reg_24_ (.o(v_paramdata_r[24]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N487));
   ms00f80 regtop_g_paramdata_r_reg_24_ (.o(regtop_g_paramdata_r[24]),
	.ck(clk),
	.d(v_paramdata_r[24]));
   ms00f80 vldtop_vld_syndec_vld_outbuf_v_paramadr_r_reg_1_ (.o(v_paramadr_r[1]),
	.ck(clk),
	.d(vldtop_vld_syndec_vld_outbuf_N46));
   ms00f80 regtop_g_paramadr_r_reg_1_ (.o(regtop_g_paramadr_r[1]),
	.ck(clk),
	.d(v_paramadr_r[1]));
   ms00f80 regtop_g_usrd_r_reg_8_ (.o(regtop_g_usrd_r[8]),
	.ck(clk),
	.d(n212287));
   ms00f80 regtop_g_usrd_r_reg_31_ (.o(regtop_g_usrd_r[31]),
	.ck(clk),
	.d(n212286));
   ms00f80 regtop_g_usrd_r_reg_30_ (.o(regtop_g_usrd_r[30]),
	.ck(clk),
	.d(n212285));
   ms00f80 regtop_g_usrd_r_reg_29_ (.o(regtop_g_usrd_r[29]),
	.ck(clk),
	.d(n212284));
   ms00f80 regtop_g_usrd_r_reg_28_ (.o(regtop_g_usrd_r[28]),
	.ck(clk),
	.d(n212283));
   ms00f80 regtop_g_usrd_r_reg_27_ (.o(regtop_g_usrd_r[27]),
	.ck(clk),
	.d(n212282));
   ms00f80 regtop_g_usrd_r_reg_26_ (.o(regtop_g_usrd_r[26]),
	.ck(clk),
	.d(n212281));
   ms00f80 regtop_g_usrd_r_reg_25_ (.o(regtop_g_usrd_r[25]),
	.ck(clk),
	.d(n212280));
   ms00f80 regtop_g_usrd_r_reg_24_ (.o(regtop_g_usrd_r[24]),
	.ck(clk),
	.d(n212279));
   ms00f80 regtop_g_usrd_r_reg_23_ (.o(regtop_g_usrd_r[23]),
	.ck(clk),
	.d(n212278));
   ms00f80 regtop_g_usrd_r_reg_22_ (.o(regtop_g_usrd_r[22]),
	.ck(clk),
	.d(n212277));
   ms00f80 regtop_g_usrd_r_reg_21_ (.o(regtop_g_usrd_r[21]),
	.ck(clk),
	.d(n212276));
   ms00f80 regtop_g_usrd_r_reg_20_ (.o(regtop_g_usrd_r[20]),
	.ck(clk),
	.d(n212275));
   ms00f80 regtop_g_usrd_r_reg_19_ (.o(regtop_g_usrd_r[19]),
	.ck(clk),
	.d(n212274));
   ms00f80 regtop_g_usrd_r_reg_18_ (.o(regtop_g_usrd_r[18]),
	.ck(clk),
	.d(n212273));
   ms00f80 regtop_g_usrd_r_reg_17_ (.o(regtop_g_usrd_r[17]),
	.ck(clk),
	.d(n212272));
   ms00f80 regtop_g_usrd_r_reg_16_ (.o(regtop_g_usrd_r[16]),
	.ck(clk),
	.d(n212271));
   ms00f80 regtop_g_usrd_r_reg_15_ (.o(regtop_g_usrd_r[15]),
	.ck(clk),
	.d(n212270));
   ms00f80 regtop_g_usrd_r_reg_14_ (.o(regtop_g_usrd_r[14]),
	.ck(clk),
	.d(n212269));
   ms00f80 regtop_g_usrd_r_reg_13_ (.o(regtop_g_usrd_r[13]),
	.ck(clk),
	.d(n212268));
   ms00f80 regtop_g_usrd_r_reg_12_ (.o(regtop_g_usrd_r[12]),
	.ck(clk),
	.d(n212267));
   ms00f80 regtop_g_usrd_r_reg_11_ (.o(regtop_g_usrd_r[11]),
	.ck(clk),
	.d(n212266));
   ms00f80 regtop_g_usrd_r_reg_10_ (.o(regtop_g_usrd_r[10]),
	.ck(clk),
	.d(n212265));
   ms00f80 regtop_g_usrd_r_reg_9_ (.o(regtop_g_usrd_r[9]),
	.ck(clk),
	.d(n212264));
   ms00f80 regtop_g_cg_r_reg (.o(regtop_g_cg_r),
	.ck(clk),
	.d(n212263));
   ms00f80 regtop_g_bl_r_reg (.o(regtop_g_bl_r),
	.ck(clk),
	.d(n212262));
   ms00f80 regtop_g_mc_r_reg_0_ (.o(regtop_g_mc_r[0]),
	.ck(clk),
	.d(n212261));
   ms00f80 regtop_g_mc_r_reg_7_ (.o(regtop_g_mc_r[7]),
	.ck(clk),
	.d(n212260));
   ms00f80 regtop_g_mc_r_reg_6_ (.o(regtop_g_mc_r[6]),
	.ck(clk),
	.d(n212259));
   ms00f80 regtop_g_mc_r_reg_5_ (.o(regtop_g_mc_r[5]),
	.ck(clk),
	.d(n212258));
   ms00f80 regtop_g_mc_r_reg_4_ (.o(regtop_g_mc_r[4]),
	.ck(clk),
	.d(n212257));
   ms00f80 regtop_g_mc_r_reg_3_ (.o(regtop_g_mc_r[3]),
	.ck(clk),
	.d(n212256));
   ms00f80 regtop_g_mc_r_reg_2_ (.o(regtop_g_mc_r[2]),
	.ck(clk),
	.d(n212255));
   ms00f80 regtop_g_mc_r_reg_1_ (.o(regtop_g_mc_r[1]),
	.ck(clk),
	.d(n212254));
   ms00f80 regtop_g_vf_r_reg_0_ (.o(regtop_g_vf_r[0]),
	.ck(clk),
	.d(n212253));
   ms00f80 regtop_g_vf_r_reg_2_ (.o(regtop_g_vf_r[2]),
	.ck(clk),
	.d(n212252));
   ms00f80 regtop_g_vf_r_reg_1_ (.o(regtop_g_vf_r[1]),
	.ck(clk),
	.d(n212251));
   ms00f80 regtop_g_ps_r_reg (.o(regtop_g_ps_r),
	.ck(clk),
	.d(n212250));
   ms00f80 regtop_g_fpst02_r_reg (.o(regtop_g_fpst_r[1]),
	.ck(clk),
	.d(n212249));
   ms00f80 regtop_g_fcvo2_r_reg_0_ (.o(regtop_g_fcvo2_r[0]),
	.ck(clk),
	.d(n212248));
   ms00f80 regtop_g_fcvo2_r_reg_15_ (.o(regtop_g_fcvo2_r[15]),
	.ck(clk),
	.d(n212247));
   ms00f80 regtop_g_fcvo2_r_reg_14_ (.o(regtop_g_fcvo2_r[14]),
	.ck(clk),
	.d(n212246));
   ms00f80 regtop_g_fcvo2_r_reg_13_ (.o(regtop_g_fcvo2_r[13]),
	.ck(clk),
	.d(n212245));
   ms00f80 regtop_g_fcvo2_r_reg_12_ (.o(regtop_g_fcvo2_r[12]),
	.ck(clk),
	.d(n212244));
   ms00f80 regtop_g_fcvo2_r_reg_11_ (.o(regtop_g_fcvo2_r[11]),
	.ck(clk),
	.d(n212243));
   ms00f80 regtop_g_fcvo2_r_reg_10_ (.o(regtop_g_fcvo2_r[10]),
	.ck(clk),
	.d(n212242));
   ms00f80 regtop_g_fcvo2_r_reg_9_ (.o(regtop_g_fcvo2_r[9]),
	.ck(clk),
	.d(n212241));
   ms00f80 regtop_g_fcvo2_r_reg_8_ (.o(regtop_g_fcvo2_r[8]),
	.ck(clk),
	.d(n212240));
   ms00f80 regtop_g_fcvo2_r_reg_7_ (.o(regtop_g_fcvo2_r[7]),
	.ck(clk),
	.d(n212239));
   ms00f80 regtop_g_fcvo2_r_reg_6_ (.o(regtop_g_fcvo2_r[6]),
	.ck(clk),
	.d(n212238));
   ms00f80 regtop_g_fcvo2_r_reg_5_ (.o(regtop_g_fcvo2_r[5]),
	.ck(clk),
	.d(n212237));
   ms00f80 regtop_g_fcvo2_r_reg_4_ (.o(regtop_g_fcvo2_r[4]),
	.ck(clk),
	.d(n212236));
   ms00f80 regtop_g_fcvo2_r_reg_3_ (.o(regtop_g_fcvo2_r[3]),
	.ck(clk),
	.d(n212235));
   ms00f80 regtop_g_fcvo2_r_reg_2_ (.o(regtop_g_fcvo2_r[2]),
	.ck(clk),
	.d(n212234));
   ms00f80 regtop_g_fcvo2_r_reg_1_ (.o(regtop_g_fcvo2_r[1]),
	.ck(clk),
	.d(n212233));
   ms00f80 regtop_g_fcvo0_r_reg_0_ (.o(regtop_g_fcvo0_r[0]),
	.ck(clk),
	.d(n212232));
   ms00f80 regtop_g_fcvo0_r_reg_15_ (.o(regtop_g_fcvo0_r[15]),
	.ck(clk),
	.d(n212231));
   ms00f80 regtop_g_fcvo0_r_reg_14_ (.o(regtop_g_fcvo0_r[14]),
	.ck(clk),
	.d(n212230));
   ms00f80 regtop_g_fcvo0_r_reg_13_ (.o(regtop_g_fcvo0_r[13]),
	.ck(clk),
	.d(n212229));
   ms00f80 regtop_g_fcvo0_r_reg_12_ (.o(regtop_g_fcvo0_r[12]),
	.ck(clk),
	.d(n212228));
   ms00f80 regtop_g_fcvo0_r_reg_11_ (.o(regtop_g_fcvo0_r[11]),
	.ck(clk),
	.d(n212227));
   ms00f80 regtop_g_fcvo0_r_reg_10_ (.o(regtop_g_fcvo0_r[10]),
	.ck(clk),
	.d(n212226));
   ms00f80 regtop_g_fcvo0_r_reg_9_ (.o(regtop_g_fcvo0_r[9]),
	.ck(clk),
	.d(n212225));
   ms00f80 regtop_g_fcvo0_r_reg_8_ (.o(regtop_g_fcvo0_r[8]),
	.ck(clk),
	.d(n212224));
   ms00f80 regtop_g_fcvo0_r_reg_7_ (.o(regtop_g_fcvo0_r[7]),
	.ck(clk),
	.d(n212223));
   ms00f80 regtop_g_fcvo0_r_reg_6_ (.o(regtop_g_fcvo0_r[6]),
	.ck(clk),
	.d(n212222));
   ms00f80 regtop_g_fcvo0_r_reg_5_ (.o(regtop_g_fcvo0_r[5]),
	.ck(clk),
	.d(n212221));
   ms00f80 regtop_g_fcvo0_r_reg_4_ (.o(regtop_g_fcvo0_r[4]),
	.ck(clk),
	.d(n212220));
   ms00f80 regtop_g_fcvo0_r_reg_3_ (.o(regtop_g_fcvo0_r[3]),
	.ck(clk),
	.d(n212219));
   ms00f80 regtop_g_fcvo0_r_reg_2_ (.o(regtop_g_fcvo0_r[2]),
	.ck(clk),
	.d(n212218));
   ms00f80 regtop_g_fcvo0_r_reg_1_ (.o(regtop_g_fcvo0_r[1]),
	.ck(clk),
	.d(n212217));
   ms00f80 regtop_g_pis_r_reg_0_ (.o(regtop_g_pis_r[0]),
	.ck(clk),
	.d(n212216));
   ms00f80 regtop_g_pis_r_reg_1_ (.o(regtop_g_pis_r[1]),
	.ck(clk),
	.d(n212215));
   ms00f80 regtop_g_pct_r_reg_0_ (.o(regtop_g_pct_r[0]),
	.ck(clk),
	.d(n212214));
   ms00f80 regtop_g_pct_r_reg_2_ (.o(regtop_g_pct_r[2]),
	.ck(clk),
	.d(n212213));
   ms00f80 regtop_g_pct_r_reg_1_ (.o(regtop_g_pct_r[1]),
	.ck(clk),
	.d(n212212));
   ms00f80 regtop_g_vbsv_r_reg_0_ (.o(regtop_g_vbsv_r[0]),
	.ck(clk),
	.d(n212211));
   ms00f80 regtop_g_vbsv_r_reg_9_ (.o(regtop_g_vbsv_r[9]),
	.ck(clk),
	.d(n212210));
   ms00f80 regtop_g_vbsv_r_reg_8_ (.o(regtop_g_vbsv_r[8]),
	.ck(clk),
	.d(n212209));
   ms00f80 regtop_g_vbsv_r_reg_7_ (.o(regtop_g_vbsv_r[7]),
	.ck(clk),
	.d(n212208));
   ms00f80 regtop_g_vbsv_r_reg_6_ (.o(regtop_g_vbsv_r[6]),
	.ck(clk),
	.d(n212207));
   ms00f80 regtop_g_vbsv_r_reg_5_ (.o(regtop_g_vbsv_r[5]),
	.ck(clk),
	.d(n212206));
   ms00f80 regtop_g_vbsv_r_reg_4_ (.o(regtop_g_vbsv_r[4]),
	.ck(clk),
	.d(n212205));
   ms00f80 regtop_g_vbsv_r_reg_3_ (.o(regtop_g_vbsv_r[3]),
	.ck(clk),
	.d(n212204));
   ms00f80 regtop_g_vbsv_r_reg_2_ (.o(regtop_g_vbsv_r[2]),
	.ck(clk),
	.d(n212203));
   ms00f80 regtop_g_vbsv_r_reg_1_ (.o(regtop_g_vbsv_r[1]),
	.ck(clk),
	.d(n212202));
   ms00f80 regtop_g_nfst03_r_reg (.o(regtop_g_nfst_r[2]),
	.ck(clk),
	.d(n212201));
   ms00f80 regtop_g_nfst08_r_reg (.o(regtop_g_nfst_r[7]),
	.ck(clk),
	.d(n212200));
   ms00f80 regtop_g_fpst06_r_reg (.o(regtop_g_fpst_r[5]),
	.ck(clk),
	.d(n212199));
   ms00f80 regtop_g_nfst17_r_reg (.o(regtop_g_nfst_r[16]),
	.ck(clk),
	.d(n212198));
   ms00f80 regtop_g_dvs_r_reg_0_ (.o(regtop_g_dvs_r[0]),
	.ck(clk),
	.d(n212197));
   ms00f80 regtop_g_dvs_r_reg_13_ (.o(regtop_g_dvs_r[13]),
	.ck(clk),
	.d(n212196));
   ms00f80 regtop_g_dvs_r_reg_12_ (.o(regtop_g_dvs_r[12]),
	.ck(clk),
	.d(n212195));
   ms00f80 regtop_g_dvs_r_reg_11_ (.o(regtop_g_dvs_r[11]),
	.ck(clk),
	.d(n212194));
   ms00f80 regtop_g_dvs_r_reg_10_ (.o(regtop_g_dvs_r[10]),
	.ck(clk),
	.d(n212193));
   ms00f80 regtop_g_dvs_r_reg_9_ (.o(regtop_g_dvs_r[9]),
	.ck(clk),
	.d(n212192));
   ms00f80 regtop_g_dvs_r_reg_8_ (.o(regtop_g_dvs_r[8]),
	.ck(clk),
	.d(n212191));
   ms00f80 regtop_g_dvs_r_reg_7_ (.o(regtop_g_dvs_r[7]),
	.ck(clk),
	.d(n212190));
   ms00f80 regtop_g_dvs_r_reg_6_ (.o(regtop_g_dvs_r[6]),
	.ck(clk),
	.d(n212189));
   ms00f80 regtop_g_dvs_r_reg_5_ (.o(regtop_g_dvs_r[5]),
	.ck(clk),
	.d(n212188));
   ms00f80 regtop_g_dvs_r_reg_4_ (.o(regtop_g_dvs_r[4]),
	.ck(clk),
	.d(n212187));
   ms00f80 regtop_g_dvs_r_reg_3_ (.o(regtop_g_dvs_r[3]),
	.ck(clk),
	.d(n212186));
   ms00f80 regtop_g_dvs_r_reg_2_ (.o(regtop_g_dvs_r[2]),
	.ck(clk),
	.d(n212185));
   ms00f80 regtop_g_dvs_r_reg_1_ (.o(regtop_g_dvs_r[1]),
	.ck(clk),
	.d(n212184));
   ms00f80 regtop_g_cp_r_reg_0_ (.o(regtop_g_cp_r[0]),
	.ck(clk),
	.d(n212183));
   ms00f80 regtop_g_cp_r_reg_7_ (.o(regtop_g_cp_r[7]),
	.ck(clk),
	.d(n212182));
   ms00f80 regtop_g_cp_r_reg_6_ (.o(regtop_g_cp_r[6]),
	.ck(clk),
	.d(n212181));
   ms00f80 regtop_g_cp_r_reg_5_ (.o(regtop_g_cp_r[5]),
	.ck(clk),
	.d(n212180));
   ms00f80 regtop_g_cp_r_reg_4_ (.o(regtop_g_cp_r[4]),
	.ck(clk),
	.d(n212179));
   ms00f80 regtop_g_cp_r_reg_3_ (.o(regtop_g_cp_r[3]),
	.ck(clk),
	.d(n212178));
   ms00f80 regtop_g_cp_r_reg_2_ (.o(regtop_g_cp_r[2]),
	.ck(clk),
	.d(n212177));
   ms00f80 regtop_g_cp_r_reg_1_ (.o(regtop_g_cp_r[1]),
	.ck(clk),
	.d(n212176));
   ms00f80 regtop_g_ld_r_reg (.o(regtop_g_ld_r),
	.ck(clk),
	.d(n212175));
   ms00f80 regtop_g_fcvo1_r_reg_0_ (.o(regtop_g_fcvo1_r[0]),
	.ck(clk),
	.d(n212174));
   ms00f80 regtop_g_fcvo1_r_reg_15_ (.o(regtop_g_fcvo1_r[15]),
	.ck(clk),
	.d(n212173));
   ms00f80 regtop_g_fcvo1_r_reg_14_ (.o(regtop_g_fcvo1_r[14]),
	.ck(clk),
	.d(n212172));
   ms00f80 regtop_g_fcvo1_r_reg_13_ (.o(regtop_g_fcvo1_r[13]),
	.ck(clk),
	.d(n212171));
   ms00f80 regtop_g_fcvo1_r_reg_12_ (.o(regtop_g_fcvo1_r[12]),
	.ck(clk),
	.d(n212170));
   ms00f80 regtop_g_fcvo1_r_reg_11_ (.o(regtop_g_fcvo1_r[11]),
	.ck(clk),
	.d(n212169));
   ms00f80 regtop_g_fcvo1_r_reg_10_ (.o(regtop_g_fcvo1_r[10]),
	.ck(clk),
	.d(n212168));
   ms00f80 regtop_g_fcvo1_r_reg_9_ (.o(regtop_g_fcvo1_r[9]),
	.ck(clk),
	.d(n212167));
   ms00f80 regtop_g_fcvo1_r_reg_8_ (.o(regtop_g_fcvo1_r[8]),
	.ck(clk),
	.d(n212166));
   ms00f80 regtop_g_fcvo1_r_reg_7_ (.o(regtop_g_fcvo1_r[7]),
	.ck(clk),
	.d(n212165));
   ms00f80 regtop_g_fcvo1_r_reg_6_ (.o(regtop_g_fcvo1_r[6]),
	.ck(clk),
	.d(n212164));
   ms00f80 regtop_g_fcvo1_r_reg_5_ (.o(regtop_g_fcvo1_r[5]),
	.ck(clk),
	.d(n212163));
   ms00f80 regtop_g_fcvo1_r_reg_4_ (.o(regtop_g_fcvo1_r[4]),
	.ck(clk),
	.d(n212162));
   ms00f80 regtop_g_fcvo1_r_reg_3_ (.o(regtop_g_fcvo1_r[3]),
	.ck(clk),
	.d(n212161));
   ms00f80 regtop_g_fcvo1_r_reg_2_ (.o(regtop_g_fcvo1_r[2]),
	.ck(clk),
	.d(n212160));
   ms00f80 regtop_g_fcvo1_r_reg_1_ (.o(regtop_g_fcvo1_r[1]),
	.ck(clk),
	.d(n212159));
   ms00f80 regtop_g_cdf_r_reg (.o(regtop_g_cdf_r),
	.ck(clk),
	.d(n212158));
   ms00f80 regtop_g_mpeg_r_reg (.o(regtop_g_mpeg_r),
	.ck(clk),
	.d(n212157));
   ms00f80 regtop_g_nfst13_r_reg (.o(regtop_g_nfst_r[12]),
	.ck(clk),
	.d(n212156));
   ms00f80 regtop_g_nfst19_r_reg (.o(regtop_g_nfst_r[18]),
	.ck(clk),
	.d(n212155));
   ms00f80 regtop_g_nfst11_r_reg (.o(regtop_g_nfst_r[10]),
	.ck(clk),
	.d(n212154));
   ms00f80 regtop_g_adb_r_reg_0_ (.o(regtop_g_adb_r[0]),
	.ck(clk),
	.d(n212153));
   ms00f80 regtop_g_adb_r_reg_1_ (.o(regtop_g_adb_r[1]),
	.ck(clk),
	.d(n212152));
   ms00f80 regtop_g_adb_r_reg_2_ (.o(regtop_g_adb_r[2]),
	.ck(clk),
	.d(n212151));
   ms00f80 regtop_g_adb_r_reg_3_ (.o(regtop_g_adb_r[3]),
	.ck(clk),
	.d(n212150));
   ms00f80 regtop_g_adb_r_reg_4_ (.o(regtop_g_adb_r[4]),
	.ck(clk),
	.d(n212149));
   ms00f80 regtop_g_adb_r_reg_5_ (.o(regtop_g_adb_r[5]),
	.ck(clk),
	.d(n212148));
   ms00f80 regtop_g_adb_r_reg_6_ (.o(regtop_g_adb_r[6]),
	.ck(clk),
	.d(n212147));
   ms00f80 regtop_g_frc_r_reg_0_ (.o(regtop_g_frc_r[0]),
	.ck(clk),
	.d(n212146));
   ms00f80 regtop_g_frc_r_reg_3_ (.o(regtop_g_frc_r[3]),
	.ck(clk),
	.d(n212145));
   ms00f80 regtop_g_frc_r_reg_2_ (.o(regtop_g_frc_r[2]),
	.ck(clk),
	.d(n212144));
   ms00f80 regtop_g_frc_r_reg_1_ (.o(regtop_g_frc_r[1]),
	.ck(clk),
	.d(n212143));
   ms00f80 regtop_g_ari_r_reg_1_ (.o(regtop_g_ari_r[1]),
	.ck(clk),
	.d(n212142));
   ms00f80 regtop_g_ari_r_reg_2_ (.o(regtop_g_ari_r[2]),
	.ck(clk),
	.d(n212141));
   ms00f80 regtop_g_ari_r_reg_3_ (.o(regtop_g_ari_r[3]),
	.ck(clk),
	.d(n212140));
   ms00f80 regtop_g_ari_r_reg_0_ (.o(regtop_g_ari_r[0]),
	.ck(clk),
	.d(n212139));
   ms00f80 regtop_g_cf_r_reg_0_ (.o(regtop_g_cf_r[0]),
	.ck(clk),
	.d(n212138));
   ms00f80 regtop_g_cf_r_reg_1_ (.o(regtop_g_cf_r[1]),
	.ck(clk),
	.d(n212137));
   ms00f80 regtop_g_cd_r_reg (.o(regtop_g_cd_r),
	.ck(clk),
	.d(n212136));
   ms00f80 regtop_g_dhs_r_reg_0_ (.o(regtop_g_dhs_r[0]),
	.ck(clk),
	.d(n212135));
   ms00f80 regtop_g_dhs_r_reg_13_ (.o(regtop_g_dhs_r[13]),
	.ck(clk),
	.d(n212134));
   ms00f80 regtop_g_dhs_r_reg_12_ (.o(regtop_g_dhs_r[12]),
	.ck(clk),
	.d(n212133));
   ms00f80 regtop_g_dhs_r_reg_11_ (.o(regtop_g_dhs_r[11]),
	.ck(clk),
	.d(n212132));
   ms00f80 regtop_g_dhs_r_reg_10_ (.o(regtop_g_dhs_r[10]),
	.ck(clk),
	.d(n212131));
   ms00f80 regtop_g_dhs_r_reg_9_ (.o(regtop_g_dhs_r[9]),
	.ck(clk),
	.d(n212130));
   ms00f80 regtop_g_dhs_r_reg_8_ (.o(regtop_g_dhs_r[8]),
	.ck(clk),
	.d(n212129));
   ms00f80 regtop_g_dhs_r_reg_7_ (.o(regtop_g_dhs_r[7]),
	.ck(clk),
	.d(n212128));
   ms00f80 regtop_g_dhs_r_reg_6_ (.o(regtop_g_dhs_r[6]),
	.ck(clk),
	.d(n212127));
   ms00f80 regtop_g_dhs_r_reg_5_ (.o(regtop_g_dhs_r[5]),
	.ck(clk),
	.d(n212126));
   ms00f80 regtop_g_dhs_r_reg_4_ (.o(regtop_g_dhs_r[4]),
	.ck(clk),
	.d(n212125));
   ms00f80 regtop_g_dhs_r_reg_3_ (.o(regtop_g_dhs_r[3]),
	.ck(clk),
	.d(n212124));
   ms00f80 regtop_g_dhs_r_reg_2_ (.o(regtop_g_dhs_r[2]),
	.ck(clk),
	.d(n212123));
   ms00f80 regtop_g_dhs_r_reg_1_ (.o(regtop_g_dhs_r[1]),
	.ck(clk),
	.d(n212122));
   ms00f80 regtop_g_atscd_r_reg_8_ (.o(regtop_g_atscd_r[8]),
	.ck(clk),
	.d(n212121));
   ms00f80 regtop_g_atscd_r_reg_31_ (.o(regtop_g_atscd_r[31]),
	.ck(clk),
	.d(n212120));
   ms00f80 regtop_g_atscd_r_reg_30_ (.o(regtop_g_atscd_r[30]),
	.ck(clk),
	.d(n212119));
   ms00f80 regtop_g_atscd_r_reg_29_ (.o(regtop_g_atscd_r[29]),
	.ck(clk),
	.d(n212118));
   ms00f80 regtop_g_atscd_r_reg_28_ (.o(regtop_g_atscd_r[28]),
	.ck(clk),
	.d(n212117));
   ms00f80 regtop_g_atscd_r_reg_27_ (.o(regtop_g_atscd_r[27]),
	.ck(clk),
	.d(n212116));
   ms00f80 regtop_g_atscd_r_reg_26_ (.o(regtop_g_atscd_r[26]),
	.ck(clk),
	.d(n212115));
   ms00f80 regtop_g_atscd_r_reg_25_ (.o(regtop_g_atscd_r[25]),
	.ck(clk),
	.d(n212114));
   ms00f80 regtop_g_atscd_r_reg_24_ (.o(regtop_g_atscd_r[24]),
	.ck(clk),
	.d(n212113));
   ms00f80 regtop_g_atscd_r_reg_23_ (.o(regtop_g_atscd_r[23]),
	.ck(clk),
	.d(n212112));
   ms00f80 regtop_g_atscd_r_reg_22_ (.o(regtop_g_atscd_r[22]),
	.ck(clk),
	.d(n212111));
   ms00f80 regtop_g_atscd_r_reg_21_ (.o(regtop_g_atscd_r[21]),
	.ck(clk),
	.d(n212110));
   ms00f80 regtop_g_atscd_r_reg_20_ (.o(regtop_g_atscd_r[20]),
	.ck(clk),
	.d(n212109));
   ms00f80 regtop_g_atscd_r_reg_19_ (.o(regtop_g_atscd_r[19]),
	.ck(clk),
	.d(n212108));
   ms00f80 regtop_g_atscd_r_reg_18_ (.o(regtop_g_atscd_r[18]),
	.ck(clk),
	.d(n212107));
   ms00f80 regtop_g_atscd_r_reg_17_ (.o(regtop_g_atscd_r[17]),
	.ck(clk),
	.d(n212106));
   ms00f80 regtop_g_atscd_r_reg_16_ (.o(regtop_g_atscd_r[16]),
	.ck(clk),
	.d(n212105));
   ms00f80 regtop_g_atscd_r_reg_15_ (.o(regtop_g_atscd_r[15]),
	.ck(clk),
	.d(n212104));
   ms00f80 regtop_g_atscd_r_reg_14_ (.o(regtop_g_atscd_r[14]),
	.ck(clk),
	.d(n212103));
   ms00f80 regtop_g_atscd_r_reg_13_ (.o(regtop_g_atscd_r[13]),
	.ck(clk),
	.d(n212102));
   ms00f80 regtop_g_atscd_r_reg_12_ (.o(regtop_g_atscd_r[12]),
	.ck(clk),
	.d(n212101));
   ms00f80 regtop_g_atscd_r_reg_11_ (.o(regtop_g_atscd_r[11]),
	.ck(clk),
	.d(n212100));
   ms00f80 regtop_g_atscd_r_reg_10_ (.o(regtop_g_atscd_r[10]),
	.ck(clk),
	.d(n212099));
   ms00f80 regtop_g_atscd_r_reg_9_ (.o(regtop_g_atscd_r[9]),
	.ck(clk),
	.d(n212098));
   ms00f80 regtop_g_nfst16_r_reg (.o(regtop_g_nfst_r[15]),
	.ck(clk),
	.d(n212097));
   ms00f80 regtop_g_cpf_r_reg (.o(regtop_g_cpf_r),
	.ck(clk),
	.d(n212096));
   ms00f80 regtop_g_vd_r_reg_0_ (.o(regtop_g_vd_r[0]),
	.ck(clk),
	.d(n212095));
   ms00f80 regtop_g_vd_r_reg_15_ (.o(regtop_g_vd_r[15]),
	.ck(clk),
	.d(n212094));
   ms00f80 regtop_g_vd_r_reg_14_ (.o(regtop_g_vd_r[14]),
	.ck(clk),
	.d(n212093));
   ms00f80 regtop_g_vd_r_reg_13_ (.o(regtop_g_vd_r[13]),
	.ck(clk),
	.d(n212092));
   ms00f80 regtop_g_vd_r_reg_12_ (.o(regtop_g_vd_r[12]),
	.ck(clk),
	.d(n212091));
   ms00f80 regtop_g_vd_r_reg_11_ (.o(regtop_g_vd_r[11]),
	.ck(clk),
	.d(n212090));
   ms00f80 regtop_g_vd_r_reg_10_ (.o(regtop_g_vd_r[10]),
	.ck(clk),
	.d(n212089));
   ms00f80 regtop_g_vd_r_reg_9_ (.o(regtop_g_vd_r[9]),
	.ck(clk),
	.d(n212088));
   ms00f80 regtop_g_vd_r_reg_8_ (.o(regtop_g_vd_r[8]),
	.ck(clk),
	.d(n212087));
   ms00f80 regtop_g_vd_r_reg_7_ (.o(regtop_g_vd_r[7]),
	.ck(clk),
	.d(n212086));
   ms00f80 regtop_g_vd_r_reg_6_ (.o(regtop_g_vd_r[6]),
	.ck(clk),
	.d(n212085));
   ms00f80 regtop_g_vd_r_reg_5_ (.o(regtop_g_vd_r[5]),
	.ck(clk),
	.d(n212084));
   ms00f80 regtop_g_vd_r_reg_4_ (.o(regtop_g_vd_r[4]),
	.ck(clk),
	.d(n212083));
   ms00f80 regtop_g_vd_r_reg_3_ (.o(regtop_g_vd_r[3]),
	.ck(clk),
	.d(n212082));
   ms00f80 regtop_g_vd_r_reg_2_ (.o(regtop_g_vd_r[2]),
	.ck(clk),
	.d(n212081));
   ms00f80 regtop_g_vd_r_reg_1_ (.o(regtop_g_vd_r[1]),
	.ck(clk),
	.d(n212080));
   ms00f80 regtop_g_pf_r_reg (.o(regtop_g_pf_r),
	.ck(clk),
	.d(n212079));
   ms00f80 regtop_g_rff_r_reg (.o(regtop_g_rff_r),
	.ck(clk),
	.d(n212078));
   ms00f80 regtop_g_tff_r_reg (.o(regtop_g_tff_r),
	.ck(clk),
	.d(n212077));
   ms00f80 regtop_g_nfco_r_reg_0_ (.o(regtop_g_nfco_r[0]),
	.ck(clk),
	.d(n212076));
   ms00f80 regtop_g_nfco_r_reg_1_ (.o(regtop_g_nfco_r[1]),
	.ck(clk),
	.d(n212075));
   ms00f80 regtop_g_fcho1_r_reg_0_ (.o(regtop_g_fcho1_r[0]),
	.ck(clk),
	.d(n212074));
   ms00f80 regtop_g_fcho1_r_reg_15_ (.o(regtop_g_fcho1_r[15]),
	.ck(clk),
	.d(n212073));
   ms00f80 regtop_g_fcho1_r_reg_14_ (.o(regtop_g_fcho1_r[14]),
	.ck(clk),
	.d(n212072));
   ms00f80 regtop_g_fcho1_r_reg_13_ (.o(regtop_g_fcho1_r[13]),
	.ck(clk),
	.d(n212071));
   ms00f80 regtop_g_fcho1_r_reg_12_ (.o(regtop_g_fcho1_r[12]),
	.ck(clk),
	.d(n212070));
   ms00f80 regtop_g_fcho1_r_reg_11_ (.o(regtop_g_fcho1_r[11]),
	.ck(clk),
	.d(n212069));
   ms00f80 regtop_g_fcho1_r_reg_10_ (.o(regtop_g_fcho1_r[10]),
	.ck(clk),
	.d(n212068));
   ms00f80 regtop_g_fcho1_r_reg_9_ (.o(regtop_g_fcho1_r[9]),
	.ck(clk),
	.d(n212067));
   ms00f80 regtop_g_fcho1_r_reg_8_ (.o(regtop_g_fcho1_r[8]),
	.ck(clk),
	.d(n212066));
   ms00f80 regtop_g_fcho1_r_reg_7_ (.o(regtop_g_fcho1_r[7]),
	.ck(clk),
	.d(n212065));
   ms00f80 regtop_g_fcho1_r_reg_6_ (.o(regtop_g_fcho1_r[6]),
	.ck(clk),
	.d(n212064));
   ms00f80 regtop_g_fcho1_r_reg_5_ (.o(regtop_g_fcho1_r[5]),
	.ck(clk),
	.d(n212063));
   ms00f80 regtop_g_fcho1_r_reg_4_ (.o(regtop_g_fcho1_r[4]),
	.ck(clk),
	.d(n212062));
   ms00f80 regtop_g_fcho1_r_reg_3_ (.o(regtop_g_fcho1_r[3]),
	.ck(clk),
	.d(n212061));
   ms00f80 regtop_g_fcho1_r_reg_2_ (.o(regtop_g_fcho1_r[2]),
	.ck(clk),
	.d(n212060));
   ms00f80 regtop_g_fcho1_r_reg_1_ (.o(regtop_g_fcho1_r[1]),
	.ck(clk),
	.d(n212059));
   ms00f80 regtop_g_nfst01_r_reg (.o(regtop_g_nfst_r[0]),
	.ck(clk),
	.d(n212058));
   ms00f80 regtop_g_nfst06_r_reg (.o(regtop_g_nfst_r[5]),
	.ck(clk),
	.d(n212057));
   ms00f80 regtop_g_nfst09_r_reg (.o(regtop_g_nfst_r[8]),
	.ck(clk),
	.d(n212056));
   ms00f80 regtop_g_udb1_r_reg_0_ (.o(regtop_g_udb1_r[0]),
	.ck(clk),
	.d(n212055));
   ms00f80 regtop_g_udb1_r_reg_1_ (.o(regtop_g_udb1_r[1]),
	.ck(clk),
	.d(n212054));
   ms00f80 regtop_g_udb1_r_reg_2_ (.o(regtop_g_udb1_r[2]),
	.ck(clk),
	.d(n212053));
   ms00f80 regtop_g_udb1_r_reg_3_ (.o(regtop_g_udb1_r[3]),
	.ck(clk),
	.d(n212052));
   ms00f80 regtop_g_udb1_r_reg_4_ (.o(regtop_g_udb1_r[4]),
	.ck(clk),
	.d(n212051));
   ms00f80 regtop_g_udb1_r_reg_5_ (.o(regtop_g_udb1_r[5]),
	.ck(clk),
	.d(n212050));
   ms00f80 regtop_g_udb1_r_reg_6_ (.o(regtop_g_udb1_r[6]),
	.ck(clk),
	.d(n212049));
   ms00f80 regtop_g_brv_r_reg_0_ (.o(regtop_g_brv_r[0]),
	.ck(clk),
	.d(n212048));
   ms00f80 regtop_g_brv_r_reg_17_ (.o(regtop_g_brv_r[17]),
	.ck(clk),
	.d(n212047));
   ms00f80 regtop_g_brv_r_reg_16_ (.o(regtop_g_brv_r[16]),
	.ck(clk),
	.d(n212046));
   ms00f80 regtop_g_brv_r_reg_15_ (.o(regtop_g_brv_r[15]),
	.ck(clk),
	.d(n212045));
   ms00f80 regtop_g_brv_r_reg_14_ (.o(regtop_g_brv_r[14]),
	.ck(clk),
	.d(n212044));
   ms00f80 regtop_g_brv_r_reg_13_ (.o(regtop_g_brv_r[13]),
	.ck(clk),
	.d(n212043));
   ms00f80 regtop_g_brv_r_reg_12_ (.o(regtop_g_brv_r[12]),
	.ck(clk),
	.d(n212042));
   ms00f80 regtop_g_brv_r_reg_11_ (.o(regtop_g_brv_r[11]),
	.ck(clk),
	.d(n212041));
   ms00f80 regtop_g_brv_r_reg_10_ (.o(regtop_g_brv_r[10]),
	.ck(clk),
	.d(n212040));
   ms00f80 regtop_g_brv_r_reg_9_ (.o(regtop_g_brv_r[9]),
	.ck(clk),
	.d(n212039));
   ms00f80 regtop_g_brv_r_reg_8_ (.o(regtop_g_brv_r[8]),
	.ck(clk),
	.d(n212038));
   ms00f80 regtop_g_brv_r_reg_7_ (.o(regtop_g_brv_r[7]),
	.ck(clk),
	.d(n212037));
   ms00f80 regtop_g_brv_r_reg_6_ (.o(regtop_g_brv_r[6]),
	.ck(clk),
	.d(n212036));
   ms00f80 regtop_g_brv_r_reg_5_ (.o(regtop_g_brv_r[5]),
	.ck(clk),
	.d(n212035));
   ms00f80 regtop_g_brv_r_reg_4_ (.o(regtop_g_brv_r[4]),
	.ck(clk),
	.d(n212034));
   ms00f80 regtop_g_brv_r_reg_3_ (.o(regtop_g_brv_r[3]),
	.ck(clk),
	.d(n212033));
   ms00f80 regtop_g_brv_r_reg_2_ (.o(regtop_g_brv_r[2]),
	.ck(clk),
	.d(n212032));
   ms00f80 regtop_g_brv_r_reg_1_ (.o(regtop_g_brv_r[1]),
	.ck(clk),
	.d(n212031));
   ms00f80 regtop_g_tr_r_reg_0_ (.o(regtop_g_tr_r[0]),
	.ck(clk),
	.d(n212030));
   ms00f80 regtop_g_tr_r_reg_9_ (.o(regtop_g_tr_r[9]),
	.ck(clk),
	.d(n212029));
   ms00f80 regtop_g_tr_r_reg_8_ (.o(regtop_g_tr_r[8]),
	.ck(clk),
	.d(n212028));
   ms00f80 regtop_g_tr_r_reg_7_ (.o(regtop_g_tr_r[7]),
	.ck(clk),
	.d(n212027));
   ms00f80 regtop_g_tr_r_reg_6_ (.o(regtop_g_tr_r[6]),
	.ck(clk),
	.d(n212026));
   ms00f80 regtop_g_tr_r_reg_5_ (.o(regtop_g_tr_r[5]),
	.ck(clk),
	.d(n212025));
   ms00f80 regtop_g_tr_r_reg_4_ (.o(regtop_g_tr_r[4]),
	.ck(clk),
	.d(n212024));
   ms00f80 regtop_g_tr_r_reg_3_ (.o(regtop_g_tr_r[3]),
	.ck(clk),
	.d(n212023));
   ms00f80 regtop_g_tr_r_reg_2_ (.o(regtop_g_tr_r[2]),
	.ck(clk),
	.d(n212022));
   ms00f80 regtop_g_tr_r_reg_1_ (.o(regtop_g_tr_r[1]),
	.ck(clk),
	.d(n212021));
   ms00f80 regtop_g_scp_r_reg_0_ (.o(regtop_g_scp_r[0]),
	.ck(clk),
	.d(n212020));
   ms00f80 regtop_g_scp_r_reg_7_ (.o(regtop_g_scp_r[7]),
	.ck(clk),
	.d(n212019));
   ms00f80 regtop_g_scp_r_reg_6_ (.o(regtop_g_scp_r[6]),
	.ck(clk),
	.d(n212018));
   ms00f80 regtop_g_scp_r_reg_5_ (.o(regtop_g_scp_r[5]),
	.ck(clk),
	.d(n212017));
   ms00f80 regtop_g_scp_r_reg_4_ (.o(regtop_g_scp_r[4]),
	.ck(clk),
	.d(n212016));
   ms00f80 regtop_g_scp_r_reg_3_ (.o(regtop_g_scp_r[3]),
	.ck(clk),
	.d(n212015));
   ms00f80 regtop_g_scp_r_reg_2_ (.o(regtop_g_scp_r[2]),
	.ck(clk),
	.d(n212014));
   ms00f80 regtop_g_scp_r_reg_1_ (.o(regtop_g_scp_r[1]),
	.ck(clk),
	.d(n212013));
   ms00f80 regtop_g_ba_r_reg_1_ (.o(regtop_g_ba_r[1]),
	.ck(clk),
	.d(n212012));
   ms00f80 regtop_g_ba_r_reg_2_ (.o(regtop_g_ba_r[2]),
	.ck(clk),
	.d(n212011));
   ms00f80 regtop_g_ba_r_reg_3_ (.o(regtop_g_ba_r[3]),
	.ck(clk),
	.d(n212010));
   ms00f80 regtop_g_ba_r_reg_4_ (.o(regtop_g_ba_r[4]),
	.ck(clk),
	.d(n212009));
   ms00f80 regtop_g_ba_r_reg_5_ (.o(regtop_g_ba_r[5]),
	.ck(clk),
	.d(n212008));
   ms00f80 regtop_g_ba_r_reg_6_ (.o(regtop_g_ba_r[6]),
	.ck(clk),
	.d(n212007));
   ms00f80 regtop_g_ba_r_reg_0_ (.o(regtop_g_ba_r[0]),
	.ck(clk),
	.d(n212006));
   ms00f80 regtop_g_sc_r_reg (.o(regtop_g_sc_r),
	.ck(clk),
	.d(n212005));
   ms00f80 regtop_g_fs_r_reg_1_ (.o(regtop_g_fs_r[1]),
	.ck(clk),
	.d(n212004));
   ms00f80 regtop_g_fs_r_reg_2_ (.o(regtop_g_fs_r[2]),
	.ck(clk),
	.d(n212003));
   ms00f80 regtop_g_fs_r_reg_0_ (.o(regtop_g_fs_r[0]),
	.ck(clk),
	.d(n212002));
   ms00f80 regtop_g_va_r_reg (.o(regtop_g_va_r),
	.ck(clk),
	.d(n212001));
   ms00f80 regtop_g_fcho0_r_reg_0_ (.o(regtop_g_fcho0_r[0]),
	.ck(clk),
	.d(n212000));
   ms00f80 regtop_g_fcho0_r_reg_15_ (.o(regtop_g_fcho0_r[15]),
	.ck(clk),
	.d(n211999));
   ms00f80 regtop_g_fcho0_r_reg_14_ (.o(regtop_g_fcho0_r[14]),
	.ck(clk),
	.d(n211998));
   ms00f80 regtop_g_fcho0_r_reg_13_ (.o(regtop_g_fcho0_r[13]),
	.ck(clk),
	.d(n211997));
   ms00f80 regtop_g_fcho0_r_reg_12_ (.o(regtop_g_fcho0_r[12]),
	.ck(clk),
	.d(n211996));
   ms00f80 regtop_g_fcho0_r_reg_11_ (.o(regtop_g_fcho0_r[11]),
	.ck(clk),
	.d(n211995));
   ms00f80 regtop_g_fcho0_r_reg_10_ (.o(regtop_g_fcho0_r[10]),
	.ck(clk),
	.d(n211994));
   ms00f80 regtop_g_fcho0_r_reg_9_ (.o(regtop_g_fcho0_r[9]),
	.ck(clk),
	.d(n211993));
   ms00f80 regtop_g_fcho0_r_reg_8_ (.o(regtop_g_fcho0_r[8]),
	.ck(clk),
	.d(n211992));
   ms00f80 regtop_g_fcho0_r_reg_7_ (.o(regtop_g_fcho0_r[7]),
	.ck(clk),
	.d(n211991));
   ms00f80 regtop_g_fcho0_r_reg_6_ (.o(regtop_g_fcho0_r[6]),
	.ck(clk),
	.d(n211990));
   ms00f80 regtop_g_fcho0_r_reg_5_ (.o(regtop_g_fcho0_r[5]),
	.ck(clk),
	.d(n211989));
   ms00f80 regtop_g_fcho0_r_reg_4_ (.o(regtop_g_fcho0_r[4]),
	.ck(clk),
	.d(n211988));
   ms00f80 regtop_g_fcho0_r_reg_3_ (.o(regtop_g_fcho0_r[3]),
	.ck(clk),
	.d(n211987));
   ms00f80 regtop_g_fcho0_r_reg_2_ (.o(regtop_g_fcho0_r[2]),
	.ck(clk),
	.d(n211986));
   ms00f80 regtop_g_fcho0_r_reg_1_ (.o(regtop_g_fcho0_r[1]),
	.ck(clk),
	.d(n211985));
   ms00f80 regtop_g_fcho2_r_reg_0_ (.o(regtop_g_fcho2_r[0]),
	.ck(clk),
	.d(n211984));
   ms00f80 regtop_g_fcho2_r_reg_15_ (.o(regtop_g_fcho2_r[15]),
	.ck(clk),
	.d(n211983));
   ms00f80 regtop_g_fcho2_r_reg_14_ (.o(regtop_g_fcho2_r[14]),
	.ck(clk),
	.d(n211982));
   ms00f80 regtop_g_fcho2_r_reg_13_ (.o(regtop_g_fcho2_r[13]),
	.ck(clk),
	.d(n211981));
   ms00f80 regtop_g_fcho2_r_reg_12_ (.o(regtop_g_fcho2_r[12]),
	.ck(clk),
	.d(n211980));
   ms00f80 regtop_g_fcho2_r_reg_11_ (.o(regtop_g_fcho2_r[11]),
	.ck(clk),
	.d(n211979));
   ms00f80 regtop_g_fcho2_r_reg_10_ (.o(regtop_g_fcho2_r[10]),
	.ck(clk),
	.d(n211978));
   ms00f80 regtop_g_fcho2_r_reg_9_ (.o(regtop_g_fcho2_r[9]),
	.ck(clk),
	.d(n211977));
   ms00f80 regtop_g_fcho2_r_reg_8_ (.o(regtop_g_fcho2_r[8]),
	.ck(clk),
	.d(n211976));
   ms00f80 regtop_g_fcho2_r_reg_7_ (.o(regtop_g_fcho2_r[7]),
	.ck(clk),
	.d(n211975));
   ms00f80 regtop_g_fcho2_r_reg_6_ (.o(regtop_g_fcho2_r[6]),
	.ck(clk),
	.d(n211974));
   ms00f80 regtop_g_fcho2_r_reg_5_ (.o(regtop_g_fcho2_r[5]),
	.ck(clk),
	.d(n211973));
   ms00f80 regtop_g_fcho2_r_reg_4_ (.o(regtop_g_fcho2_r[4]),
	.ck(clk),
	.d(n211972));
   ms00f80 regtop_g_fcho2_r_reg_3_ (.o(regtop_g_fcho2_r[3]),
	.ck(clk),
	.d(n211971));
   ms00f80 regtop_g_fcho2_r_reg_2_ (.o(regtop_g_fcho2_r[2]),
	.ck(clk),
	.d(n211970));
   ms00f80 regtop_g_fcho2_r_reg_1_ (.o(regtop_g_fcho2_r[1]),
	.ck(clk),
	.d(n211969));
   ms00f80 regtop_g_nfst10_r_reg (.o(regtop_g_nfst_r[9]),
	.ck(clk),
	.d(n211968));
   ms00f80 regtop_g_nfst02_r_reg (.o(regtop_g_nfst_r[1]),
	.ck(clk),
	.d(n211967));
   ms00f80 regtop_g_nfst12_r_reg (.o(regtop_g_nfst_r[11]),
	.ck(clk),
	.d(n211966));
   ms00f80 regtop_g_nfst05_r_reg (.o(regtop_g_nfst_r[4]),
	.ck(clk),
	.d(n211965));
   ms00f80 regtop_g_nfst18_r_reg (.o(regtop_g_nfst_r[17]),
	.ck(clk),
	.d(n211964));
   ms00f80 regtop_g_nfst07_r_reg (.o(regtop_g_nfst_r[6]),
	.ck(clk),
	.d(n211963));
   ms00f80 regtop_g_fpst05_r_reg (.o(regtop_g_fpst_r[4]),
	.ck(clk),
	.d(n211962));
   ms00f80 regtop_g_udb2_r_reg_0_ (.o(regtop_g_udb2_r[0]),
	.ck(clk),
	.d(n211961));
   ms00f80 regtop_g_udb2_r_reg_1_ (.o(regtop_g_udb2_r[1]),
	.ck(clk),
	.d(n211960));
   ms00f80 regtop_g_udb2_r_reg_2_ (.o(regtop_g_udb2_r[2]),
	.ck(clk),
	.d(n211959));
   ms00f80 regtop_g_udb2_r_reg_3_ (.o(regtop_g_udb2_r[3]),
	.ck(clk),
	.d(n211958));
   ms00f80 regtop_g_udb2_r_reg_4_ (.o(regtop_g_udb2_r[4]),
	.ck(clk),
	.d(n211957));
   ms00f80 regtop_g_udb2_r_reg_5_ (.o(regtop_g_udb2_r[5]),
	.ck(clk),
	.d(n211956));
   ms00f80 regtop_g_udb2_r_reg_6_ (.o(regtop_g_udb2_r[6]),
	.ck(clk),
	.d(n211955));
   ms00f80 regtop_g_udb0_r_reg_0_ (.o(regtop_g_udb0_r[0]),
	.ck(clk),
	.d(n211954));
   ms00f80 regtop_g_udb0_r_reg_1_ (.o(regtop_g_udb0_r[1]),
	.ck(clk),
	.d(n211953));
   ms00f80 regtop_g_udb0_r_reg_2_ (.o(regtop_g_udb0_r[2]),
	.ck(clk),
	.d(n211952));
   ms00f80 regtop_g_udb0_r_reg_3_ (.o(regtop_g_udb0_r[3]),
	.ck(clk),
	.d(n211951));
   ms00f80 regtop_g_udb0_r_reg_4_ (.o(regtop_g_udb0_r[4]),
	.ck(clk),
	.d(n211950));
   ms00f80 regtop_g_udb0_r_reg_5_ (.o(regtop_g_udb0_r[5]),
	.ck(clk),
	.d(n211949));
   ms00f80 regtop_g_udb0_r_reg_6_ (.o(regtop_g_udb0_r[6]),
	.ck(clk),
	.d(n211948));
   ms00f80 regtop_g_vsv_r_reg_0_ (.o(regtop_g_vsv_r[0]),
	.ck(clk),
	.d(n211940));
   ms00f80 regtop_g_vsv_r_reg_11_ (.o(regtop_g_vsv_r[11]),
	.ck(clk),
	.d(n211939));
   ms00f80 regtop_g_vsv_r_reg_10_ (.o(regtop_g_vsv_r[10]),
	.ck(clk),
	.d(n211938));
   ms00f80 regtop_g_vsv_r_reg_9_ (.o(regtop_g_vsv_r[9]),
	.ck(clk),
	.d(n211937));
   ms00f80 regtop_g_vsv_r_reg_8_ (.o(regtop_g_vsv_r[8]),
	.ck(clk),
	.d(n211936));
   ms00f80 regtop_g_vsv_r_reg_7_ (.o(regtop_g_vsv_r[7]),
	.ck(clk),
	.d(n211935));
   ms00f80 regtop_g_vsv_r_reg_6_ (.o(regtop_g_vsv_r[6]),
	.ck(clk),
	.d(n211934));
   ms00f80 regtop_g_vsv_r_reg_5_ (.o(regtop_g_vsv_r[5]),
	.ck(clk),
	.d(n211933));
   ms00f80 regtop_g_vsv_r_reg_4_ (.o(regtop_g_vsv_r[4]),
	.ck(clk),
	.d(n211932));
   ms00f80 regtop_g_vsv_r_reg_3_ (.o(regtop_g_vsv_r[3]),
	.ck(clk),
	.d(n211931));
   ms00f80 regtop_g_vsv_r_reg_2_ (.o(regtop_g_vsv_r[2]),
	.ck(clk),
	.d(n211930));
   ms00f80 regtop_g_vsv_r_reg_1_ (.o(regtop_g_vsv_r[1]),
	.ck(clk),
	.d(n211929));
   ms00f80 regtop_g_hsv_r_reg_1_ (.o(regtop_g_hsv_r[1]),
	.ck(clk),
	.d(n211928));
   ms00f80 regtop_g_hsv_r_reg_2_ (.o(regtop_g_hsv_r[2]),
	.ck(clk),
	.d(n211927));
   ms00f80 regtop_g_hsv_r_reg_3_ (.o(regtop_g_hsv_r[3]),
	.ck(clk),
	.d(n211926));
   ms00f80 regtop_g_hsv_r_reg_4_ (.o(regtop_g_hsv_r[4]),
	.ck(clk),
	.d(n211925));
   ms00f80 regtop_g_hsv_r_reg_5_ (.o(regtop_g_hsv_r[5]),
	.ck(clk),
	.d(n211924));
   ms00f80 regtop_g_hsv_r_reg_6_ (.o(regtop_g_hsv_r[6]),
	.ck(clk),
	.d(n211923));
   ms00f80 regtop_g_hsv_r_reg_7_ (.o(regtop_g_hsv_r[7]),
	.ck(clk),
	.d(n211922));
   ms00f80 regtop_g_hsv_r_reg_8_ (.o(regtop_g_hsv_r[8]),
	.ck(clk),
	.d(n211921));
   ms00f80 regtop_g_hsv_r_reg_9_ (.o(regtop_g_hsv_r[9]),
	.ck(clk),
	.d(n211920));
   ms00f80 regtop_g_hsv_r_reg_10_ (.o(regtop_g_hsv_r[10]),
	.ck(clk),
	.d(n211919));
   ms00f80 regtop_g_hsv_r_reg_11_ (.o(regtop_g_hsv_r[11]),
	.ck(clk),
	.d(n211918));
   ms00f80 regtop_g_hsv_r_reg_0_ (.o(regtop_g_hsv_r[0]),
	.ck(clk),
	.d(n211917));
   ms00f80 regtop_g_pali_r_reg_0_ (.o(regtop_g_pali_r[0]),
	.ck(clk),
	.d(n211916));
   ms00f80 regtop_g_pali_r_reg_7_ (.o(regtop_g_pali_r[7]),
	.ck(clk),
	.d(n211915));
   ms00f80 regtop_g_pali_r_reg_6_ (.o(regtop_g_pali_r[6]),
	.ck(clk),
	.d(n211914));
   ms00f80 regtop_g_pali_r_reg_5_ (.o(regtop_g_pali_r[5]),
	.ck(clk),
	.d(n211913));
   ms00f80 regtop_g_pali_r_reg_4_ (.o(regtop_g_pali_r[4]),
	.ck(clk),
	.d(n211912));
   ms00f80 regtop_g_pali_r_reg_3_ (.o(regtop_g_pali_r[3]),
	.ck(clk),
	.d(n211911));
   ms00f80 regtop_g_pali_r_reg_2_ (.o(regtop_g_pali_r[2]),
	.ck(clk),
	.d(n211910));
   ms00f80 regtop_g_pali_r_reg_1_ (.o(regtop_g_pali_r[1]),
	.ck(clk),
	.d(n211909));
   ms00f80 regtop_g_tc_r_reg_0_ (.o(regtop_g_tc_r[0]),
	.ck(clk),
	.d(n211908));
   ms00f80 regtop_g_tc_r_reg_7_ (.o(regtop_g_tc_r[7]),
	.ck(clk),
	.d(n211907));
   ms00f80 regtop_g_tc_r_reg_6_ (.o(regtop_g_tc_r[6]),
	.ck(clk),
	.d(n211906));
   ms00f80 regtop_g_tc_r_reg_5_ (.o(regtop_g_tc_r[5]),
	.ck(clk),
	.d(n211905));
   ms00f80 regtop_g_tc_r_reg_4_ (.o(regtop_g_tc_r[4]),
	.ck(clk),
	.d(n211904));
   ms00f80 regtop_g_tc_r_reg_3_ (.o(regtop_g_tc_r[3]),
	.ck(clk),
	.d(n211903));
   ms00f80 regtop_g_tc_r_reg_2_ (.o(regtop_g_tc_r[2]),
	.ck(clk),
	.d(n211902));
   ms00f80 regtop_g_tc_r_reg_1_ (.o(regtop_g_tc_r[1]),
	.ck(clk),
	.d(n211901));
   ms00f80 regtop_g_tmc_r_reg_0_ (.o(regtop_g_tmc_r[0]),
	.ck(clk),
	.d(n211900));
   ms00f80 regtop_g_tmc_r_reg_23_ (.o(regtop_g_tmc_r[23]),
	.ck(clk),
	.d(n211899));
   ms00f80 regtop_g_tmc_r_reg_22_ (.o(regtop_g_tmc_r[22]),
	.ck(clk),
	.d(n211898));
   ms00f80 regtop_g_tmc_r_reg_21_ (.o(regtop_g_tmc_r[21]),
	.ck(clk),
	.d(n211897));
   ms00f80 regtop_g_tmc_r_reg_20_ (.o(regtop_g_tmc_r[20]),
	.ck(clk),
	.d(n211896));
   ms00f80 regtop_g_tmc_r_reg_19_ (.o(regtop_g_tmc_r[19]),
	.ck(clk),
	.d(n211895));
   ms00f80 regtop_g_tmc_r_reg_18_ (.o(regtop_g_tmc_r[18]),
	.ck(clk),
	.d(n211894));
   ms00f80 regtop_g_tmc_r_reg_17_ (.o(regtop_g_tmc_r[17]),
	.ck(clk),
	.d(n211893));
   ms00f80 regtop_g_tmc_r_reg_16_ (.o(regtop_g_tmc_r[16]),
	.ck(clk),
	.d(n211892));
   ms00f80 regtop_g_tmc_r_reg_15_ (.o(regtop_g_tmc_r[15]),
	.ck(clk),
	.d(n211891));
   ms00f80 regtop_g_tmc_r_reg_14_ (.o(regtop_g_tmc_r[14]),
	.ck(clk),
	.d(n211890));
   ms00f80 regtop_g_tmc_r_reg_13_ (.o(regtop_g_tmc_r[13]),
	.ck(clk),
	.d(n211889));
   ms00f80 regtop_g_tmc_r_reg_12_ (.o(regtop_g_tmc_r[12]),
	.ck(clk),
	.d(n211888));
   ms00f80 regtop_g_tmc_r_reg_11_ (.o(regtop_g_tmc_r[11]),
	.ck(clk),
	.d(n211887));
   ms00f80 regtop_g_tmc_r_reg_10_ (.o(regtop_g_tmc_r[10]),
	.ck(clk),
	.d(n211886));
   ms00f80 regtop_g_tmc_r_reg_9_ (.o(regtop_g_tmc_r[9]),
	.ck(clk),
	.d(n211885));
   ms00f80 regtop_g_tmc_r_reg_8_ (.o(regtop_g_tmc_r[8]),
	.ck(clk),
	.d(n211884));
   ms00f80 regtop_g_tmc_r_reg_7_ (.o(regtop_g_tmc_r[7]),
	.ck(clk),
	.d(n211883));
   ms00f80 regtop_g_tmc_r_reg_6_ (.o(regtop_g_tmc_r[6]),
	.ck(clk),
	.d(n211882));
   ms00f80 regtop_g_tmc_r_reg_5_ (.o(regtop_g_tmc_r[5]),
	.ck(clk),
	.d(n211881));
   ms00f80 regtop_g_tmc_r_reg_4_ (.o(regtop_g_tmc_r[4]),
	.ck(clk),
	.d(n211880));
   ms00f80 regtop_g_tmc_r_reg_3_ (.o(regtop_g_tmc_r[3]),
	.ck(clk),
	.d(n211879));
   ms00f80 regtop_g_tmc_r_reg_2_ (.o(regtop_g_tmc_r[2]),
	.ck(clk),
	.d(n211878));
   ms00f80 regtop_g_tmc_r_reg_1_ (.o(regtop_g_tmc_r[1]),
	.ck(clk),
	.d(n211877));
   ms00f80 regtop_g_fpst01_r_reg (.o(regtop_g_fpst_r[0]),
	.ck(clk),
	.d(n211876));
   ms00f80 regtop_g_nfst23_r_reg (.o(regtop_g_nfst_r[22]),
	.ck(clk),
	.d(n186732));
   ms00f80 regtop_g_fbst08_r_reg (.o(regtop_g_fbst_r[7]),
	.ck(clk),
	.d(n186726));
   ms00f80 regtop_g_fbst07_r_reg (.o(regtop_g_fbst_r[6]),
	.ck(clk),
	.d(n186725));
   ms00f80 regtop_g_fbst06_r_reg (.o(regtop_g_fbst_r[5]),
	.ck(clk),
	.d(n186724));
   ms00f80 regtop_g_fbst05_r_reg (.o(regtop_g_fbst_r[4]),
	.ck(clk),
	.d(n186723));
   ms00f80 regtop_g_fbst04_r_reg (.o(regtop_g_fbst_r[3]),
	.ck(clk),
	.d(n186722));
   ms00f80 regtop_g_fbst02_r_reg (.o(regtop_g_fbst_r[1]),
	.ck(clk),
	.d(n186721));
   ms00f80 regtop_g_fbst01_r_reg (.o(regtop_g_fbst_r[0]),
	.ck(clk),
	.d(n186720));
   ms00f80 cntrltop_ctmg_ctpedet_c_bigpictdet_r_reg (.o(cntrltop_ctmg_ctpedet_c_bigpictdet_r),
	.ck(clk),
	.d(n186718));
   ms00f80 cntrltop_ctmg_ctpedet_c_tmg_ferr_pre_d1_r_reg (.o(cntrltop_ctmg_ctpedet_c_tmg_ferr_pre_d1_r),
	.ck(clk),
	.d(cntrltop_ctmg_ctpedet_c_tmg_ferr_pre));
   ms00f80 cntrltop_ctmg_ctpedet_c_tmg_ferr_hit_r_reg (.o(c_tmg_ferr_hit_r),
	.ck(clk),
	.d(cntrltop_ctmg_ctpedet_N22));
   ms00f80 regtop_g_tmg_ferr_hit_r_reg (.o(regtop_g_tmg_ferr_hit_r),
	.ck(clk),
	.d(c_tmg_ferr_hit_r));
   ms00f80 regtop_g_fbst10_r_reg (.o(regtop_g_fbst_r[9]),
	.ck(clk),
	.d(n186717));
   ms00f80 regtop_g_prev_efbst_r_reg (.o(regtop_g_prev_efbst_r),
	.ck(clk),
	.d(regtop_N1267));
   ms00f80 regtop_g_dsts_r_reg (.o(regtop_g_dsts_r),
	.ck(clk),
	.d(n186714));
   ms00f80 regtop_v1_dmareq8_n_reg (.o(v1_dmareq8_n),
	.ck(clk),
	.d(n245083));
   ms00f80 regtop_g_hclr_r_s_reg (.o(regtop_g_hclr_r_s),
	.ck(clk),
	.d(n186713));
   ms00f80 regtop_g_udb_cpu_r_reg_6_ (.o(regtop_g_udb_cpu_r[6]),
	.ck(clk),
	.d(n186699));
   ms00f80 regtop_g_udb_cpu_r_reg_5_ (.o(regtop_g_udb_cpu_r[5]),
	.ck(clk),
	.d(n186698));
   ms00f80 regtop_g_udb_cpu_r_reg_4_ (.o(regtop_g_udb_cpu_r[4]),
	.ck(clk),
	.d(n186697));
   ms00f80 regtop_g_udb_cpu_r_reg_3_ (.o(regtop_g_udb_cpu_r[3]),
	.ck(clk),
	.d(n186696));
   ms00f80 regtop_g_udb_cpu_r_reg_2_ (.o(regtop_g_udb_cpu_r[2]),
	.ck(clk),
	.d(n186695));
   ms00f80 regtop_g_udb_cpu_r_reg_1_ (.o(regtop_g_udb_cpu_r[1]),
	.ck(clk),
	.d(n186694));
   ms00f80 regtop_g_udb_cpu_r_reg_0_ (.o(regtop_g_udb_cpu_r[0]),
	.ck(clk),
	.d(n186693));
   ms00f80 regtop_g_adb_cpu_r_reg_6_ (.o(regtop_g_adb_cpu_r[6]),
	.ck(clk),
	.d(n186692));
   ms00f80 regtop_g_adb_cpu_r_reg_5_ (.o(regtop_g_adb_cpu_r[5]),
	.ck(clk),
	.d(n186691));
   ms00f80 regtop_g_adb_cpu_r_reg_4_ (.o(regtop_g_adb_cpu_r[4]),
	.ck(clk),
	.d(n186690));
   ms00f80 regtop_g_adb_cpu_r_reg_3_ (.o(regtop_g_adb_cpu_r[3]),
	.ck(clk),
	.d(n186689));
   ms00f80 regtop_g_adb_cpu_r_reg_2_ (.o(regtop_g_adb_cpu_r[2]),
	.ck(clk),
	.d(n186688));
   ms00f80 regtop_g_adb_cpu_r_reg_1_ (.o(regtop_g_adb_cpu_r[1]),
	.ck(clk),
	.d(n186687));
   ms00f80 regtop_g_adb_cpu_r_reg_0_ (.o(regtop_g_adb_cpu_r[0]),
	.ck(clk),
	.d(n186686));
   ms00f80 regtop_g_ispi_r_reg (.o(regtop_g_ispi_r),
	.ck(clk),
	.d(n186685));
   ms00f80 regtop_g_isph_r_reg (.o(regtop_g_isph_r),
	.ck(clk),
	.d(n186684));
   ms00f80 regtop_g_issw_r_reg (.o(regtop_g_issw_r),
	.ck(clk),
	.d(n186682));
   ms00f80 regtop_g_issr_r_reg (.o(regtop_g_issr_r),
	.ck(clk),
	.d(n186681));
   ms00f80 regtop_g_isfb_r_reg (.o(regtop_g_isfb_r),
	.ck(clk),
	.d(n186680));
   ms00f80 regtop_g_isfp_r_reg (.o(regtop_g_isfp_r),
	.ck(clk),
	.d(n186679));
   ms00f80 regtop_g_memr_ok_r_reg (.o(regtop_g_memr_ok_r),
	.ck(clk),
	.d(regtop_N1990));
   ms00f80 regtop_v1_hpb_wait_n_reg (.o(wbb_ack_o),
	.ck(clk),
	.d(n186678));
   ms00f80 regtop_v1_hdi00_d_reg_17_ (.o(regtop_v1_hdi00_d[17]),
	.ck(clk),
	.d(n245011));
   ms00f80 regtop_v1_hdi00_d_reg_16_ (.o(regtop_v1_hdi00_d[16]),
	.ck(clk),
	.d(n245010));
   ms00f80 regtop_v1_hdi00_d_reg_31_ (.o(regtop_v1_hdi00_d[31]),
	.ck(clk),
	.d(n245025));
   ms00f80 regtop_v1_hdi00_d_reg_30_ (.o(regtop_v1_hdi00_d[30]),
	.ck(clk),
	.d(n245024));
   ms00f80 regtop_v1_hdi00_d_reg_29_ (.o(regtop_v1_hdi00_d[29]),
	.ck(clk),
	.d(n245023));
   ms00f80 regtop_v1_hdi00_d_reg_28_ (.o(regtop_v1_hdi00_d[28]),
	.ck(clk),
	.d(n245022));
   ms00f80 regtop_v1_hdi00_d_reg_27_ (.o(regtop_v1_hdi00_d[27]),
	.ck(clk),
	.d(n245021));
   ms00f80 regtop_v1_hdi00_d_reg_26_ (.o(regtop_v1_hdi00_d[26]),
	.ck(clk),
	.d(n245020));
   ms00f80 regtop_v1_hdi00_d_reg_25_ (.o(regtop_v1_hdi00_d[25]),
	.ck(clk),
	.d(n245019));
   ms00f80 regtop_v1_hdi00_d_reg_24_ (.o(regtop_v1_hdi00_d[24]),
	.ck(clk),
	.d(n245018));
   ms00f80 regtop_v1_hdi00_d_reg_23_ (.o(regtop_v1_hdi00_d[23]),
	.ck(clk),
	.d(n245017));
   ms00f80 regtop_v1_hdi00_d_reg_22_ (.o(regtop_v1_hdi00_d[22]),
	.ck(clk),
	.d(n245016));
   ms00f80 regtop_v1_hdi00_d_reg_21_ (.o(regtop_v1_hdi00_d[21]),
	.ck(clk),
	.d(n245015));
   ms00f80 regtop_v1_hdi00_d_reg_20_ (.o(regtop_v1_hdi00_d[20]),
	.ck(clk),
	.d(n245014));
   ms00f80 regtop_v1_hdi00_d_reg_19_ (.o(regtop_v1_hdi00_d[19]),
	.ck(clk),
	.d(n245013));
   ms00f80 regtop_v1_hdi00_d_reg_18_ (.o(regtop_v1_hdi00_d[18]),
	.ck(clk),
	.d(n245012));
   ms00f80 regtop_v1_hdi00_d_reg_15_ (.o(regtop_v1_hdi00_d[15]),
	.ck(clk),
	.d(n245009));
   ms00f80 regtop_v1_hdi00_d_reg_14_ (.o(regtop_v1_hdi00_d[14]),
	.ck(clk),
	.d(n245008));
   ms00f80 regtop_v1_hdi00_d_reg_13_ (.o(regtop_v1_hdi00_d[13]),
	.ck(clk),
	.d(n245007));
   ms00f80 regtop_v1_hdi00_d_reg_12_ (.o(regtop_v1_hdi00_d[12]),
	.ck(clk),
	.d(n245006));
   ms00f80 regtop_v1_hdi00_d_reg_11_ (.o(regtop_v1_hdi00_d[11]),
	.ck(clk),
	.d(n245005));
   ms00f80 regtop_v1_hdi00_d_reg_10_ (.o(regtop_v1_hdi00_d[10]),
	.ck(clk),
	.d(n245004));
   ms00f80 regtop_v1_hdi00_d_reg_9_ (.o(regtop_v1_hdi00_d[9]),
	.ck(clk),
	.d(n245003));
   ms00f80 regtop_v1_hdi00_d_reg_8_ (.o(regtop_v1_hdi00_d[8]),
	.ck(clk),
	.d(n245002));
   ms00f80 regtop_v1_hdi00_d_reg_7_ (.o(regtop_v1_hdi00_d[7]),
	.ck(clk),
	.d(n245001));
   ms00f80 regtop_v1_hdi00_d_reg_6_ (.o(regtop_v1_hdi00_d[6]),
	.ck(clk),
	.d(n245000));
   ms00f80 regtop_v1_hdi00_d_reg_5_ (.o(regtop_v1_hdi00_d[5]),
	.ck(clk),
	.d(n244999));
   ms00f80 regtop_v1_hdi00_d_reg_4_ (.o(regtop_v1_hdi00_d[4]),
	.ck(clk),
	.d(n244998));
   ms00f80 regtop_v1_hdi00_d_reg_3_ (.o(regtop_v1_hdi00_d[3]),
	.ck(clk),
	.d(n244997));
   ms00f80 regtop_v1_hdi00_d_reg_2_ (.o(regtop_v1_hdi00_d[2]),
	.ck(clk),
	.d(n244996));
   ms00f80 regtop_v1_hdi00_d_reg_1_ (.o(regtop_v1_hdi00_d[1]),
	.ck(clk),
	.d(n244995));
   ms00f80 regtop_v1_hdi00_d_reg_0_ (.o(regtop_v1_hdi00_d[0]),
	.ck(clk),
	.d(n244994));
   ms00f80 regtop_v1_hdi00_a_reg_0_ (.o(regtop_v1_hdi00_a[0]),
	.ck(clk),
	.d(n244992));
   ms00f80 regtop_v1_hdi00_a_reg_1_ (.o(regtop_v1_hdi00_a[1]),
	.ck(clk),
	.d(n244991));
   ms00f80 regtop_v1_hdi00_a_reg_2_ (.o(regtop_v1_hdi00_a[2]),
	.ck(clk),
	.d(n244990));
   ms00f80 regtop_v1_hdi00_a_reg_3_ (.o(regtop_v1_hdi00_a[3]),
	.ck(clk),
	.d(n244989));
   ms00f80 regtop_v1_hdi00_a_reg_4_ (.o(regtop_v1_hdi00_a[4]),
	.ck(clk),
	.d(n244988));
   ms00f80 regtop_v1_hdi00_a_reg_5_ (.o(regtop_v1_hdi00_a[5]),
	.ck(clk),
	.d(n244987));
   ms00f80 regtop_v1_hdi00_we_reg (.o(regtop_v1_hdi00_we),
	.ck(clk),
	.d(n245026));
   ms00f80 regtop_v1_hdi00_bs_reg (.o(regtop_v1_hdi00_bs),
	.ck(clk),
	.d(n244986));
   ms00f80 regtop_g_rd_en_r_reg (.o(regtop_g_rd_en_r),
	.ck(clk),
	.d(regtop_N1991));
   ms00f80 regtop_g_rd_en2_r_reg (.o(regtop_g_rd_en2_r),
	.ck(clk),
	.d(regtop_g_rd_en_r));
   ms00f80 regtop_g_mem_rd2_r_reg_0_ (.o(regtop_g_mem_rd2_r[0]),
	.ck(clk),
	.d(regtop_N1993));
   ms00f80 regtop_g_mem_rd2_r_reg_1_ (.o(regtop_g_mem_rd2_r[1]),
	.ck(clk),
	.d(regtop_N1994));
   ms00f80 regtop_g_mem_rd2_r_reg_2_ (.o(regtop_g_mem_rd2_r[2]),
	.ck(clk),
	.d(regtop_N1995));
   ms00f80 regtop_g_mem_rd2_r_reg_3_ (.o(regtop_g_mem_rd2_r[3]),
	.ck(clk),
	.d(regtop_N1996));
   ms00f80 regtop_g_mem_rd2_r_reg_4_ (.o(regtop_g_mem_rd2_r[4]),
	.ck(clk),
	.d(regtop_N1997));
   ms00f80 regtop_g_mem_rd2_r_reg_5_ (.o(regtop_g_mem_rd2_r[5]),
	.ck(clk),
	.d(regtop_N1998));
   ms00f80 regtop_g_mem_rd2_r_reg_6_ (.o(regtop_g_mem_rd2_r[6]),
	.ck(clk),
	.d(regtop_N1999));
   ms00f80 regtop_g_mem_rd2_r_reg_7_ (.o(regtop_g_mem_rd2_r[7]),
	.ck(clk),
	.d(regtop_N2000));
   ms00f80 regtop_g_mem_rd2_r_reg_8_ (.o(regtop_g_mem_rd2_r[8]),
	.ck(clk),
	.d(regtop_N2001));
   ms00f80 regtop_g_mem_rd2_r_reg_9_ (.o(regtop_g_mem_rd2_r[9]),
	.ck(clk),
	.d(regtop_N2002));
   ms00f80 regtop_g_mem_rd2_r_reg_10_ (.o(regtop_g_mem_rd2_r[10]),
	.ck(clk),
	.d(regtop_N2003));
   ms00f80 regtop_g_mem_rd2_r_reg_11_ (.o(regtop_g_mem_rd2_r[11]),
	.ck(clk),
	.d(regtop_N2004));
   ms00f80 regtop_g_mem_rd2_r_reg_12_ (.o(regtop_g_mem_rd2_r[12]),
	.ck(clk),
	.d(regtop_N2005));
   ms00f80 regtop_g_mem_rd2_r_reg_13_ (.o(regtop_g_mem_rd2_r[13]),
	.ck(clk),
	.d(regtop_N2006));
   ms00f80 regtop_g_mem_rd2_r_reg_14_ (.o(regtop_g_mem_rd2_r[14]),
	.ck(clk),
	.d(regtop_N2007));
   ms00f80 regtop_g_mem_rd2_r_reg_15_ (.o(regtop_g_mem_rd2_r[15]),
	.ck(clk),
	.d(regtop_N2008));
   ms00f80 regtop_g_mem_rd2_r_reg_16_ (.o(regtop_g_mem_rd2_r[16]),
	.ck(clk),
	.d(regtop_N2009));
   ms00f80 regtop_g_mem_rd2_r_reg_17_ (.o(regtop_g_mem_rd2_r[17]),
	.ck(clk),
	.d(regtop_N2010));
   ms00f80 regtop_g_mem_rd2_r_reg_18_ (.o(regtop_g_mem_rd2_r[18]),
	.ck(clk),
	.d(regtop_N2011));
   ms00f80 regtop_g_mem_rd2_r_reg_19_ (.o(regtop_g_mem_rd2_r[19]),
	.ck(clk),
	.d(regtop_N2012));
   ms00f80 regtop_g_mem_rd2_r_reg_20_ (.o(regtop_g_mem_rd2_r[20]),
	.ck(clk),
	.d(regtop_N2013));
   ms00f80 regtop_g_mem_rd2_r_reg_21_ (.o(regtop_g_mem_rd2_r[21]),
	.ck(clk),
	.d(regtop_N2014));
   ms00f80 regtop_g_mem_rd2_r_reg_22_ (.o(regtop_g_mem_rd2_r[22]),
	.ck(clk),
	.d(regtop_N2015));
   ms00f80 regtop_g_mem_rd2_r_reg_23_ (.o(regtop_g_mem_rd2_r[23]),
	.ck(clk),
	.d(regtop_N2016));
   ms00f80 regtop_g_mem_rd2_r_reg_24_ (.o(regtop_g_mem_rd2_r[24]),
	.ck(clk),
	.d(regtop_N2017));
   ms00f80 regtop_g_mem_rd2_r_reg_25_ (.o(regtop_g_mem_rd2_r[25]),
	.ck(clk),
	.d(regtop_N2018));
   ms00f80 regtop_g_mem_rd2_r_reg_26_ (.o(regtop_g_mem_rd2_r[26]),
	.ck(clk),
	.d(regtop_N2019));
   ms00f80 regtop_g_mem_rd2_r_reg_27_ (.o(regtop_g_mem_rd2_r[27]),
	.ck(clk),
	.d(regtop_N2020));
   ms00f80 regtop_g_mem_rd2_r_reg_28_ (.o(regtop_g_mem_rd2_r[28]),
	.ck(clk),
	.d(regtop_N2021));
   ms00f80 regtop_g_mem_rd2_r_reg_29_ (.o(regtop_g_mem_rd2_r[29]),
	.ck(clk),
	.d(regtop_N2022));
   ms00f80 regtop_g_mem_rd2_r_reg_30_ (.o(regtop_g_mem_rd2_r[30]),
	.ck(clk),
	.d(regtop_N2023));
   ms00f80 regtop_g_mem_rd2_r_reg_31_ (.o(regtop_g_mem_rd2_r[31]),
	.ck(clk),
	.d(regtop_N2024));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__0_ (.o(regtop_dchdi_w1_hdi00[1536]),
	.ck(clk),
	.d(n186677));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__1_ (.o(regtop_dchdi_w1_hdi00[1537]),
	.ck(clk),
	.d(n186676));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__2_ (.o(regtop_dchdi_w1_hdi00[1538]),
	.ck(clk),
	.d(n186675));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__3_ (.o(regtop_dchdi_w1_hdi00[1539]),
	.ck(clk),
	.d(n186674));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__4_ (.o(regtop_dchdi_w1_hdi00[1540]),
	.ck(clk),
	.d(n186673));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__5_ (.o(regtop_dchdi_w1_hdi00[1541]),
	.ck(clk),
	.d(n186672));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__6_ (.o(regtop_dchdi_w1_hdi00[1542]),
	.ck(clk),
	.d(n186671));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__7_ (.o(regtop_dchdi_w1_hdi00[1543]),
	.ck(clk),
	.d(n186670));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__8_ (.o(regtop_dchdi_w1_hdi00[1544]),
	.ck(clk),
	.d(n186669));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__9_ (.o(regtop_dchdi_w1_hdi00[1545]),
	.ck(clk),
	.d(n186668));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__10_ (.o(regtop_dchdi_w1_hdi00[1546]),
	.ck(clk),
	.d(n186667));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__11_ (.o(regtop_dchdi_w1_hdi00[1547]),
	.ck(clk),
	.d(n186666));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__12_ (.o(regtop_dchdi_w1_hdi00[1548]),
	.ck(clk),
	.d(n186665));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__13_ (.o(regtop_dchdi_w1_hdi00[1549]),
	.ck(clk),
	.d(n186664));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__14_ (.o(regtop_dchdi_w1_hdi00[1550]),
	.ck(clk),
	.d(n186663));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__15_ (.o(regtop_dchdi_w1_hdi00[1551]),
	.ck(clk),
	.d(n186662));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__16_ (.o(regtop_dchdi_w1_hdi00[1552]),
	.ck(clk),
	.d(n186661));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__17_ (.o(regtop_dchdi_w1_hdi00[1553]),
	.ck(clk),
	.d(n186660));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__18_ (.o(regtop_dchdi_w1_hdi00[1554]),
	.ck(clk),
	.d(n186659));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__19_ (.o(regtop_dchdi_w1_hdi00[1555]),
	.ck(clk),
	.d(n186658));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__20_ (.o(regtop_dchdi_w1_hdi00[1556]),
	.ck(clk),
	.d(n186657));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__21_ (.o(regtop_dchdi_w1_hdi00[1557]),
	.ck(clk),
	.d(n186656));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__22_ (.o(regtop_dchdi_w1_hdi00[1558]),
	.ck(clk),
	.d(n186655));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__23_ (.o(regtop_dchdi_w1_hdi00[1559]),
	.ck(clk),
	.d(n186654));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__24_ (.o(regtop_dchdi_w1_hdi00[1560]),
	.ck(clk),
	.d(n186653));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__25_ (.o(regtop_dchdi_w1_hdi00[1561]),
	.ck(clk),
	.d(n186652));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__26_ (.o(regtop_dchdi_w1_hdi00[1562]),
	.ck(clk),
	.d(n186651));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__27_ (.o(regtop_dchdi_w1_hdi00[1563]),
	.ck(clk),
	.d(n186650));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__28_ (.o(regtop_dchdi_w1_hdi00[1564]),
	.ck(clk),
	.d(n186649));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__29_ (.o(regtop_dchdi_w1_hdi00[1565]),
	.ck(clk),
	.d(n186648));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__30_ (.o(regtop_dchdi_w1_hdi00[1566]),
	.ck(clk),
	.d(n186647));
   ms00f80 regtop_dchdi_w1_hdi00_reg_0__31_ (.o(regtop_dchdi_w1_hdi00[1567]),
	.ck(clk),
	.d(n186646));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__0_ (.o(regtop_dchdi_w1_hdi00[1568]),
	.ck(clk),
	.d(n186645));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__1_ (.o(regtop_dchdi_w1_hdi00[1569]),
	.ck(clk),
	.d(n186644));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__2_ (.o(regtop_dchdi_w1_hdi00[1570]),
	.ck(clk),
	.d(n186643));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__3_ (.o(regtop_dchdi_w1_hdi00[1571]),
	.ck(clk),
	.d(n186642));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__4_ (.o(regtop_dchdi_w1_hdi00[1572]),
	.ck(clk),
	.d(n186641));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__5_ (.o(regtop_dchdi_w1_hdi00[1573]),
	.ck(clk),
	.d(n186640));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__6_ (.o(regtop_dchdi_w1_hdi00[1574]),
	.ck(clk),
	.d(n186639));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__7_ (.o(regtop_dchdi_w1_hdi00[1575]),
	.ck(clk),
	.d(n186638));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__8_ (.o(regtop_dchdi_w1_hdi00[1576]),
	.ck(clk),
	.d(n186637));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__9_ (.o(regtop_dchdi_w1_hdi00[1577]),
	.ck(clk),
	.d(n186636));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__10_ (.o(regtop_dchdi_w1_hdi00[1578]),
	.ck(clk),
	.d(n186635));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__11_ (.o(regtop_dchdi_w1_hdi00[1579]),
	.ck(clk),
	.d(n186634));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__12_ (.o(regtop_dchdi_w1_hdi00[1580]),
	.ck(clk),
	.d(n186633));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__13_ (.o(regtop_dchdi_w1_hdi00[1581]),
	.ck(clk),
	.d(n186632));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__14_ (.o(regtop_dchdi_w1_hdi00[1582]),
	.ck(clk),
	.d(n186631));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__15_ (.o(regtop_dchdi_w1_hdi00[1583]),
	.ck(clk),
	.d(n186630));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__16_ (.o(regtop_dchdi_w1_hdi00[1584]),
	.ck(clk),
	.d(n186629));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__17_ (.o(regtop_dchdi_w1_hdi00[1585]),
	.ck(clk),
	.d(n186628));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__18_ (.o(regtop_dchdi_w1_hdi00[1586]),
	.ck(clk),
	.d(n186627));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__19_ (.o(regtop_dchdi_w1_hdi00[1587]),
	.ck(clk),
	.d(n186626));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__20_ (.o(regtop_dchdi_w1_hdi00[1588]),
	.ck(clk),
	.d(n186625));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__21_ (.o(regtop_dchdi_w1_hdi00[1589]),
	.ck(clk),
	.d(n186624));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__22_ (.o(regtop_dchdi_w1_hdi00[1590]),
	.ck(clk),
	.d(n186623));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__23_ (.o(regtop_dchdi_w1_hdi00[1591]),
	.ck(clk),
	.d(n186622));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__24_ (.o(regtop_dchdi_w1_hdi00[1592]),
	.ck(clk),
	.d(n186621));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__25_ (.o(regtop_dchdi_w1_hdi00[1593]),
	.ck(clk),
	.d(n186620));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__26_ (.o(regtop_dchdi_w1_hdi00[1594]),
	.ck(clk),
	.d(n186619));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__27_ (.o(regtop_dchdi_w1_hdi00[1595]),
	.ck(clk),
	.d(n186618));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__28_ (.o(regtop_dchdi_w1_hdi00[1596]),
	.ck(clk),
	.d(n186617));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__29_ (.o(regtop_dchdi_w1_hdi00[1597]),
	.ck(clk),
	.d(n186616));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__30_ (.o(regtop_dchdi_w1_hdi00[1598]),
	.ck(clk),
	.d(n186615));
   ms00f80 regtop_dchdi_w1_hdi00_reg_1__31_ (.o(regtop_dchdi_w1_hdi00[1599]),
	.ck(clk),
	.d(n186614));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__0_ (.o(regtop_dchdi_w1_hdi00[1600]),
	.ck(clk),
	.d(n186613));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__1_ (.o(regtop_dchdi_w1_hdi00[1601]),
	.ck(clk),
	.d(n186612));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__2_ (.o(regtop_dchdi_w1_hdi00[1602]),
	.ck(clk),
	.d(n186611));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__3_ (.o(regtop_dchdi_w1_hdi00[1603]),
	.ck(clk),
	.d(n186610));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__4_ (.o(regtop_dchdi_w1_hdi00[1604]),
	.ck(clk),
	.d(n186609));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__5_ (.o(regtop_dchdi_w1_hdi00[1605]),
	.ck(clk),
	.d(n186608));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__6_ (.o(regtop_dchdi_w1_hdi00[1606]),
	.ck(clk),
	.d(n186607));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__7_ (.o(regtop_dchdi_w1_hdi00[1607]),
	.ck(clk),
	.d(n186606));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__8_ (.o(regtop_dchdi_w1_hdi00[1608]),
	.ck(clk),
	.d(n186605));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__9_ (.o(regtop_dchdi_w1_hdi00[1609]),
	.ck(clk),
	.d(n186604));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__10_ (.o(regtop_dchdi_w1_hdi00[1610]),
	.ck(clk),
	.d(n186603));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__11_ (.o(regtop_dchdi_w1_hdi00[1611]),
	.ck(clk),
	.d(n186602));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__12_ (.o(regtop_dchdi_w1_hdi00[1612]),
	.ck(clk),
	.d(n186601));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__13_ (.o(regtop_dchdi_w1_hdi00[1613]),
	.ck(clk),
	.d(n186600));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__14_ (.o(regtop_dchdi_w1_hdi00[1614]),
	.ck(clk),
	.d(n186599));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__15_ (.o(regtop_dchdi_w1_hdi00[1615]),
	.ck(clk),
	.d(n186598));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__16_ (.o(regtop_dchdi_w1_hdi00[1616]),
	.ck(clk),
	.d(n186597));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__17_ (.o(regtop_dchdi_w1_hdi00[1617]),
	.ck(clk),
	.d(n186596));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__18_ (.o(regtop_dchdi_w1_hdi00[1618]),
	.ck(clk),
	.d(n186595));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__19_ (.o(regtop_dchdi_w1_hdi00[1619]),
	.ck(clk),
	.d(n186594));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__20_ (.o(regtop_dchdi_w1_hdi00[1620]),
	.ck(clk),
	.d(n186593));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__21_ (.o(regtop_dchdi_w1_hdi00[1621]),
	.ck(clk),
	.d(n186592));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__22_ (.o(regtop_dchdi_w1_hdi00[1622]),
	.ck(clk),
	.d(n186591));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__23_ (.o(regtop_dchdi_w1_hdi00[1623]),
	.ck(clk),
	.d(n186590));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__24_ (.o(regtop_dchdi_w1_hdi00[1624]),
	.ck(clk),
	.d(n186589));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__25_ (.o(regtop_dchdi_w1_hdi00[1625]),
	.ck(clk),
	.d(n186588));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__26_ (.o(regtop_dchdi_w1_hdi00[1626]),
	.ck(clk),
	.d(n186587));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__27_ (.o(regtop_dchdi_w1_hdi00[1627]),
	.ck(clk),
	.d(n186586));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__28_ (.o(regtop_dchdi_w1_hdi00[1628]),
	.ck(clk),
	.d(n186585));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__29_ (.o(regtop_dchdi_w1_hdi00[1629]),
	.ck(clk),
	.d(n186584));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__30_ (.o(regtop_dchdi_w1_hdi00[1630]),
	.ck(clk),
	.d(n186583));
   ms00f80 regtop_dchdi_w1_hdi00_reg_2__31_ (.o(regtop_dchdi_w1_hdi00[1631]),
	.ck(clk),
	.d(n186582));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__0_ (.o(regtop_dchdi_w1_hdi00[1632]),
	.ck(clk),
	.d(n186581));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__1_ (.o(regtop_dchdi_w1_hdi00[1633]),
	.ck(clk),
	.d(n186580));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__2_ (.o(regtop_dchdi_w1_hdi00[1634]),
	.ck(clk),
	.d(n186579));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__3_ (.o(regtop_dchdi_w1_hdi00[1635]),
	.ck(clk),
	.d(n186578));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__4_ (.o(regtop_dchdi_w1_hdi00[1636]),
	.ck(clk),
	.d(n186577));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__5_ (.o(regtop_dchdi_w1_hdi00[1637]),
	.ck(clk),
	.d(n186576));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__6_ (.o(regtop_dchdi_w1_hdi00[1638]),
	.ck(clk),
	.d(n186575));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__7_ (.o(regtop_dchdi_w1_hdi00[1639]),
	.ck(clk),
	.d(n186574));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__8_ (.o(regtop_dchdi_w1_hdi00[1640]),
	.ck(clk),
	.d(n186573));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__9_ (.o(regtop_dchdi_w1_hdi00[1641]),
	.ck(clk),
	.d(n186572));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__10_ (.o(regtop_dchdi_w1_hdi00[1642]),
	.ck(clk),
	.d(n186571));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__11_ (.o(regtop_dchdi_w1_hdi00[1643]),
	.ck(clk),
	.d(n186570));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__12_ (.o(regtop_dchdi_w1_hdi00[1644]),
	.ck(clk),
	.d(n186569));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__13_ (.o(regtop_dchdi_w1_hdi00[1645]),
	.ck(clk),
	.d(n186568));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__14_ (.o(regtop_dchdi_w1_hdi00[1646]),
	.ck(clk),
	.d(n186567));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__15_ (.o(regtop_dchdi_w1_hdi00[1647]),
	.ck(clk),
	.d(n186566));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__16_ (.o(regtop_dchdi_w1_hdi00[1648]),
	.ck(clk),
	.d(n186565));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__17_ (.o(regtop_dchdi_w1_hdi00[1649]),
	.ck(clk),
	.d(n186564));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__18_ (.o(regtop_dchdi_w1_hdi00[1650]),
	.ck(clk),
	.d(n186563));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__19_ (.o(regtop_dchdi_w1_hdi00[1651]),
	.ck(clk),
	.d(n186562));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__20_ (.o(regtop_dchdi_w1_hdi00[1652]),
	.ck(clk),
	.d(n186561));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__21_ (.o(regtop_dchdi_w1_hdi00[1653]),
	.ck(clk),
	.d(n186560));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__22_ (.o(regtop_dchdi_w1_hdi00[1654]),
	.ck(clk),
	.d(n186559));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__23_ (.o(regtop_dchdi_w1_hdi00[1655]),
	.ck(clk),
	.d(n186558));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__24_ (.o(regtop_dchdi_w1_hdi00[1656]),
	.ck(clk),
	.d(n186557));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__25_ (.o(regtop_dchdi_w1_hdi00[1657]),
	.ck(clk),
	.d(n186556));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__26_ (.o(regtop_dchdi_w1_hdi00[1658]),
	.ck(clk),
	.d(n186555));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__27_ (.o(regtop_dchdi_w1_hdi00[1659]),
	.ck(clk),
	.d(n186554));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__28_ (.o(regtop_dchdi_w1_hdi00[1660]),
	.ck(clk),
	.d(n186553));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__29_ (.o(regtop_dchdi_w1_hdi00[1661]),
	.ck(clk),
	.d(n186552));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__30_ (.o(regtop_dchdi_w1_hdi00[1662]),
	.ck(clk),
	.d(n186551));
   ms00f80 regtop_dchdi_w1_hdi00_reg_3__31_ (.o(regtop_dchdi_w1_hdi00[1663]),
	.ck(clk),
	.d(n186550));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__0_ (.o(regtop_dchdi_w1_hdi00[1664]),
	.ck(clk),
	.d(n186549));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__1_ (.o(regtop_dchdi_w1_hdi00[1665]),
	.ck(clk),
	.d(n186548));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__2_ (.o(regtop_dchdi_w1_hdi00[1666]),
	.ck(clk),
	.d(n186547));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__3_ (.o(regtop_dchdi_w1_hdi00[1667]),
	.ck(clk),
	.d(n186546));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__4_ (.o(regtop_dchdi_w1_hdi00[1668]),
	.ck(clk),
	.d(n186545));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__5_ (.o(regtop_dchdi_w1_hdi00[1669]),
	.ck(clk),
	.d(n186544));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__6_ (.o(regtop_dchdi_w1_hdi00[1670]),
	.ck(clk),
	.d(n186543));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__7_ (.o(regtop_dchdi_w1_hdi00[1671]),
	.ck(clk),
	.d(n186542));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__8_ (.o(regtop_dchdi_w1_hdi00[1672]),
	.ck(clk),
	.d(n186541));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__9_ (.o(regtop_dchdi_w1_hdi00[1673]),
	.ck(clk),
	.d(n186540));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__10_ (.o(regtop_dchdi_w1_hdi00[1674]),
	.ck(clk),
	.d(n186539));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__11_ (.o(regtop_dchdi_w1_hdi00[1675]),
	.ck(clk),
	.d(n186538));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__12_ (.o(regtop_dchdi_w1_hdi00[1676]),
	.ck(clk),
	.d(n186537));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__13_ (.o(regtop_dchdi_w1_hdi00[1677]),
	.ck(clk),
	.d(n186536));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__14_ (.o(regtop_dchdi_w1_hdi00[1678]),
	.ck(clk),
	.d(n186535));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__15_ (.o(regtop_dchdi_w1_hdi00[1679]),
	.ck(clk),
	.d(n186534));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__16_ (.o(regtop_dchdi_w1_hdi00[1680]),
	.ck(clk),
	.d(n186533));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__17_ (.o(regtop_dchdi_w1_hdi00[1681]),
	.ck(clk),
	.d(n186532));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__18_ (.o(regtop_dchdi_w1_hdi00[1682]),
	.ck(clk),
	.d(n186531));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__19_ (.o(regtop_dchdi_w1_hdi00[1683]),
	.ck(clk),
	.d(n186530));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__20_ (.o(regtop_dchdi_w1_hdi00[1684]),
	.ck(clk),
	.d(n186529));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__21_ (.o(regtop_dchdi_w1_hdi00[1685]),
	.ck(clk),
	.d(n186528));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__22_ (.o(regtop_dchdi_w1_hdi00[1686]),
	.ck(clk),
	.d(n186527));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__23_ (.o(regtop_dchdi_w1_hdi00[1687]),
	.ck(clk),
	.d(n186526));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__24_ (.o(regtop_dchdi_w1_hdi00[1688]),
	.ck(clk),
	.d(n186525));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__25_ (.o(regtop_dchdi_w1_hdi00[1689]),
	.ck(clk),
	.d(n186524));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__26_ (.o(regtop_dchdi_w1_hdi00[1690]),
	.ck(clk),
	.d(n186523));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__27_ (.o(regtop_dchdi_w1_hdi00[1691]),
	.ck(clk),
	.d(n186522));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__28_ (.o(regtop_dchdi_w1_hdi00[1692]),
	.ck(clk),
	.d(n186521));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__29_ (.o(regtop_dchdi_w1_hdi00[1693]),
	.ck(clk),
	.d(n186520));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__30_ (.o(regtop_dchdi_w1_hdi00[1694]),
	.ck(clk),
	.d(n186519));
   ms00f80 regtop_dchdi_w1_hdi00_reg_4__31_ (.o(regtop_dchdi_w1_hdi00[1695]),
	.ck(clk),
	.d(n186518));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__0_ (.o(regtop_dchdi_w1_hdi00[1696]),
	.ck(clk),
	.d(n186517));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__1_ (.o(regtop_dchdi_w1_hdi00[1697]),
	.ck(clk),
	.d(n186516));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__2_ (.o(regtop_dchdi_w1_hdi00[1698]),
	.ck(clk),
	.d(n186515));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__3_ (.o(regtop_dchdi_w1_hdi00[1699]),
	.ck(clk),
	.d(n186514));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__4_ (.o(regtop_dchdi_w1_hdi00[1700]),
	.ck(clk),
	.d(n186513));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__5_ (.o(regtop_dchdi_w1_hdi00[1701]),
	.ck(clk),
	.d(n186512));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__6_ (.o(regtop_dchdi_w1_hdi00[1702]),
	.ck(clk),
	.d(n186511));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__7_ (.o(regtop_dchdi_w1_hdi00[1703]),
	.ck(clk),
	.d(n186510));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__8_ (.o(regtop_dchdi_w1_hdi00[1704]),
	.ck(clk),
	.d(n186509));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__9_ (.o(regtop_dchdi_w1_hdi00[1705]),
	.ck(clk),
	.d(n186508));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__10_ (.o(regtop_dchdi_w1_hdi00[1706]),
	.ck(clk),
	.d(n186507));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__11_ (.o(regtop_dchdi_w1_hdi00[1707]),
	.ck(clk),
	.d(n186506));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__12_ (.o(regtop_dchdi_w1_hdi00[1708]),
	.ck(clk),
	.d(n186505));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__13_ (.o(regtop_dchdi_w1_hdi00[1709]),
	.ck(clk),
	.d(n186504));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__14_ (.o(regtop_dchdi_w1_hdi00[1710]),
	.ck(clk),
	.d(n186503));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__15_ (.o(regtop_dchdi_w1_hdi00[1711]),
	.ck(clk),
	.d(n186502));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__16_ (.o(regtop_dchdi_w1_hdi00[1712]),
	.ck(clk),
	.d(n186501));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__17_ (.o(regtop_dchdi_w1_hdi00[1713]),
	.ck(clk),
	.d(n186500));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__18_ (.o(regtop_dchdi_w1_hdi00[1714]),
	.ck(clk),
	.d(n186499));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__19_ (.o(regtop_dchdi_w1_hdi00[1715]),
	.ck(clk),
	.d(n186498));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__20_ (.o(regtop_dchdi_w1_hdi00[1716]),
	.ck(clk),
	.d(n186497));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__21_ (.o(regtop_dchdi_w1_hdi00[1717]),
	.ck(clk),
	.d(n186496));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__22_ (.o(regtop_dchdi_w1_hdi00[1718]),
	.ck(clk),
	.d(n186495));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__23_ (.o(regtop_dchdi_w1_hdi00[1719]),
	.ck(clk),
	.d(n186494));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__24_ (.o(regtop_dchdi_w1_hdi00[1720]),
	.ck(clk),
	.d(n186493));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__25_ (.o(regtop_dchdi_w1_hdi00[1721]),
	.ck(clk),
	.d(n186492));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__26_ (.o(regtop_dchdi_w1_hdi00[1722]),
	.ck(clk),
	.d(n186491));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__27_ (.o(regtop_dchdi_w1_hdi00[1723]),
	.ck(clk),
	.d(n186490));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__28_ (.o(regtop_dchdi_w1_hdi00[1724]),
	.ck(clk),
	.d(n186489));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__29_ (.o(regtop_dchdi_w1_hdi00[1725]),
	.ck(clk),
	.d(n186488));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__30_ (.o(regtop_dchdi_w1_hdi00[1726]),
	.ck(clk),
	.d(n186487));
   ms00f80 regtop_dchdi_w1_hdi00_reg_5__31_ (.o(regtop_dchdi_w1_hdi00[1727]),
	.ck(clk),
	.d(n186486));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__0_ (.o(regtop_dchdi_w1_hdi00[1728]),
	.ck(clk),
	.d(n186485));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__1_ (.o(regtop_dchdi_w1_hdi00[1729]),
	.ck(clk),
	.d(n186484));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__2_ (.o(regtop_dchdi_w1_hdi00[1730]),
	.ck(clk),
	.d(n186483));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__3_ (.o(regtop_dchdi_w1_hdi00[1731]),
	.ck(clk),
	.d(n186482));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__4_ (.o(regtop_dchdi_w1_hdi00[1732]),
	.ck(clk),
	.d(n186481));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__5_ (.o(regtop_dchdi_w1_hdi00[1733]),
	.ck(clk),
	.d(n186480));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__6_ (.o(regtop_dchdi_w1_hdi00[1734]),
	.ck(clk),
	.d(n186479));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__7_ (.o(regtop_dchdi_w1_hdi00[1735]),
	.ck(clk),
	.d(n186478));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__8_ (.o(regtop_dchdi_w1_hdi00[1736]),
	.ck(clk),
	.d(n186477));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__9_ (.o(regtop_dchdi_w1_hdi00[1737]),
	.ck(clk),
	.d(n186476));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__10_ (.o(regtop_dchdi_w1_hdi00[1738]),
	.ck(clk),
	.d(n186475));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__11_ (.o(regtop_dchdi_w1_hdi00[1739]),
	.ck(clk),
	.d(n186474));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__12_ (.o(regtop_dchdi_w1_hdi00[1740]),
	.ck(clk),
	.d(n186473));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__13_ (.o(regtop_dchdi_w1_hdi00[1741]),
	.ck(clk),
	.d(n186472));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__14_ (.o(regtop_dchdi_w1_hdi00[1742]),
	.ck(clk),
	.d(n186471));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__15_ (.o(regtop_dchdi_w1_hdi00[1743]),
	.ck(clk),
	.d(n186470));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__16_ (.o(regtop_dchdi_w1_hdi00[1744]),
	.ck(clk),
	.d(n186469));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__17_ (.o(regtop_dchdi_w1_hdi00[1745]),
	.ck(clk),
	.d(n186468));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__18_ (.o(regtop_dchdi_w1_hdi00[1746]),
	.ck(clk),
	.d(n186467));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__19_ (.o(regtop_dchdi_w1_hdi00[1747]),
	.ck(clk),
	.d(n186466));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__20_ (.o(regtop_dchdi_w1_hdi00[1748]),
	.ck(clk),
	.d(n186465));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__21_ (.o(regtop_dchdi_w1_hdi00[1749]),
	.ck(clk),
	.d(n186464));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__22_ (.o(regtop_dchdi_w1_hdi00[1750]),
	.ck(clk),
	.d(n186463));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__23_ (.o(regtop_dchdi_w1_hdi00[1751]),
	.ck(clk),
	.d(n186462));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__24_ (.o(regtop_dchdi_w1_hdi00[1752]),
	.ck(clk),
	.d(n186461));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__25_ (.o(regtop_dchdi_w1_hdi00[1753]),
	.ck(clk),
	.d(n186460));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__26_ (.o(regtop_dchdi_w1_hdi00[1754]),
	.ck(clk),
	.d(n186459));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__27_ (.o(regtop_dchdi_w1_hdi00[1755]),
	.ck(clk),
	.d(n186458));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__28_ (.o(regtop_dchdi_w1_hdi00[1756]),
	.ck(clk),
	.d(n186457));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__29_ (.o(regtop_dchdi_w1_hdi00[1757]),
	.ck(clk),
	.d(n186456));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__30_ (.o(regtop_dchdi_w1_hdi00[1758]),
	.ck(clk),
	.d(n186455));
   ms00f80 regtop_dchdi_w1_hdi00_reg_6__31_ (.o(regtop_dchdi_w1_hdi00[1759]),
	.ck(clk),
	.d(n186454));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__0_ (.o(regtop_dchdi_w1_hdi00[1760]),
	.ck(clk),
	.d(n186453));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__1_ (.o(regtop_dchdi_w1_hdi00[1761]),
	.ck(clk),
	.d(n186452));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__2_ (.o(regtop_dchdi_w1_hdi00[1762]),
	.ck(clk),
	.d(n186451));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__3_ (.o(regtop_dchdi_w1_hdi00[1763]),
	.ck(clk),
	.d(n186450));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__4_ (.o(regtop_dchdi_w1_hdi00[1764]),
	.ck(clk),
	.d(n186449));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__5_ (.o(regtop_dchdi_w1_hdi00[1765]),
	.ck(clk),
	.d(n186448));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__6_ (.o(regtop_dchdi_w1_hdi00[1766]),
	.ck(clk),
	.d(n186447));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__7_ (.o(regtop_dchdi_w1_hdi00[1767]),
	.ck(clk),
	.d(n186446));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__8_ (.o(regtop_dchdi_w1_hdi00[1768]),
	.ck(clk),
	.d(n186445));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__9_ (.o(regtop_dchdi_w1_hdi00[1769]),
	.ck(clk),
	.d(n186444));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__10_ (.o(regtop_dchdi_w1_hdi00[1770]),
	.ck(clk),
	.d(n186443));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__11_ (.o(regtop_dchdi_w1_hdi00[1771]),
	.ck(clk),
	.d(n186442));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__12_ (.o(regtop_dchdi_w1_hdi00[1772]),
	.ck(clk),
	.d(n186441));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__13_ (.o(regtop_dchdi_w1_hdi00[1773]),
	.ck(clk),
	.d(n186440));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__14_ (.o(regtop_dchdi_w1_hdi00[1774]),
	.ck(clk),
	.d(n186439));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__15_ (.o(regtop_dchdi_w1_hdi00[1775]),
	.ck(clk),
	.d(n186438));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__16_ (.o(regtop_dchdi_w1_hdi00[1776]),
	.ck(clk),
	.d(n186437));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__17_ (.o(regtop_dchdi_w1_hdi00[1777]),
	.ck(clk),
	.d(n186436));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__18_ (.o(regtop_dchdi_w1_hdi00[1778]),
	.ck(clk),
	.d(n186435));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__19_ (.o(regtop_dchdi_w1_hdi00[1779]),
	.ck(clk),
	.d(n186434));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__20_ (.o(regtop_dchdi_w1_hdi00[1780]),
	.ck(clk),
	.d(n186433));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__21_ (.o(regtop_dchdi_w1_hdi00[1781]),
	.ck(clk),
	.d(n186432));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__22_ (.o(regtop_dchdi_w1_hdi00[1782]),
	.ck(clk),
	.d(n186431));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__23_ (.o(regtop_dchdi_w1_hdi00[1783]),
	.ck(clk),
	.d(n186430));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__24_ (.o(regtop_dchdi_w1_hdi00[1784]),
	.ck(clk),
	.d(n186429));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__25_ (.o(regtop_dchdi_w1_hdi00[1785]),
	.ck(clk),
	.d(n186428));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__26_ (.o(regtop_dchdi_w1_hdi00[1786]),
	.ck(clk),
	.d(n186427));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__27_ (.o(regtop_dchdi_w1_hdi00[1787]),
	.ck(clk),
	.d(n186426));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__28_ (.o(regtop_dchdi_w1_hdi00[1788]),
	.ck(clk),
	.d(n186425));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__29_ (.o(regtop_dchdi_w1_hdi00[1789]),
	.ck(clk),
	.d(n186424));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__30_ (.o(regtop_dchdi_w1_hdi00[1790]),
	.ck(clk),
	.d(n186423));
   ms00f80 regtop_dchdi_w1_hdi00_reg_7__31_ (.o(regtop_dchdi_w1_hdi00[1791]),
	.ck(clk),
	.d(n186422));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__0_ (.o(regtop_dchdi_w1_hdi00[1792]),
	.ck(clk),
	.d(n186421));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__1_ (.o(regtop_dchdi_w1_hdi00[1793]),
	.ck(clk),
	.d(n186420));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__2_ (.o(regtop_dchdi_w1_hdi00[1794]),
	.ck(clk),
	.d(n186419));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__3_ (.o(regtop_dchdi_w1_hdi00[1795]),
	.ck(clk),
	.d(n186418));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__4_ (.o(regtop_dchdi_w1_hdi00[1796]),
	.ck(clk),
	.d(n186417));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__5_ (.o(regtop_dchdi_w1_hdi00[1797]),
	.ck(clk),
	.d(n186416));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__6_ (.o(regtop_dchdi_w1_hdi00[1798]),
	.ck(clk),
	.d(n186415));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__7_ (.o(regtop_dchdi_w1_hdi00[1799]),
	.ck(clk),
	.d(n186414));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__8_ (.o(regtop_dchdi_w1_hdi00[1800]),
	.ck(clk),
	.d(n186413));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__9_ (.o(regtop_dchdi_w1_hdi00[1801]),
	.ck(clk),
	.d(n186412));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__10_ (.o(regtop_dchdi_w1_hdi00[1802]),
	.ck(clk),
	.d(n186411));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__11_ (.o(regtop_dchdi_w1_hdi00[1803]),
	.ck(clk),
	.d(n186410));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__12_ (.o(regtop_dchdi_w1_hdi00[1804]),
	.ck(clk),
	.d(n186409));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__13_ (.o(regtop_dchdi_w1_hdi00[1805]),
	.ck(clk),
	.d(n186408));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__14_ (.o(regtop_dchdi_w1_hdi00[1806]),
	.ck(clk),
	.d(n186407));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__15_ (.o(regtop_dchdi_w1_hdi00[1807]),
	.ck(clk),
	.d(n186406));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__16_ (.o(regtop_dchdi_w1_hdi00[1808]),
	.ck(clk),
	.d(n186405));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__17_ (.o(regtop_dchdi_w1_hdi00[1809]),
	.ck(clk),
	.d(n186404));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__18_ (.o(regtop_dchdi_w1_hdi00[1810]),
	.ck(clk),
	.d(n186403));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__19_ (.o(regtop_dchdi_w1_hdi00[1811]),
	.ck(clk),
	.d(n186402));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__20_ (.o(regtop_dchdi_w1_hdi00[1812]),
	.ck(clk),
	.d(n186401));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__21_ (.o(regtop_dchdi_w1_hdi00[1813]),
	.ck(clk),
	.d(n186400));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__22_ (.o(regtop_dchdi_w1_hdi00[1814]),
	.ck(clk),
	.d(n186399));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__23_ (.o(regtop_dchdi_w1_hdi00[1815]),
	.ck(clk),
	.d(n186398));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__24_ (.o(regtop_dchdi_w1_hdi00[1816]),
	.ck(clk),
	.d(n186397));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__25_ (.o(regtop_dchdi_w1_hdi00[1817]),
	.ck(clk),
	.d(n186396));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__26_ (.o(regtop_dchdi_w1_hdi00[1818]),
	.ck(clk),
	.d(n186395));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__27_ (.o(regtop_dchdi_w1_hdi00[1819]),
	.ck(clk),
	.d(n186394));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__28_ (.o(regtop_dchdi_w1_hdi00[1820]),
	.ck(clk),
	.d(n186393));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__29_ (.o(regtop_dchdi_w1_hdi00[1821]),
	.ck(clk),
	.d(n186392));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__30_ (.o(regtop_dchdi_w1_hdi00[1822]),
	.ck(clk),
	.d(n186391));
   ms00f80 regtop_dchdi_w1_hdi00_reg_8__31_ (.o(regtop_dchdi_w1_hdi00[1823]),
	.ck(clk),
	.d(n186390));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__0_ (.o(regtop_dchdi_w1_hdi00[1824]),
	.ck(clk),
	.d(n186389));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__1_ (.o(regtop_dchdi_w1_hdi00[1825]),
	.ck(clk),
	.d(n186388));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__2_ (.o(regtop_dchdi_w1_hdi00[1826]),
	.ck(clk),
	.d(n186387));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__3_ (.o(regtop_dchdi_w1_hdi00[1827]),
	.ck(clk),
	.d(n186386));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__4_ (.o(regtop_dchdi_w1_hdi00[1828]),
	.ck(clk),
	.d(n186385));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__5_ (.o(regtop_dchdi_w1_hdi00[1829]),
	.ck(clk),
	.d(n186384));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__6_ (.o(regtop_dchdi_w1_hdi00[1830]),
	.ck(clk),
	.d(n186383));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__7_ (.o(regtop_dchdi_w1_hdi00[1831]),
	.ck(clk),
	.d(n186382));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__8_ (.o(regtop_dchdi_w1_hdi00[1832]),
	.ck(clk),
	.d(n186381));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__9_ (.o(regtop_dchdi_w1_hdi00[1833]),
	.ck(clk),
	.d(n186380));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__10_ (.o(regtop_dchdi_w1_hdi00[1834]),
	.ck(clk),
	.d(n186379));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__11_ (.o(regtop_dchdi_w1_hdi00[1835]),
	.ck(clk),
	.d(n186378));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__12_ (.o(regtop_dchdi_w1_hdi00[1836]),
	.ck(clk),
	.d(n186377));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__13_ (.o(regtop_dchdi_w1_hdi00[1837]),
	.ck(clk),
	.d(n186376));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__14_ (.o(regtop_dchdi_w1_hdi00[1838]),
	.ck(clk),
	.d(n186375));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__15_ (.o(regtop_dchdi_w1_hdi00[1839]),
	.ck(clk),
	.d(n186374));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__16_ (.o(regtop_dchdi_w1_hdi00[1840]),
	.ck(clk),
	.d(n186373));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__17_ (.o(regtop_dchdi_w1_hdi00[1841]),
	.ck(clk),
	.d(n186372));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__18_ (.o(regtop_dchdi_w1_hdi00[1842]),
	.ck(clk),
	.d(n186371));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__19_ (.o(regtop_dchdi_w1_hdi00[1843]),
	.ck(clk),
	.d(n186370));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__20_ (.o(regtop_dchdi_w1_hdi00[1844]),
	.ck(clk),
	.d(n186369));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__21_ (.o(regtop_dchdi_w1_hdi00[1845]),
	.ck(clk),
	.d(n186368));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__22_ (.o(regtop_dchdi_w1_hdi00[1846]),
	.ck(clk),
	.d(n186367));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__23_ (.o(regtop_dchdi_w1_hdi00[1847]),
	.ck(clk),
	.d(n186366));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__24_ (.o(regtop_dchdi_w1_hdi00[1848]),
	.ck(clk),
	.d(n186365));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__25_ (.o(regtop_dchdi_w1_hdi00[1849]),
	.ck(clk),
	.d(n186364));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__26_ (.o(regtop_dchdi_w1_hdi00[1850]),
	.ck(clk),
	.d(n186363));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__27_ (.o(regtop_dchdi_w1_hdi00[1851]),
	.ck(clk),
	.d(n186362));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__28_ (.o(regtop_dchdi_w1_hdi00[1852]),
	.ck(clk),
	.d(n186361));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__29_ (.o(regtop_dchdi_w1_hdi00[1853]),
	.ck(clk),
	.d(n186360));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__30_ (.o(regtop_dchdi_w1_hdi00[1854]),
	.ck(clk),
	.d(n186359));
   ms00f80 regtop_dchdi_w1_hdi00_reg_9__31_ (.o(regtop_dchdi_w1_hdi00[1855]),
	.ck(clk),
	.d(n186358));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__0_ (.o(regtop_dchdi_w1_hdi00[1856]),
	.ck(clk),
	.d(n186357));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__1_ (.o(regtop_dchdi_w1_hdi00[1857]),
	.ck(clk),
	.d(n186356));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__2_ (.o(regtop_dchdi_w1_hdi00[1858]),
	.ck(clk),
	.d(n186355));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__3_ (.o(regtop_dchdi_w1_hdi00[1859]),
	.ck(clk),
	.d(n186354));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__4_ (.o(regtop_dchdi_w1_hdi00[1860]),
	.ck(clk),
	.d(n186353));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__5_ (.o(regtop_dchdi_w1_hdi00[1861]),
	.ck(clk),
	.d(n186352));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__6_ (.o(regtop_dchdi_w1_hdi00[1862]),
	.ck(clk),
	.d(n186351));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__7_ (.o(regtop_dchdi_w1_hdi00[1863]),
	.ck(clk),
	.d(n186350));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__8_ (.o(regtop_dchdi_w1_hdi00[1864]),
	.ck(clk),
	.d(n186349));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__9_ (.o(regtop_dchdi_w1_hdi00[1865]),
	.ck(clk),
	.d(n186348));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__10_ (.o(regtop_dchdi_w1_hdi00[1866]),
	.ck(clk),
	.d(n186347));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__11_ (.o(regtop_dchdi_w1_hdi00[1867]),
	.ck(clk),
	.d(n186346));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__12_ (.o(regtop_dchdi_w1_hdi00[1868]),
	.ck(clk),
	.d(n186345));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__13_ (.o(regtop_dchdi_w1_hdi00[1869]),
	.ck(clk),
	.d(n186344));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__14_ (.o(regtop_dchdi_w1_hdi00[1870]),
	.ck(clk),
	.d(n186343));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__15_ (.o(regtop_dchdi_w1_hdi00[1871]),
	.ck(clk),
	.d(n186342));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__16_ (.o(regtop_dchdi_w1_hdi00[1872]),
	.ck(clk),
	.d(n186341));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__17_ (.o(regtop_dchdi_w1_hdi00[1873]),
	.ck(clk),
	.d(n186340));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__18_ (.o(regtop_dchdi_w1_hdi00[1874]),
	.ck(clk),
	.d(n186339));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__19_ (.o(regtop_dchdi_w1_hdi00[1875]),
	.ck(clk),
	.d(n186338));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__20_ (.o(regtop_dchdi_w1_hdi00[1876]),
	.ck(clk),
	.d(n186337));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__21_ (.o(regtop_dchdi_w1_hdi00[1877]),
	.ck(clk),
	.d(n186336));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__22_ (.o(regtop_dchdi_w1_hdi00[1878]),
	.ck(clk),
	.d(n186335));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__23_ (.o(regtop_dchdi_w1_hdi00[1879]),
	.ck(clk),
	.d(n186334));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__24_ (.o(regtop_dchdi_w1_hdi00[1880]),
	.ck(clk),
	.d(n186333));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__25_ (.o(regtop_dchdi_w1_hdi00[1881]),
	.ck(clk),
	.d(n186332));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__26_ (.o(regtop_dchdi_w1_hdi00[1882]),
	.ck(clk),
	.d(n186331));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__27_ (.o(regtop_dchdi_w1_hdi00[1883]),
	.ck(clk),
	.d(n186330));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__28_ (.o(regtop_dchdi_w1_hdi00[1884]),
	.ck(clk),
	.d(n186329));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__29_ (.o(regtop_dchdi_w1_hdi00[1885]),
	.ck(clk),
	.d(n186328));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__30_ (.o(regtop_dchdi_w1_hdi00[1886]),
	.ck(clk),
	.d(n186327));
   ms00f80 regtop_dchdi_w1_hdi00_reg_10__31_ (.o(regtop_dchdi_w1_hdi00[1887]),
	.ck(clk),
	.d(n186326));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__0_ (.o(regtop_dchdi_w1_hdi00[1888]),
	.ck(clk),
	.d(n186325));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__1_ (.o(regtop_dchdi_w1_hdi00[1889]),
	.ck(clk),
	.d(n186324));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__2_ (.o(regtop_dchdi_w1_hdi00[1890]),
	.ck(clk),
	.d(n186323));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__3_ (.o(regtop_dchdi_w1_hdi00[1891]),
	.ck(clk),
	.d(n186322));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__4_ (.o(regtop_dchdi_w1_hdi00[1892]),
	.ck(clk),
	.d(n186321));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__5_ (.o(regtop_dchdi_w1_hdi00[1893]),
	.ck(clk),
	.d(n186320));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__6_ (.o(regtop_dchdi_w1_hdi00[1894]),
	.ck(clk),
	.d(n186319));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__7_ (.o(regtop_dchdi_w1_hdi00[1895]),
	.ck(clk),
	.d(n186318));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__8_ (.o(regtop_dchdi_w1_hdi00[1896]),
	.ck(clk),
	.d(n186317));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__9_ (.o(regtop_dchdi_w1_hdi00[1897]),
	.ck(clk),
	.d(n186316));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__10_ (.o(regtop_dchdi_w1_hdi00[1898]),
	.ck(clk),
	.d(n186315));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__11_ (.o(regtop_dchdi_w1_hdi00[1899]),
	.ck(clk),
	.d(n186314));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__12_ (.o(regtop_dchdi_w1_hdi00[1900]),
	.ck(clk),
	.d(n186313));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__13_ (.o(regtop_dchdi_w1_hdi00[1901]),
	.ck(clk),
	.d(n186312));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__14_ (.o(regtop_dchdi_w1_hdi00[1902]),
	.ck(clk),
	.d(n186311));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__15_ (.o(regtop_dchdi_w1_hdi00[1903]),
	.ck(clk),
	.d(n186310));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__16_ (.o(regtop_dchdi_w1_hdi00[1904]),
	.ck(clk),
	.d(n186309));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__17_ (.o(regtop_dchdi_w1_hdi00[1905]),
	.ck(clk),
	.d(n186308));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__18_ (.o(regtop_dchdi_w1_hdi00[1906]),
	.ck(clk),
	.d(n186307));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__19_ (.o(regtop_dchdi_w1_hdi00[1907]),
	.ck(clk),
	.d(n186306));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__20_ (.o(regtop_dchdi_w1_hdi00[1908]),
	.ck(clk),
	.d(n186305));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__21_ (.o(regtop_dchdi_w1_hdi00[1909]),
	.ck(clk),
	.d(n186304));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__22_ (.o(regtop_dchdi_w1_hdi00[1910]),
	.ck(clk),
	.d(n186303));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__23_ (.o(regtop_dchdi_w1_hdi00[1911]),
	.ck(clk),
	.d(n186302));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__24_ (.o(regtop_dchdi_w1_hdi00[1912]),
	.ck(clk),
	.d(n186301));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__25_ (.o(regtop_dchdi_w1_hdi00[1913]),
	.ck(clk),
	.d(n186300));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__26_ (.o(regtop_dchdi_w1_hdi00[1914]),
	.ck(clk),
	.d(n186299));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__27_ (.o(regtop_dchdi_w1_hdi00[1915]),
	.ck(clk),
	.d(n186298));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__28_ (.o(regtop_dchdi_w1_hdi00[1916]),
	.ck(clk),
	.d(n186297));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__29_ (.o(regtop_dchdi_w1_hdi00[1917]),
	.ck(clk),
	.d(n186296));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__30_ (.o(regtop_dchdi_w1_hdi00[1918]),
	.ck(clk),
	.d(n186295));
   ms00f80 regtop_dchdi_w1_hdi00_reg_11__31_ (.o(regtop_dchdi_w1_hdi00[1919]),
	.ck(clk),
	.d(n186294));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__0_ (.o(regtop_dchdi_w1_hdi00[1920]),
	.ck(clk),
	.d(n186293));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__1_ (.o(regtop_dchdi_w1_hdi00[1921]),
	.ck(clk),
	.d(n186292));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__2_ (.o(regtop_dchdi_w1_hdi00[1922]),
	.ck(clk),
	.d(n186291));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__3_ (.o(regtop_dchdi_w1_hdi00[1923]),
	.ck(clk),
	.d(n186290));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__4_ (.o(regtop_dchdi_w1_hdi00[1924]),
	.ck(clk),
	.d(n186289));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__5_ (.o(regtop_dchdi_w1_hdi00[1925]),
	.ck(clk),
	.d(n186288));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__6_ (.o(regtop_dchdi_w1_hdi00[1926]),
	.ck(clk),
	.d(n186287));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__7_ (.o(regtop_dchdi_w1_hdi00[1927]),
	.ck(clk),
	.d(n186286));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__8_ (.o(regtop_dchdi_w1_hdi00[1928]),
	.ck(clk),
	.d(n186285));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__9_ (.o(regtop_dchdi_w1_hdi00[1929]),
	.ck(clk),
	.d(n186284));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__10_ (.o(regtop_dchdi_w1_hdi00[1930]),
	.ck(clk),
	.d(n186283));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__11_ (.o(regtop_dchdi_w1_hdi00[1931]),
	.ck(clk),
	.d(n186282));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__12_ (.o(regtop_dchdi_w1_hdi00[1932]),
	.ck(clk),
	.d(n186281));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__13_ (.o(regtop_dchdi_w1_hdi00[1933]),
	.ck(clk),
	.d(n186280));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__14_ (.o(regtop_dchdi_w1_hdi00[1934]),
	.ck(clk),
	.d(n186279));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__15_ (.o(regtop_dchdi_w1_hdi00[1935]),
	.ck(clk),
	.d(n186278));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__16_ (.o(regtop_dchdi_w1_hdi00[1936]),
	.ck(clk),
	.d(n186277));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__17_ (.o(regtop_dchdi_w1_hdi00[1937]),
	.ck(clk),
	.d(n186276));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__18_ (.o(regtop_dchdi_w1_hdi00[1938]),
	.ck(clk),
	.d(n186275));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__19_ (.o(regtop_dchdi_w1_hdi00[1939]),
	.ck(clk),
	.d(n186274));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__20_ (.o(regtop_dchdi_w1_hdi00[1940]),
	.ck(clk),
	.d(n186273));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__21_ (.o(regtop_dchdi_w1_hdi00[1941]),
	.ck(clk),
	.d(n186272));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__22_ (.o(regtop_dchdi_w1_hdi00[1942]),
	.ck(clk),
	.d(n186271));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__23_ (.o(regtop_dchdi_w1_hdi00[1943]),
	.ck(clk),
	.d(n186270));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__24_ (.o(regtop_dchdi_w1_hdi00[1944]),
	.ck(clk),
	.d(n186269));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__25_ (.o(regtop_dchdi_w1_hdi00[1945]),
	.ck(clk),
	.d(n186268));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__26_ (.o(regtop_dchdi_w1_hdi00[1946]),
	.ck(clk),
	.d(n186267));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__27_ (.o(regtop_dchdi_w1_hdi00[1947]),
	.ck(clk),
	.d(n186266));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__28_ (.o(regtop_dchdi_w1_hdi00[1948]),
	.ck(clk),
	.d(n186265));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__29_ (.o(regtop_dchdi_w1_hdi00[1949]),
	.ck(clk),
	.d(n186264));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__30_ (.o(regtop_dchdi_w1_hdi00[1950]),
	.ck(clk),
	.d(n186263));
   ms00f80 regtop_dchdi_w1_hdi00_reg_12__31_ (.o(regtop_dchdi_w1_hdi00[1951]),
	.ck(clk),
	.d(n186262));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__0_ (.o(regtop_dchdi_w1_hdi00[1952]),
	.ck(clk),
	.d(n186261));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__1_ (.o(regtop_dchdi_w1_hdi00[1953]),
	.ck(clk),
	.d(n186260));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__2_ (.o(regtop_dchdi_w1_hdi00[1954]),
	.ck(clk),
	.d(n186259));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__3_ (.o(regtop_dchdi_w1_hdi00[1955]),
	.ck(clk),
	.d(n186258));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__4_ (.o(regtop_dchdi_w1_hdi00[1956]),
	.ck(clk),
	.d(n186257));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__5_ (.o(regtop_dchdi_w1_hdi00[1957]),
	.ck(clk),
	.d(n186256));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__6_ (.o(regtop_dchdi_w1_hdi00[1958]),
	.ck(clk),
	.d(n186255));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__7_ (.o(regtop_dchdi_w1_hdi00[1959]),
	.ck(clk),
	.d(n186254));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__8_ (.o(regtop_dchdi_w1_hdi00[1960]),
	.ck(clk),
	.d(n186253));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__9_ (.o(regtop_dchdi_w1_hdi00[1961]),
	.ck(clk),
	.d(n186252));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__10_ (.o(regtop_dchdi_w1_hdi00[1962]),
	.ck(clk),
	.d(n186251));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__11_ (.o(regtop_dchdi_w1_hdi00[1963]),
	.ck(clk),
	.d(n186250));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__12_ (.o(regtop_dchdi_w1_hdi00[1964]),
	.ck(clk),
	.d(n186249));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__13_ (.o(regtop_dchdi_w1_hdi00[1965]),
	.ck(clk),
	.d(n186248));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__14_ (.o(regtop_dchdi_w1_hdi00[1966]),
	.ck(clk),
	.d(n186247));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__15_ (.o(regtop_dchdi_w1_hdi00[1967]),
	.ck(clk),
	.d(n186246));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__16_ (.o(regtop_dchdi_w1_hdi00[1968]),
	.ck(clk),
	.d(n186245));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__17_ (.o(regtop_dchdi_w1_hdi00[1969]),
	.ck(clk),
	.d(n186244));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__18_ (.o(regtop_dchdi_w1_hdi00[1970]),
	.ck(clk),
	.d(n186243));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__19_ (.o(regtop_dchdi_w1_hdi00[1971]),
	.ck(clk),
	.d(n186242));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__20_ (.o(regtop_dchdi_w1_hdi00[1972]),
	.ck(clk),
	.d(n186241));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__21_ (.o(regtop_dchdi_w1_hdi00[1973]),
	.ck(clk),
	.d(n186240));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__22_ (.o(regtop_dchdi_w1_hdi00[1974]),
	.ck(clk),
	.d(n186239));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__23_ (.o(regtop_dchdi_w1_hdi00[1975]),
	.ck(clk),
	.d(n186238));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__24_ (.o(regtop_dchdi_w1_hdi00[1976]),
	.ck(clk),
	.d(n186237));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__25_ (.o(regtop_dchdi_w1_hdi00[1977]),
	.ck(clk),
	.d(n186236));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__26_ (.o(regtop_dchdi_w1_hdi00[1978]),
	.ck(clk),
	.d(n186235));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__27_ (.o(regtop_dchdi_w1_hdi00[1979]),
	.ck(clk),
	.d(n186234));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__28_ (.o(regtop_dchdi_w1_hdi00[1980]),
	.ck(clk),
	.d(n186233));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__29_ (.o(regtop_dchdi_w1_hdi00[1981]),
	.ck(clk),
	.d(n186232));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__30_ (.o(regtop_dchdi_w1_hdi00[1982]),
	.ck(clk),
	.d(n186231));
   ms00f80 regtop_dchdi_w1_hdi00_reg_13__31_ (.o(regtop_dchdi_w1_hdi00[1983]),
	.ck(clk),
	.d(n186230));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__0_ (.o(regtop_dchdi_w1_hdi00[1984]),
	.ck(clk),
	.d(n186229));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__1_ (.o(regtop_dchdi_w1_hdi00[1985]),
	.ck(clk),
	.d(n186228));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__2_ (.o(regtop_dchdi_w1_hdi00[1986]),
	.ck(clk),
	.d(n186227));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__3_ (.o(regtop_dchdi_w1_hdi00[1987]),
	.ck(clk),
	.d(n186226));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__4_ (.o(regtop_dchdi_w1_hdi00[1988]),
	.ck(clk),
	.d(n186225));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__5_ (.o(regtop_dchdi_w1_hdi00[1989]),
	.ck(clk),
	.d(n186224));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__6_ (.o(regtop_dchdi_w1_hdi00[1990]),
	.ck(clk),
	.d(n186223));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__7_ (.o(regtop_dchdi_w1_hdi00[1991]),
	.ck(clk),
	.d(n186222));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__8_ (.o(regtop_dchdi_w1_hdi00[1992]),
	.ck(clk),
	.d(n186221));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__9_ (.o(regtop_dchdi_w1_hdi00[1993]),
	.ck(clk),
	.d(n186220));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__10_ (.o(regtop_dchdi_w1_hdi00[1994]),
	.ck(clk),
	.d(n186219));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__11_ (.o(regtop_dchdi_w1_hdi00[1995]),
	.ck(clk),
	.d(n186218));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__12_ (.o(regtop_dchdi_w1_hdi00[1996]),
	.ck(clk),
	.d(n186217));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__13_ (.o(regtop_dchdi_w1_hdi00[1997]),
	.ck(clk),
	.d(n186216));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__14_ (.o(regtop_dchdi_w1_hdi00[1998]),
	.ck(clk),
	.d(n186215));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__15_ (.o(regtop_dchdi_w1_hdi00[1999]),
	.ck(clk),
	.d(n186214));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__16_ (.o(regtop_dchdi_w1_hdi00[2000]),
	.ck(clk),
	.d(n186213));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__17_ (.o(regtop_dchdi_w1_hdi00[2001]),
	.ck(clk),
	.d(n186212));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__18_ (.o(regtop_dchdi_w1_hdi00[2002]),
	.ck(clk),
	.d(n186211));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__19_ (.o(regtop_dchdi_w1_hdi00[2003]),
	.ck(clk),
	.d(n186210));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__20_ (.o(regtop_dchdi_w1_hdi00[2004]),
	.ck(clk),
	.d(n186209));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__21_ (.o(regtop_dchdi_w1_hdi00[2005]),
	.ck(clk),
	.d(n186208));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__22_ (.o(regtop_dchdi_w1_hdi00[2006]),
	.ck(clk),
	.d(n186207));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__23_ (.o(regtop_dchdi_w1_hdi00[2007]),
	.ck(clk),
	.d(n186206));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__24_ (.o(regtop_dchdi_w1_hdi00[2008]),
	.ck(clk),
	.d(n186205));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__25_ (.o(regtop_dchdi_w1_hdi00[2009]),
	.ck(clk),
	.d(n186204));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__26_ (.o(regtop_dchdi_w1_hdi00[2010]),
	.ck(clk),
	.d(n186203));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__27_ (.o(regtop_dchdi_w1_hdi00[2011]),
	.ck(clk),
	.d(n186202));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__28_ (.o(regtop_dchdi_w1_hdi00[2012]),
	.ck(clk),
	.d(n186201));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__29_ (.o(regtop_dchdi_w1_hdi00[2013]),
	.ck(clk),
	.d(n186200));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__30_ (.o(regtop_dchdi_w1_hdi00[2014]),
	.ck(clk),
	.d(n186199));
   ms00f80 regtop_dchdi_w1_hdi00_reg_14__31_ (.o(regtop_dchdi_w1_hdi00[2015]),
	.ck(clk),
	.d(n186198));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__0_ (.o(regtop_dchdi_w1_hdi00[2016]),
	.ck(clk),
	.d(n186197));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__1_ (.o(regtop_dchdi_w1_hdi00[2017]),
	.ck(clk),
	.d(n186196));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__2_ (.o(regtop_dchdi_w1_hdi00[2018]),
	.ck(clk),
	.d(n186195));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__3_ (.o(regtop_dchdi_w1_hdi00[2019]),
	.ck(clk),
	.d(n186194));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__4_ (.o(regtop_dchdi_w1_hdi00[2020]),
	.ck(clk),
	.d(n186193));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__5_ (.o(regtop_dchdi_w1_hdi00[2021]),
	.ck(clk),
	.d(n186192));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__6_ (.o(regtop_dchdi_w1_hdi00[2022]),
	.ck(clk),
	.d(n186191));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__7_ (.o(regtop_dchdi_w1_hdi00[2023]),
	.ck(clk),
	.d(n186190));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__8_ (.o(regtop_dchdi_w1_hdi00[2024]),
	.ck(clk),
	.d(n186189));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__9_ (.o(regtop_dchdi_w1_hdi00[2025]),
	.ck(clk),
	.d(n186188));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__10_ (.o(regtop_dchdi_w1_hdi00[2026]),
	.ck(clk),
	.d(n186187));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__11_ (.o(regtop_dchdi_w1_hdi00[2027]),
	.ck(clk),
	.d(n186186));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__12_ (.o(regtop_dchdi_w1_hdi00[2028]),
	.ck(clk),
	.d(n186185));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__13_ (.o(regtop_dchdi_w1_hdi00[2029]),
	.ck(clk),
	.d(n186184));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__14_ (.o(regtop_dchdi_w1_hdi00[2030]),
	.ck(clk),
	.d(n186183));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__15_ (.o(regtop_dchdi_w1_hdi00[2031]),
	.ck(clk),
	.d(n186182));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__16_ (.o(regtop_dchdi_w1_hdi00[2032]),
	.ck(clk),
	.d(n186181));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__17_ (.o(regtop_dchdi_w1_hdi00[2033]),
	.ck(clk),
	.d(n186180));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__18_ (.o(regtop_dchdi_w1_hdi00[2034]),
	.ck(clk),
	.d(n186179));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__19_ (.o(regtop_dchdi_w1_hdi00[2035]),
	.ck(clk),
	.d(n186178));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__20_ (.o(regtop_dchdi_w1_hdi00[2036]),
	.ck(clk),
	.d(n186177));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__21_ (.o(regtop_dchdi_w1_hdi00[2037]),
	.ck(clk),
	.d(n186176));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__22_ (.o(regtop_dchdi_w1_hdi00[2038]),
	.ck(clk),
	.d(n186175));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__23_ (.o(regtop_dchdi_w1_hdi00[2039]),
	.ck(clk),
	.d(n186174));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__24_ (.o(regtop_dchdi_w1_hdi00[2040]),
	.ck(clk),
	.d(n186173));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__25_ (.o(regtop_dchdi_w1_hdi00[2041]),
	.ck(clk),
	.d(n186172));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__26_ (.o(regtop_dchdi_w1_hdi00[2042]),
	.ck(clk),
	.d(n186171));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__27_ (.o(regtop_dchdi_w1_hdi00[2043]),
	.ck(clk),
	.d(n186170));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__28_ (.o(regtop_dchdi_w1_hdi00[2044]),
	.ck(clk),
	.d(n186169));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__29_ (.o(regtop_dchdi_w1_hdi00[2045]),
	.ck(clk),
	.d(n186168));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__30_ (.o(regtop_dchdi_w1_hdi00[2046]),
	.ck(clk),
	.d(n186167));
   ms00f80 regtop_dchdi_w1_hdi00_reg_15__31_ (.o(regtop_dchdi_w1_hdi00[2047]),
	.ck(clk),
	.d(n186166));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__0_ (.o(regtop_dchdi_w1_hdi00[1024]),
	.ck(clk),
	.d(n186165));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__1_ (.o(regtop_dchdi_w1_hdi00[1025]),
	.ck(clk),
	.d(n186164));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__2_ (.o(regtop_dchdi_w1_hdi00[1026]),
	.ck(clk),
	.d(n186163));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__3_ (.o(regtop_dchdi_w1_hdi00[1027]),
	.ck(clk),
	.d(n186162));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__4_ (.o(regtop_dchdi_w1_hdi00[1028]),
	.ck(clk),
	.d(n186161));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__5_ (.o(regtop_dchdi_w1_hdi00[1029]),
	.ck(clk),
	.d(n186160));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__6_ (.o(regtop_dchdi_w1_hdi00[1030]),
	.ck(clk),
	.d(n186159));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__7_ (.o(regtop_dchdi_w1_hdi00[1031]),
	.ck(clk),
	.d(n186158));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__8_ (.o(regtop_dchdi_w1_hdi00[1032]),
	.ck(clk),
	.d(n186157));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__9_ (.o(regtop_dchdi_w1_hdi00[1033]),
	.ck(clk),
	.d(n186156));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__10_ (.o(regtop_dchdi_w1_hdi00[1034]),
	.ck(clk),
	.d(n186155));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__11_ (.o(regtop_dchdi_w1_hdi00[1035]),
	.ck(clk),
	.d(n186154));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__12_ (.o(regtop_dchdi_w1_hdi00[1036]),
	.ck(clk),
	.d(n186153));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__13_ (.o(regtop_dchdi_w1_hdi00[1037]),
	.ck(clk),
	.d(n186152));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__14_ (.o(regtop_dchdi_w1_hdi00[1038]),
	.ck(clk),
	.d(n186151));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__15_ (.o(regtop_dchdi_w1_hdi00[1039]),
	.ck(clk),
	.d(n186150));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__16_ (.o(regtop_dchdi_w1_hdi00[1040]),
	.ck(clk),
	.d(n186149));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__17_ (.o(regtop_dchdi_w1_hdi00[1041]),
	.ck(clk),
	.d(n186148));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__18_ (.o(regtop_dchdi_w1_hdi00[1042]),
	.ck(clk),
	.d(n186147));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__19_ (.o(regtop_dchdi_w1_hdi00[1043]),
	.ck(clk),
	.d(n186146));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__20_ (.o(regtop_dchdi_w1_hdi00[1044]),
	.ck(clk),
	.d(n186145));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__21_ (.o(regtop_dchdi_w1_hdi00[1045]),
	.ck(clk),
	.d(n186144));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__22_ (.o(regtop_dchdi_w1_hdi00[1046]),
	.ck(clk),
	.d(n186143));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__23_ (.o(regtop_dchdi_w1_hdi00[1047]),
	.ck(clk),
	.d(n186142));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__24_ (.o(regtop_dchdi_w1_hdi00[1048]),
	.ck(clk),
	.d(n186141));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__25_ (.o(regtop_dchdi_w1_hdi00[1049]),
	.ck(clk),
	.d(n186140));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__26_ (.o(regtop_dchdi_w1_hdi00[1050]),
	.ck(clk),
	.d(n186139));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__27_ (.o(regtop_dchdi_w1_hdi00[1051]),
	.ck(clk),
	.d(n186138));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__28_ (.o(regtop_dchdi_w1_hdi00[1052]),
	.ck(clk),
	.d(n186137));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__29_ (.o(regtop_dchdi_w1_hdi00[1053]),
	.ck(clk),
	.d(n186136));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__30_ (.o(regtop_dchdi_w1_hdi00[1054]),
	.ck(clk),
	.d(n186135));
   ms00f80 regtop_dchdi_w1_hdi00_reg_16__31_ (.o(regtop_dchdi_w1_hdi00[1055]),
	.ck(clk),
	.d(n186134));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__0_ (.o(regtop_dchdi_w1_hdi00[1056]),
	.ck(clk),
	.d(n186133));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__1_ (.o(regtop_dchdi_w1_hdi00[1057]),
	.ck(clk),
	.d(n186132));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__2_ (.o(regtop_dchdi_w1_hdi00[1058]),
	.ck(clk),
	.d(n186131));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__3_ (.o(regtop_dchdi_w1_hdi00[1059]),
	.ck(clk),
	.d(n186130));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__4_ (.o(regtop_dchdi_w1_hdi00[1060]),
	.ck(clk),
	.d(n186129));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__5_ (.o(regtop_dchdi_w1_hdi00[1061]),
	.ck(clk),
	.d(n186128));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__6_ (.o(regtop_dchdi_w1_hdi00[1062]),
	.ck(clk),
	.d(n186127));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__7_ (.o(regtop_dchdi_w1_hdi00[1063]),
	.ck(clk),
	.d(n186126));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__8_ (.o(regtop_dchdi_w1_hdi00[1064]),
	.ck(clk),
	.d(n186125));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__9_ (.o(regtop_dchdi_w1_hdi00[1065]),
	.ck(clk),
	.d(n186124));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__10_ (.o(regtop_dchdi_w1_hdi00[1066]),
	.ck(clk),
	.d(n186123));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__11_ (.o(regtop_dchdi_w1_hdi00[1067]),
	.ck(clk),
	.d(n186122));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__12_ (.o(regtop_dchdi_w1_hdi00[1068]),
	.ck(clk),
	.d(n186121));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__13_ (.o(regtop_dchdi_w1_hdi00[1069]),
	.ck(clk),
	.d(n186120));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__14_ (.o(regtop_dchdi_w1_hdi00[1070]),
	.ck(clk),
	.d(n186119));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__15_ (.o(regtop_dchdi_w1_hdi00[1071]),
	.ck(clk),
	.d(n186118));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__16_ (.o(regtop_dchdi_w1_hdi00[1072]),
	.ck(clk),
	.d(n186117));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__17_ (.o(regtop_dchdi_w1_hdi00[1073]),
	.ck(clk),
	.d(n186116));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__18_ (.o(regtop_dchdi_w1_hdi00[1074]),
	.ck(clk),
	.d(n186115));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__19_ (.o(regtop_dchdi_w1_hdi00[1075]),
	.ck(clk),
	.d(n186114));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__20_ (.o(regtop_dchdi_w1_hdi00[1076]),
	.ck(clk),
	.d(n186113));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__21_ (.o(regtop_dchdi_w1_hdi00[1077]),
	.ck(clk),
	.d(n186112));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__22_ (.o(regtop_dchdi_w1_hdi00[1078]),
	.ck(clk),
	.d(n186111));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__23_ (.o(regtop_dchdi_w1_hdi00[1079]),
	.ck(clk),
	.d(n186110));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__24_ (.o(regtop_dchdi_w1_hdi00[1080]),
	.ck(clk),
	.d(n186109));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__25_ (.o(regtop_dchdi_w1_hdi00[1081]),
	.ck(clk),
	.d(n186108));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__26_ (.o(regtop_dchdi_w1_hdi00[1082]),
	.ck(clk),
	.d(n186107));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__27_ (.o(regtop_dchdi_w1_hdi00[1083]),
	.ck(clk),
	.d(n186106));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__28_ (.o(regtop_dchdi_w1_hdi00[1084]),
	.ck(clk),
	.d(n186105));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__29_ (.o(regtop_dchdi_w1_hdi00[1085]),
	.ck(clk),
	.d(n186104));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__30_ (.o(regtop_dchdi_w1_hdi00[1086]),
	.ck(clk),
	.d(n186103));
   ms00f80 regtop_dchdi_w1_hdi00_reg_17__31_ (.o(regtop_dchdi_w1_hdi00[1087]),
	.ck(clk),
	.d(n186102));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__0_ (.o(regtop_dchdi_w1_hdi00[1088]),
	.ck(clk),
	.d(n186101));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__1_ (.o(regtop_dchdi_w1_hdi00[1089]),
	.ck(clk),
	.d(n186100));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__2_ (.o(regtop_dchdi_w1_hdi00[1090]),
	.ck(clk),
	.d(n186099));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__3_ (.o(regtop_dchdi_w1_hdi00[1091]),
	.ck(clk),
	.d(n186098));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__4_ (.o(regtop_dchdi_w1_hdi00[1092]),
	.ck(clk),
	.d(n186097));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__5_ (.o(regtop_dchdi_w1_hdi00[1093]),
	.ck(clk),
	.d(n186096));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__6_ (.o(regtop_dchdi_w1_hdi00[1094]),
	.ck(clk),
	.d(n186095));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__7_ (.o(regtop_dchdi_w1_hdi00[1095]),
	.ck(clk),
	.d(n186094));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__8_ (.o(regtop_dchdi_w1_hdi00[1096]),
	.ck(clk),
	.d(n186093));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__9_ (.o(regtop_dchdi_w1_hdi00[1097]),
	.ck(clk),
	.d(n186092));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__10_ (.o(regtop_dchdi_w1_hdi00[1098]),
	.ck(clk),
	.d(n186091));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__11_ (.o(regtop_dchdi_w1_hdi00[1099]),
	.ck(clk),
	.d(n186090));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__12_ (.o(regtop_dchdi_w1_hdi00[1100]),
	.ck(clk),
	.d(n186089));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__13_ (.o(regtop_dchdi_w1_hdi00[1101]),
	.ck(clk),
	.d(n186088));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__14_ (.o(regtop_dchdi_w1_hdi00[1102]),
	.ck(clk),
	.d(n186087));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__15_ (.o(regtop_dchdi_w1_hdi00[1103]),
	.ck(clk),
	.d(n186086));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__16_ (.o(regtop_dchdi_w1_hdi00[1104]),
	.ck(clk),
	.d(n186085));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__17_ (.o(regtop_dchdi_w1_hdi00[1105]),
	.ck(clk),
	.d(n186084));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__18_ (.o(regtop_dchdi_w1_hdi00[1106]),
	.ck(clk),
	.d(n186083));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__19_ (.o(regtop_dchdi_w1_hdi00[1107]),
	.ck(clk),
	.d(n186082));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__20_ (.o(regtop_dchdi_w1_hdi00[1108]),
	.ck(clk),
	.d(n186081));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__21_ (.o(regtop_dchdi_w1_hdi00[1109]),
	.ck(clk),
	.d(n186080));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__22_ (.o(regtop_dchdi_w1_hdi00[1110]),
	.ck(clk),
	.d(n186079));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__23_ (.o(regtop_dchdi_w1_hdi00[1111]),
	.ck(clk),
	.d(n186078));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__24_ (.o(regtop_dchdi_w1_hdi00[1112]),
	.ck(clk),
	.d(n186077));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__25_ (.o(regtop_dchdi_w1_hdi00[1113]),
	.ck(clk),
	.d(n186076));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__26_ (.o(regtop_dchdi_w1_hdi00[1114]),
	.ck(clk),
	.d(n186075));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__27_ (.o(regtop_dchdi_w1_hdi00[1115]),
	.ck(clk),
	.d(n186074));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__28_ (.o(regtop_dchdi_w1_hdi00[1116]),
	.ck(clk),
	.d(n186073));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__29_ (.o(regtop_dchdi_w1_hdi00[1117]),
	.ck(clk),
	.d(n186072));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__30_ (.o(regtop_dchdi_w1_hdi00[1118]),
	.ck(clk),
	.d(n186071));
   ms00f80 regtop_dchdi_w1_hdi00_reg_18__31_ (.o(regtop_dchdi_w1_hdi00[1119]),
	.ck(clk),
	.d(n186070));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__0_ (.o(regtop_dchdi_w1_hdi00[1120]),
	.ck(clk),
	.d(n186069));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__1_ (.o(regtop_dchdi_w1_hdi00[1121]),
	.ck(clk),
	.d(n186068));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__2_ (.o(regtop_dchdi_w1_hdi00[1122]),
	.ck(clk),
	.d(n186067));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__3_ (.o(regtop_dchdi_w1_hdi00[1123]),
	.ck(clk),
	.d(n186066));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__4_ (.o(regtop_dchdi_w1_hdi00[1124]),
	.ck(clk),
	.d(n186065));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__5_ (.o(regtop_dchdi_w1_hdi00[1125]),
	.ck(clk),
	.d(n186064));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__6_ (.o(regtop_dchdi_w1_hdi00[1126]),
	.ck(clk),
	.d(n186063));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__7_ (.o(regtop_dchdi_w1_hdi00[1127]),
	.ck(clk),
	.d(n186062));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__8_ (.o(regtop_dchdi_w1_hdi00[1128]),
	.ck(clk),
	.d(n186061));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__9_ (.o(regtop_dchdi_w1_hdi00[1129]),
	.ck(clk),
	.d(n186060));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__10_ (.o(regtop_dchdi_w1_hdi00[1130]),
	.ck(clk),
	.d(n186059));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__11_ (.o(regtop_dchdi_w1_hdi00[1131]),
	.ck(clk),
	.d(n186058));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__12_ (.o(regtop_dchdi_w1_hdi00[1132]),
	.ck(clk),
	.d(n186057));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__13_ (.o(regtop_dchdi_w1_hdi00[1133]),
	.ck(clk),
	.d(n186056));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__14_ (.o(regtop_dchdi_w1_hdi00[1134]),
	.ck(clk),
	.d(n186055));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__15_ (.o(regtop_dchdi_w1_hdi00[1135]),
	.ck(clk),
	.d(n186054));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__16_ (.o(regtop_dchdi_w1_hdi00[1136]),
	.ck(clk),
	.d(n186053));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__17_ (.o(regtop_dchdi_w1_hdi00[1137]),
	.ck(clk),
	.d(n186052));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__18_ (.o(regtop_dchdi_w1_hdi00[1138]),
	.ck(clk),
	.d(n186051));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__19_ (.o(regtop_dchdi_w1_hdi00[1139]),
	.ck(clk),
	.d(n186050));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__20_ (.o(regtop_dchdi_w1_hdi00[1140]),
	.ck(clk),
	.d(n186049));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__21_ (.o(regtop_dchdi_w1_hdi00[1141]),
	.ck(clk),
	.d(n186048));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__22_ (.o(regtop_dchdi_w1_hdi00[1142]),
	.ck(clk),
	.d(n186047));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__23_ (.o(regtop_dchdi_w1_hdi00[1143]),
	.ck(clk),
	.d(n186046));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__24_ (.o(regtop_dchdi_w1_hdi00[1144]),
	.ck(clk),
	.d(n186045));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__25_ (.o(regtop_dchdi_w1_hdi00[1145]),
	.ck(clk),
	.d(n186044));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__26_ (.o(regtop_dchdi_w1_hdi00[1146]),
	.ck(clk),
	.d(n186043));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__27_ (.o(regtop_dchdi_w1_hdi00[1147]),
	.ck(clk),
	.d(n186042));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__28_ (.o(regtop_dchdi_w1_hdi00[1148]),
	.ck(clk),
	.d(n186041));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__29_ (.o(regtop_dchdi_w1_hdi00[1149]),
	.ck(clk),
	.d(n186040));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__30_ (.o(regtop_dchdi_w1_hdi00[1150]),
	.ck(clk),
	.d(n186039));
   ms00f80 regtop_dchdi_w1_hdi00_reg_19__31_ (.o(regtop_dchdi_w1_hdi00[1151]),
	.ck(clk),
	.d(n186038));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__0_ (.o(regtop_dchdi_w1_hdi00[1152]),
	.ck(clk),
	.d(n186037));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__1_ (.o(regtop_dchdi_w1_hdi00[1153]),
	.ck(clk),
	.d(n186036));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__2_ (.o(regtop_dchdi_w1_hdi00[1154]),
	.ck(clk),
	.d(n186035));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__3_ (.o(regtop_dchdi_w1_hdi00[1155]),
	.ck(clk),
	.d(n186034));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__4_ (.o(regtop_dchdi_w1_hdi00[1156]),
	.ck(clk),
	.d(n186033));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__5_ (.o(regtop_dchdi_w1_hdi00[1157]),
	.ck(clk),
	.d(n186032));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__6_ (.o(regtop_dchdi_w1_hdi00[1158]),
	.ck(clk),
	.d(n186031));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__7_ (.o(regtop_dchdi_w1_hdi00[1159]),
	.ck(clk),
	.d(n186030));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__8_ (.o(regtop_dchdi_w1_hdi00[1160]),
	.ck(clk),
	.d(n186029));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__9_ (.o(regtop_dchdi_w1_hdi00[1161]),
	.ck(clk),
	.d(n186028));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__10_ (.o(regtop_dchdi_w1_hdi00[1162]),
	.ck(clk),
	.d(n186027));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__11_ (.o(regtop_dchdi_w1_hdi00[1163]),
	.ck(clk),
	.d(n186026));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__12_ (.o(regtop_dchdi_w1_hdi00[1164]),
	.ck(clk),
	.d(n186025));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__13_ (.o(regtop_dchdi_w1_hdi00[1165]),
	.ck(clk),
	.d(n186024));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__14_ (.o(regtop_dchdi_w1_hdi00[1166]),
	.ck(clk),
	.d(n186023));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__15_ (.o(regtop_dchdi_w1_hdi00[1167]),
	.ck(clk),
	.d(n186022));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__16_ (.o(regtop_dchdi_w1_hdi00[1168]),
	.ck(clk),
	.d(n186021));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__17_ (.o(regtop_dchdi_w1_hdi00[1169]),
	.ck(clk),
	.d(n186020));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__18_ (.o(regtop_dchdi_w1_hdi00[1170]),
	.ck(clk),
	.d(n186019));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__19_ (.o(regtop_dchdi_w1_hdi00[1171]),
	.ck(clk),
	.d(n186018));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__20_ (.o(regtop_dchdi_w1_hdi00[1172]),
	.ck(clk),
	.d(n186017));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__21_ (.o(regtop_dchdi_w1_hdi00[1173]),
	.ck(clk),
	.d(n186016));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__22_ (.o(regtop_dchdi_w1_hdi00[1174]),
	.ck(clk),
	.d(n186015));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__23_ (.o(regtop_dchdi_w1_hdi00[1175]),
	.ck(clk),
	.d(n186014));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__24_ (.o(regtop_dchdi_w1_hdi00[1176]),
	.ck(clk),
	.d(n186013));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__25_ (.o(regtop_dchdi_w1_hdi00[1177]),
	.ck(clk),
	.d(n186012));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__26_ (.o(regtop_dchdi_w1_hdi00[1178]),
	.ck(clk),
	.d(n186011));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__27_ (.o(regtop_dchdi_w1_hdi00[1179]),
	.ck(clk),
	.d(n186010));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__28_ (.o(regtop_dchdi_w1_hdi00[1180]),
	.ck(clk),
	.d(n186009));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__29_ (.o(regtop_dchdi_w1_hdi00[1181]),
	.ck(clk),
	.d(n186008));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__30_ (.o(regtop_dchdi_w1_hdi00[1182]),
	.ck(clk),
	.d(n186007));
   ms00f80 regtop_dchdi_w1_hdi00_reg_20__31_ (.o(regtop_dchdi_w1_hdi00[1183]),
	.ck(clk),
	.d(n186006));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__0_ (.o(regtop_dchdi_w1_hdi00[1184]),
	.ck(clk),
	.d(n186005));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__1_ (.o(regtop_dchdi_w1_hdi00[1185]),
	.ck(clk),
	.d(n186004));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__2_ (.o(regtop_dchdi_w1_hdi00[1186]),
	.ck(clk),
	.d(n186003));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__3_ (.o(regtop_dchdi_w1_hdi00[1187]),
	.ck(clk),
	.d(n186002));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__4_ (.o(regtop_dchdi_w1_hdi00[1188]),
	.ck(clk),
	.d(n186001));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__5_ (.o(regtop_dchdi_w1_hdi00[1189]),
	.ck(clk),
	.d(n186000));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__6_ (.o(regtop_dchdi_w1_hdi00[1190]),
	.ck(clk),
	.d(n185999));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__7_ (.o(regtop_dchdi_w1_hdi00[1191]),
	.ck(clk),
	.d(n185998));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__8_ (.o(regtop_dchdi_w1_hdi00[1192]),
	.ck(clk),
	.d(n185997));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__9_ (.o(regtop_dchdi_w1_hdi00[1193]),
	.ck(clk),
	.d(n185996));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__10_ (.o(regtop_dchdi_w1_hdi00[1194]),
	.ck(clk),
	.d(n185995));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__11_ (.o(regtop_dchdi_w1_hdi00[1195]),
	.ck(clk),
	.d(n185994));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__12_ (.o(regtop_dchdi_w1_hdi00[1196]),
	.ck(clk),
	.d(n185993));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__13_ (.o(regtop_dchdi_w1_hdi00[1197]),
	.ck(clk),
	.d(n185992));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__14_ (.o(regtop_dchdi_w1_hdi00[1198]),
	.ck(clk),
	.d(n185991));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__15_ (.o(regtop_dchdi_w1_hdi00[1199]),
	.ck(clk),
	.d(n185990));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__16_ (.o(regtop_dchdi_w1_hdi00[1200]),
	.ck(clk),
	.d(n185989));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__17_ (.o(regtop_dchdi_w1_hdi00[1201]),
	.ck(clk),
	.d(n185988));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__18_ (.o(regtop_dchdi_w1_hdi00[1202]),
	.ck(clk),
	.d(n185987));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__19_ (.o(regtop_dchdi_w1_hdi00[1203]),
	.ck(clk),
	.d(n185986));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__20_ (.o(regtop_dchdi_w1_hdi00[1204]),
	.ck(clk),
	.d(n185985));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__21_ (.o(regtop_dchdi_w1_hdi00[1205]),
	.ck(clk),
	.d(n185984));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__22_ (.o(regtop_dchdi_w1_hdi00[1206]),
	.ck(clk),
	.d(n185983));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__23_ (.o(regtop_dchdi_w1_hdi00[1207]),
	.ck(clk),
	.d(n185982));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__24_ (.o(regtop_dchdi_w1_hdi00[1208]),
	.ck(clk),
	.d(n185981));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__25_ (.o(regtop_dchdi_w1_hdi00[1209]),
	.ck(clk),
	.d(n185980));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__26_ (.o(regtop_dchdi_w1_hdi00[1210]),
	.ck(clk),
	.d(n185979));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__27_ (.o(regtop_dchdi_w1_hdi00[1211]),
	.ck(clk),
	.d(n185978));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__28_ (.o(regtop_dchdi_w1_hdi00[1212]),
	.ck(clk),
	.d(n185977));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__29_ (.o(regtop_dchdi_w1_hdi00[1213]),
	.ck(clk),
	.d(n185976));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__30_ (.o(regtop_dchdi_w1_hdi00[1214]),
	.ck(clk),
	.d(n185975));
   ms00f80 regtop_dchdi_w1_hdi00_reg_21__31_ (.o(regtop_dchdi_w1_hdi00[1215]),
	.ck(clk),
	.d(n185974));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__0_ (.o(regtop_dchdi_w1_hdi00[1216]),
	.ck(clk),
	.d(n185973));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__1_ (.o(regtop_dchdi_w1_hdi00[1217]),
	.ck(clk),
	.d(n185972));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__2_ (.o(regtop_dchdi_w1_hdi00[1218]),
	.ck(clk),
	.d(n185971));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__3_ (.o(regtop_dchdi_w1_hdi00[1219]),
	.ck(clk),
	.d(n185970));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__4_ (.o(regtop_dchdi_w1_hdi00[1220]),
	.ck(clk),
	.d(n185969));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__5_ (.o(regtop_dchdi_w1_hdi00[1221]),
	.ck(clk),
	.d(n185968));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__6_ (.o(regtop_dchdi_w1_hdi00[1222]),
	.ck(clk),
	.d(n185967));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__7_ (.o(regtop_dchdi_w1_hdi00[1223]),
	.ck(clk),
	.d(n185966));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__8_ (.o(regtop_dchdi_w1_hdi00[1224]),
	.ck(clk),
	.d(n185965));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__9_ (.o(regtop_dchdi_w1_hdi00[1225]),
	.ck(clk),
	.d(n185964));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__10_ (.o(regtop_dchdi_w1_hdi00[1226]),
	.ck(clk),
	.d(n185963));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__11_ (.o(regtop_dchdi_w1_hdi00[1227]),
	.ck(clk),
	.d(n185962));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__12_ (.o(regtop_dchdi_w1_hdi00[1228]),
	.ck(clk),
	.d(n185961));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__13_ (.o(regtop_dchdi_w1_hdi00[1229]),
	.ck(clk),
	.d(n185960));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__14_ (.o(regtop_dchdi_w1_hdi00[1230]),
	.ck(clk),
	.d(n185959));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__15_ (.o(regtop_dchdi_w1_hdi00[1231]),
	.ck(clk),
	.d(n185958));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__16_ (.o(regtop_dchdi_w1_hdi00[1232]),
	.ck(clk),
	.d(n185957));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__17_ (.o(regtop_dchdi_w1_hdi00[1233]),
	.ck(clk),
	.d(n185956));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__18_ (.o(regtop_dchdi_w1_hdi00[1234]),
	.ck(clk),
	.d(n185955));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__19_ (.o(regtop_dchdi_w1_hdi00[1235]),
	.ck(clk),
	.d(n185954));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__20_ (.o(regtop_dchdi_w1_hdi00[1236]),
	.ck(clk),
	.d(n185953));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__21_ (.o(regtop_dchdi_w1_hdi00[1237]),
	.ck(clk),
	.d(n185952));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__22_ (.o(regtop_dchdi_w1_hdi00[1238]),
	.ck(clk),
	.d(n185951));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__23_ (.o(regtop_dchdi_w1_hdi00[1239]),
	.ck(clk),
	.d(n185950));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__24_ (.o(regtop_dchdi_w1_hdi00[1240]),
	.ck(clk),
	.d(n185949));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__25_ (.o(regtop_dchdi_w1_hdi00[1241]),
	.ck(clk),
	.d(n185948));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__26_ (.o(regtop_dchdi_w1_hdi00[1242]),
	.ck(clk),
	.d(n185947));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__27_ (.o(regtop_dchdi_w1_hdi00[1243]),
	.ck(clk),
	.d(n185946));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__28_ (.o(regtop_dchdi_w1_hdi00[1244]),
	.ck(clk),
	.d(n185945));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__29_ (.o(regtop_dchdi_w1_hdi00[1245]),
	.ck(clk),
	.d(n185944));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__30_ (.o(regtop_dchdi_w1_hdi00[1246]),
	.ck(clk),
	.d(n185943));
   ms00f80 regtop_dchdi_w1_hdi00_reg_22__31_ (.o(regtop_dchdi_w1_hdi00[1247]),
	.ck(clk),
	.d(n185942));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__0_ (.o(regtop_dchdi_w1_hdi00[1248]),
	.ck(clk),
	.d(n185941));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__1_ (.o(regtop_dchdi_w1_hdi00[1249]),
	.ck(clk),
	.d(n185940));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__2_ (.o(regtop_dchdi_w1_hdi00[1250]),
	.ck(clk),
	.d(n185939));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__3_ (.o(regtop_dchdi_w1_hdi00[1251]),
	.ck(clk),
	.d(n185938));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__4_ (.o(regtop_dchdi_w1_hdi00[1252]),
	.ck(clk),
	.d(n185937));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__5_ (.o(regtop_dchdi_w1_hdi00[1253]),
	.ck(clk),
	.d(n185936));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__6_ (.o(regtop_dchdi_w1_hdi00[1254]),
	.ck(clk),
	.d(n185935));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__7_ (.o(regtop_dchdi_w1_hdi00[1255]),
	.ck(clk),
	.d(n185934));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__8_ (.o(regtop_dchdi_w1_hdi00[1256]),
	.ck(clk),
	.d(n185933));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__9_ (.o(regtop_dchdi_w1_hdi00[1257]),
	.ck(clk),
	.d(n185932));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__10_ (.o(regtop_dchdi_w1_hdi00[1258]),
	.ck(clk),
	.d(n185931));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__11_ (.o(regtop_dchdi_w1_hdi00[1259]),
	.ck(clk),
	.d(n185930));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__12_ (.o(regtop_dchdi_w1_hdi00[1260]),
	.ck(clk),
	.d(n185929));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__13_ (.o(regtop_dchdi_w1_hdi00[1261]),
	.ck(clk),
	.d(n185928));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__14_ (.o(regtop_dchdi_w1_hdi00[1262]),
	.ck(clk),
	.d(n185927));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__15_ (.o(regtop_dchdi_w1_hdi00[1263]),
	.ck(clk),
	.d(n185926));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__16_ (.o(regtop_dchdi_w1_hdi00[1264]),
	.ck(clk),
	.d(n185925));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__17_ (.o(regtop_dchdi_w1_hdi00[1265]),
	.ck(clk),
	.d(n185924));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__18_ (.o(regtop_dchdi_w1_hdi00[1266]),
	.ck(clk),
	.d(n185923));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__19_ (.o(regtop_dchdi_w1_hdi00[1267]),
	.ck(clk),
	.d(n185922));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__20_ (.o(regtop_dchdi_w1_hdi00[1268]),
	.ck(clk),
	.d(n185921));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__21_ (.o(regtop_dchdi_w1_hdi00[1269]),
	.ck(clk),
	.d(n185920));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__22_ (.o(regtop_dchdi_w1_hdi00[1270]),
	.ck(clk),
	.d(n185919));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__23_ (.o(regtop_dchdi_w1_hdi00[1271]),
	.ck(clk),
	.d(n185918));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__24_ (.o(regtop_dchdi_w1_hdi00[1272]),
	.ck(clk),
	.d(n185917));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__25_ (.o(regtop_dchdi_w1_hdi00[1273]),
	.ck(clk),
	.d(n185916));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__26_ (.o(regtop_dchdi_w1_hdi00[1274]),
	.ck(clk),
	.d(n185915));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__27_ (.o(regtop_dchdi_w1_hdi00[1275]),
	.ck(clk),
	.d(n185914));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__28_ (.o(regtop_dchdi_w1_hdi00[1276]),
	.ck(clk),
	.d(n185913));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__29_ (.o(regtop_dchdi_w1_hdi00[1277]),
	.ck(clk),
	.d(n185912));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__30_ (.o(regtop_dchdi_w1_hdi00[1278]),
	.ck(clk),
	.d(n185911));
   ms00f80 regtop_dchdi_w1_hdi00_reg_23__31_ (.o(regtop_dchdi_w1_hdi00[1279]),
	.ck(clk),
	.d(n185910));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__0_ (.o(regtop_dchdi_w1_hdi00[1280]),
	.ck(clk),
	.d(n185909));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__1_ (.o(regtop_dchdi_w1_hdi00[1281]),
	.ck(clk),
	.d(n185908));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__2_ (.o(regtop_dchdi_w1_hdi00[1282]),
	.ck(clk),
	.d(n185907));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__3_ (.o(regtop_dchdi_w1_hdi00[1283]),
	.ck(clk),
	.d(n185906));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__4_ (.o(regtop_dchdi_w1_hdi00[1284]),
	.ck(clk),
	.d(n185905));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__5_ (.o(regtop_dchdi_w1_hdi00[1285]),
	.ck(clk),
	.d(n185904));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__6_ (.o(regtop_dchdi_w1_hdi00[1286]),
	.ck(clk),
	.d(n185903));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__7_ (.o(regtop_dchdi_w1_hdi00[1287]),
	.ck(clk),
	.d(n185902));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__8_ (.o(regtop_dchdi_w1_hdi00[1288]),
	.ck(clk),
	.d(n185901));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__9_ (.o(regtop_dchdi_w1_hdi00[1289]),
	.ck(clk),
	.d(n185900));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__10_ (.o(regtop_dchdi_w1_hdi00[1290]),
	.ck(clk),
	.d(n185899));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__11_ (.o(regtop_dchdi_w1_hdi00[1291]),
	.ck(clk),
	.d(n185898));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__12_ (.o(regtop_dchdi_w1_hdi00[1292]),
	.ck(clk),
	.d(n185897));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__13_ (.o(regtop_dchdi_w1_hdi00[1293]),
	.ck(clk),
	.d(n185896));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__14_ (.o(regtop_dchdi_w1_hdi00[1294]),
	.ck(clk),
	.d(n185895));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__15_ (.o(regtop_dchdi_w1_hdi00[1295]),
	.ck(clk),
	.d(n185894));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__16_ (.o(regtop_dchdi_w1_hdi00[1296]),
	.ck(clk),
	.d(n185893));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__17_ (.o(regtop_dchdi_w1_hdi00[1297]),
	.ck(clk),
	.d(n185892));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__18_ (.o(regtop_dchdi_w1_hdi00[1298]),
	.ck(clk),
	.d(n185891));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__19_ (.o(regtop_dchdi_w1_hdi00[1299]),
	.ck(clk),
	.d(n185890));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__20_ (.o(regtop_dchdi_w1_hdi00[1300]),
	.ck(clk),
	.d(n185889));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__21_ (.o(regtop_dchdi_w1_hdi00[1301]),
	.ck(clk),
	.d(n185888));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__22_ (.o(regtop_dchdi_w1_hdi00[1302]),
	.ck(clk),
	.d(n185887));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__23_ (.o(regtop_dchdi_w1_hdi00[1303]),
	.ck(clk),
	.d(n185886));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__24_ (.o(regtop_dchdi_w1_hdi00[1304]),
	.ck(clk),
	.d(n185885));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__25_ (.o(regtop_dchdi_w1_hdi00[1305]),
	.ck(clk),
	.d(n185884));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__26_ (.o(regtop_dchdi_w1_hdi00[1306]),
	.ck(clk),
	.d(n185883));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__27_ (.o(regtop_dchdi_w1_hdi00[1307]),
	.ck(clk),
	.d(n185882));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__28_ (.o(regtop_dchdi_w1_hdi00[1308]),
	.ck(clk),
	.d(n185881));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__29_ (.o(regtop_dchdi_w1_hdi00[1309]),
	.ck(clk),
	.d(n185880));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__30_ (.o(regtop_dchdi_w1_hdi00[1310]),
	.ck(clk),
	.d(n185879));
   ms00f80 regtop_dchdi_w1_hdi00_reg_24__31_ (.o(regtop_dchdi_w1_hdi00[1311]),
	.ck(clk),
	.d(n185878));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__0_ (.o(regtop_dchdi_w1_hdi00[1312]),
	.ck(clk),
	.d(n185877));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__1_ (.o(regtop_dchdi_w1_hdi00[1313]),
	.ck(clk),
	.d(n185876));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__2_ (.o(regtop_dchdi_w1_hdi00[1314]),
	.ck(clk),
	.d(n185875));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__3_ (.o(regtop_dchdi_w1_hdi00[1315]),
	.ck(clk),
	.d(n185874));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__4_ (.o(regtop_dchdi_w1_hdi00[1316]),
	.ck(clk),
	.d(n185873));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__5_ (.o(regtop_dchdi_w1_hdi00[1317]),
	.ck(clk),
	.d(n185872));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__6_ (.o(regtop_dchdi_w1_hdi00[1318]),
	.ck(clk),
	.d(n185871));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__7_ (.o(regtop_dchdi_w1_hdi00[1319]),
	.ck(clk),
	.d(n185870));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__8_ (.o(regtop_dchdi_w1_hdi00[1320]),
	.ck(clk),
	.d(n185869));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__9_ (.o(regtop_dchdi_w1_hdi00[1321]),
	.ck(clk),
	.d(n185868));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__10_ (.o(regtop_dchdi_w1_hdi00[1322]),
	.ck(clk),
	.d(n185867));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__11_ (.o(regtop_dchdi_w1_hdi00[1323]),
	.ck(clk),
	.d(n185866));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__12_ (.o(regtop_dchdi_w1_hdi00[1324]),
	.ck(clk),
	.d(n185865));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__13_ (.o(regtop_dchdi_w1_hdi00[1325]),
	.ck(clk),
	.d(n185864));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__14_ (.o(regtop_dchdi_w1_hdi00[1326]),
	.ck(clk),
	.d(n185863));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__15_ (.o(regtop_dchdi_w1_hdi00[1327]),
	.ck(clk),
	.d(n185862));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__16_ (.o(regtop_dchdi_w1_hdi00[1328]),
	.ck(clk),
	.d(n185861));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__17_ (.o(regtop_dchdi_w1_hdi00[1329]),
	.ck(clk),
	.d(n185860));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__18_ (.o(regtop_dchdi_w1_hdi00[1330]),
	.ck(clk),
	.d(n185859));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__19_ (.o(regtop_dchdi_w1_hdi00[1331]),
	.ck(clk),
	.d(n185858));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__20_ (.o(regtop_dchdi_w1_hdi00[1332]),
	.ck(clk),
	.d(n185857));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__21_ (.o(regtop_dchdi_w1_hdi00[1333]),
	.ck(clk),
	.d(n185856));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__22_ (.o(regtop_dchdi_w1_hdi00[1334]),
	.ck(clk),
	.d(n185855));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__23_ (.o(regtop_dchdi_w1_hdi00[1335]),
	.ck(clk),
	.d(n185854));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__24_ (.o(regtop_dchdi_w1_hdi00[1336]),
	.ck(clk),
	.d(n185853));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__25_ (.o(regtop_dchdi_w1_hdi00[1337]),
	.ck(clk),
	.d(n185852));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__26_ (.o(regtop_dchdi_w1_hdi00[1338]),
	.ck(clk),
	.d(n185851));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__27_ (.o(regtop_dchdi_w1_hdi00[1339]),
	.ck(clk),
	.d(n185850));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__28_ (.o(regtop_dchdi_w1_hdi00[1340]),
	.ck(clk),
	.d(n185849));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__29_ (.o(regtop_dchdi_w1_hdi00[1341]),
	.ck(clk),
	.d(n185848));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__30_ (.o(regtop_dchdi_w1_hdi00[1342]),
	.ck(clk),
	.d(n185847));
   ms00f80 regtop_dchdi_w1_hdi00_reg_25__31_ (.o(regtop_dchdi_w1_hdi00[1343]),
	.ck(clk),
	.d(n185846));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__0_ (.o(regtop_dchdi_w1_hdi00[1344]),
	.ck(clk),
	.d(n185845));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__1_ (.o(regtop_dchdi_w1_hdi00[1345]),
	.ck(clk),
	.d(n185844));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__2_ (.o(regtop_dchdi_w1_hdi00[1346]),
	.ck(clk),
	.d(n185843));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__3_ (.o(regtop_dchdi_w1_hdi00[1347]),
	.ck(clk),
	.d(n185842));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__4_ (.o(regtop_dchdi_w1_hdi00[1348]),
	.ck(clk),
	.d(n185841));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__5_ (.o(regtop_dchdi_w1_hdi00[1349]),
	.ck(clk),
	.d(n185840));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__6_ (.o(regtop_dchdi_w1_hdi00[1350]),
	.ck(clk),
	.d(n185839));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__7_ (.o(regtop_dchdi_w1_hdi00[1351]),
	.ck(clk),
	.d(n185838));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__8_ (.o(regtop_dchdi_w1_hdi00[1352]),
	.ck(clk),
	.d(n185837));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__9_ (.o(regtop_dchdi_w1_hdi00[1353]),
	.ck(clk),
	.d(n185836));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__10_ (.o(regtop_dchdi_w1_hdi00[1354]),
	.ck(clk),
	.d(n185835));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__11_ (.o(regtop_dchdi_w1_hdi00[1355]),
	.ck(clk),
	.d(n185834));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__12_ (.o(regtop_dchdi_w1_hdi00[1356]),
	.ck(clk),
	.d(n185833));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__13_ (.o(regtop_dchdi_w1_hdi00[1357]),
	.ck(clk),
	.d(n185832));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__14_ (.o(regtop_dchdi_w1_hdi00[1358]),
	.ck(clk),
	.d(n185831));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__15_ (.o(regtop_dchdi_w1_hdi00[1359]),
	.ck(clk),
	.d(n185830));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__16_ (.o(regtop_dchdi_w1_hdi00[1360]),
	.ck(clk),
	.d(n185829));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__17_ (.o(regtop_dchdi_w1_hdi00[1361]),
	.ck(clk),
	.d(n185828));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__18_ (.o(regtop_dchdi_w1_hdi00[1362]),
	.ck(clk),
	.d(n185827));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__19_ (.o(regtop_dchdi_w1_hdi00[1363]),
	.ck(clk),
	.d(n185826));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__20_ (.o(regtop_dchdi_w1_hdi00[1364]),
	.ck(clk),
	.d(n185825));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__21_ (.o(regtop_dchdi_w1_hdi00[1365]),
	.ck(clk),
	.d(n185824));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__22_ (.o(regtop_dchdi_w1_hdi00[1366]),
	.ck(clk),
	.d(n185823));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__23_ (.o(regtop_dchdi_w1_hdi00[1367]),
	.ck(clk),
	.d(n185822));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__24_ (.o(regtop_dchdi_w1_hdi00[1368]),
	.ck(clk),
	.d(n185821));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__25_ (.o(regtop_dchdi_w1_hdi00[1369]),
	.ck(clk),
	.d(n185820));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__26_ (.o(regtop_dchdi_w1_hdi00[1370]),
	.ck(clk),
	.d(n185819));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__27_ (.o(regtop_dchdi_w1_hdi00[1371]),
	.ck(clk),
	.d(n185818));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__28_ (.o(regtop_dchdi_w1_hdi00[1372]),
	.ck(clk),
	.d(n185817));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__29_ (.o(regtop_dchdi_w1_hdi00[1373]),
	.ck(clk),
	.d(n185816));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__30_ (.o(regtop_dchdi_w1_hdi00[1374]),
	.ck(clk),
	.d(n185815));
   ms00f80 regtop_dchdi_w1_hdi00_reg_26__31_ (.o(regtop_dchdi_w1_hdi00[1375]),
	.ck(clk),
	.d(n185814));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__0_ (.o(regtop_dchdi_w1_hdi00[1376]),
	.ck(clk),
	.d(n185813));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__1_ (.o(regtop_dchdi_w1_hdi00[1377]),
	.ck(clk),
	.d(n185812));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__2_ (.o(regtop_dchdi_w1_hdi00[1378]),
	.ck(clk),
	.d(n185811));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__3_ (.o(regtop_dchdi_w1_hdi00[1379]),
	.ck(clk),
	.d(n185810));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__4_ (.o(regtop_dchdi_w1_hdi00[1380]),
	.ck(clk),
	.d(n185809));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__5_ (.o(regtop_dchdi_w1_hdi00[1381]),
	.ck(clk),
	.d(n185808));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__6_ (.o(regtop_dchdi_w1_hdi00[1382]),
	.ck(clk),
	.d(n185807));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__7_ (.o(regtop_dchdi_w1_hdi00[1383]),
	.ck(clk),
	.d(n185806));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__8_ (.o(regtop_dchdi_w1_hdi00[1384]),
	.ck(clk),
	.d(n185805));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__9_ (.o(regtop_dchdi_w1_hdi00[1385]),
	.ck(clk),
	.d(n185804));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__10_ (.o(regtop_dchdi_w1_hdi00[1386]),
	.ck(clk),
	.d(n185803));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__11_ (.o(regtop_dchdi_w1_hdi00[1387]),
	.ck(clk),
	.d(n185802));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__12_ (.o(regtop_dchdi_w1_hdi00[1388]),
	.ck(clk),
	.d(n185801));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__13_ (.o(regtop_dchdi_w1_hdi00[1389]),
	.ck(clk),
	.d(n185800));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__14_ (.o(regtop_dchdi_w1_hdi00[1390]),
	.ck(clk),
	.d(n185799));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__15_ (.o(regtop_dchdi_w1_hdi00[1391]),
	.ck(clk),
	.d(n185798));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__16_ (.o(regtop_dchdi_w1_hdi00[1392]),
	.ck(clk),
	.d(n185797));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__17_ (.o(regtop_dchdi_w1_hdi00[1393]),
	.ck(clk),
	.d(n185796));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__18_ (.o(regtop_dchdi_w1_hdi00[1394]),
	.ck(clk),
	.d(n185795));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__19_ (.o(regtop_dchdi_w1_hdi00[1395]),
	.ck(clk),
	.d(n185794));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__20_ (.o(regtop_dchdi_w1_hdi00[1396]),
	.ck(clk),
	.d(n185793));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__21_ (.o(regtop_dchdi_w1_hdi00[1397]),
	.ck(clk),
	.d(n185792));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__22_ (.o(regtop_dchdi_w1_hdi00[1398]),
	.ck(clk),
	.d(n185791));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__23_ (.o(regtop_dchdi_w1_hdi00[1399]),
	.ck(clk),
	.d(n185790));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__24_ (.o(regtop_dchdi_w1_hdi00[1400]),
	.ck(clk),
	.d(n185789));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__25_ (.o(regtop_dchdi_w1_hdi00[1401]),
	.ck(clk),
	.d(n185788));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__26_ (.o(regtop_dchdi_w1_hdi00[1402]),
	.ck(clk),
	.d(n185787));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__27_ (.o(regtop_dchdi_w1_hdi00[1403]),
	.ck(clk),
	.d(n185786));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__28_ (.o(regtop_dchdi_w1_hdi00[1404]),
	.ck(clk),
	.d(n185785));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__29_ (.o(regtop_dchdi_w1_hdi00[1405]),
	.ck(clk),
	.d(n185784));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__30_ (.o(regtop_dchdi_w1_hdi00[1406]),
	.ck(clk),
	.d(n185783));
   ms00f80 regtop_dchdi_w1_hdi00_reg_27__31_ (.o(regtop_dchdi_w1_hdi00[1407]),
	.ck(clk),
	.d(n185782));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__0_ (.o(regtop_dchdi_w1_hdi00[1408]),
	.ck(clk),
	.d(n185781));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__1_ (.o(regtop_dchdi_w1_hdi00[1409]),
	.ck(clk),
	.d(n185780));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__2_ (.o(regtop_dchdi_w1_hdi00[1410]),
	.ck(clk),
	.d(n185779));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__3_ (.o(regtop_dchdi_w1_hdi00[1411]),
	.ck(clk),
	.d(n185778));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__4_ (.o(regtop_dchdi_w1_hdi00[1412]),
	.ck(clk),
	.d(n185777));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__5_ (.o(regtop_dchdi_w1_hdi00[1413]),
	.ck(clk),
	.d(n185776));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__6_ (.o(regtop_dchdi_w1_hdi00[1414]),
	.ck(clk),
	.d(n185775));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__7_ (.o(regtop_dchdi_w1_hdi00[1415]),
	.ck(clk),
	.d(n185774));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__8_ (.o(regtop_dchdi_w1_hdi00[1416]),
	.ck(clk),
	.d(n185773));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__9_ (.o(regtop_dchdi_w1_hdi00[1417]),
	.ck(clk),
	.d(n185772));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__10_ (.o(regtop_dchdi_w1_hdi00[1418]),
	.ck(clk),
	.d(n185771));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__11_ (.o(regtop_dchdi_w1_hdi00[1419]),
	.ck(clk),
	.d(n185770));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__12_ (.o(regtop_dchdi_w1_hdi00[1420]),
	.ck(clk),
	.d(n185769));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__13_ (.o(regtop_dchdi_w1_hdi00[1421]),
	.ck(clk),
	.d(n185768));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__14_ (.o(regtop_dchdi_w1_hdi00[1422]),
	.ck(clk),
	.d(n185767));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__15_ (.o(regtop_dchdi_w1_hdi00[1423]),
	.ck(clk),
	.d(n185766));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__16_ (.o(regtop_dchdi_w1_hdi00[1424]),
	.ck(clk),
	.d(n185765));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__17_ (.o(regtop_dchdi_w1_hdi00[1425]),
	.ck(clk),
	.d(n185764));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__18_ (.o(regtop_dchdi_w1_hdi00[1426]),
	.ck(clk),
	.d(n185763));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__19_ (.o(regtop_dchdi_w1_hdi00[1427]),
	.ck(clk),
	.d(n185762));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__20_ (.o(regtop_dchdi_w1_hdi00[1428]),
	.ck(clk),
	.d(n185761));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__21_ (.o(regtop_dchdi_w1_hdi00[1429]),
	.ck(clk),
	.d(n185760));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__22_ (.o(regtop_dchdi_w1_hdi00[1430]),
	.ck(clk),
	.d(n185759));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__23_ (.o(regtop_dchdi_w1_hdi00[1431]),
	.ck(clk),
	.d(n185758));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__24_ (.o(regtop_dchdi_w1_hdi00[1432]),
	.ck(clk),
	.d(n185757));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__25_ (.o(regtop_dchdi_w1_hdi00[1433]),
	.ck(clk),
	.d(n185756));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__26_ (.o(regtop_dchdi_w1_hdi00[1434]),
	.ck(clk),
	.d(n185755));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__27_ (.o(regtop_dchdi_w1_hdi00[1435]),
	.ck(clk),
	.d(n185754));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__28_ (.o(regtop_dchdi_w1_hdi00[1436]),
	.ck(clk),
	.d(n185753));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__29_ (.o(regtop_dchdi_w1_hdi00[1437]),
	.ck(clk),
	.d(n185752));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__30_ (.o(regtop_dchdi_w1_hdi00[1438]),
	.ck(clk),
	.d(n185751));
   ms00f80 regtop_dchdi_w1_hdi00_reg_28__31_ (.o(regtop_dchdi_w1_hdi00[1439]),
	.ck(clk),
	.d(n185750));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__0_ (.o(regtop_dchdi_w1_hdi00[1440]),
	.ck(clk),
	.d(n185749));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__1_ (.o(regtop_dchdi_w1_hdi00[1441]),
	.ck(clk),
	.d(n185748));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__2_ (.o(regtop_dchdi_w1_hdi00[1442]),
	.ck(clk),
	.d(n185747));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__3_ (.o(regtop_dchdi_w1_hdi00[1443]),
	.ck(clk),
	.d(n185746));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__4_ (.o(regtop_dchdi_w1_hdi00[1444]),
	.ck(clk),
	.d(n185745));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__5_ (.o(regtop_dchdi_w1_hdi00[1445]),
	.ck(clk),
	.d(n185744));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__6_ (.o(regtop_dchdi_w1_hdi00[1446]),
	.ck(clk),
	.d(n185743));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__7_ (.o(regtop_dchdi_w1_hdi00[1447]),
	.ck(clk),
	.d(n185742));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__8_ (.o(regtop_dchdi_w1_hdi00[1448]),
	.ck(clk),
	.d(n185741));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__9_ (.o(regtop_dchdi_w1_hdi00[1449]),
	.ck(clk),
	.d(n185740));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__10_ (.o(regtop_dchdi_w1_hdi00[1450]),
	.ck(clk),
	.d(n185739));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__11_ (.o(regtop_dchdi_w1_hdi00[1451]),
	.ck(clk),
	.d(n185738));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__12_ (.o(regtop_dchdi_w1_hdi00[1452]),
	.ck(clk),
	.d(n185737));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__13_ (.o(regtop_dchdi_w1_hdi00[1453]),
	.ck(clk),
	.d(n185736));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__14_ (.o(regtop_dchdi_w1_hdi00[1454]),
	.ck(clk),
	.d(n185735));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__15_ (.o(regtop_dchdi_w1_hdi00[1455]),
	.ck(clk),
	.d(n185734));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__16_ (.o(regtop_dchdi_w1_hdi00[1456]),
	.ck(clk),
	.d(n185733));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__17_ (.o(regtop_dchdi_w1_hdi00[1457]),
	.ck(clk),
	.d(n185732));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__18_ (.o(regtop_dchdi_w1_hdi00[1458]),
	.ck(clk),
	.d(n185731));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__19_ (.o(regtop_dchdi_w1_hdi00[1459]),
	.ck(clk),
	.d(n185730));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__20_ (.o(regtop_dchdi_w1_hdi00[1460]),
	.ck(clk),
	.d(n185729));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__21_ (.o(regtop_dchdi_w1_hdi00[1461]),
	.ck(clk),
	.d(n185728));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__22_ (.o(regtop_dchdi_w1_hdi00[1462]),
	.ck(clk),
	.d(n185727));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__23_ (.o(regtop_dchdi_w1_hdi00[1463]),
	.ck(clk),
	.d(n185726));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__24_ (.o(regtop_dchdi_w1_hdi00[1464]),
	.ck(clk),
	.d(n185725));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__25_ (.o(regtop_dchdi_w1_hdi00[1465]),
	.ck(clk),
	.d(n185724));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__26_ (.o(regtop_dchdi_w1_hdi00[1466]),
	.ck(clk),
	.d(n185723));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__27_ (.o(regtop_dchdi_w1_hdi00[1467]),
	.ck(clk),
	.d(n185722));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__28_ (.o(regtop_dchdi_w1_hdi00[1468]),
	.ck(clk),
	.d(n185721));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__29_ (.o(regtop_dchdi_w1_hdi00[1469]),
	.ck(clk),
	.d(n185720));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__30_ (.o(regtop_dchdi_w1_hdi00[1470]),
	.ck(clk),
	.d(n185719));
   ms00f80 regtop_dchdi_w1_hdi00_reg_29__31_ (.o(regtop_dchdi_w1_hdi00[1471]),
	.ck(clk),
	.d(n185718));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__0_ (.o(regtop_dchdi_w1_hdi00[1472]),
	.ck(clk),
	.d(n185717));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__1_ (.o(regtop_dchdi_w1_hdi00[1473]),
	.ck(clk),
	.d(n185716));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__2_ (.o(regtop_dchdi_w1_hdi00[1474]),
	.ck(clk),
	.d(n185715));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__3_ (.o(regtop_dchdi_w1_hdi00[1475]),
	.ck(clk),
	.d(n185714));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__4_ (.o(regtop_dchdi_w1_hdi00[1476]),
	.ck(clk),
	.d(n185713));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__5_ (.o(regtop_dchdi_w1_hdi00[1477]),
	.ck(clk),
	.d(n185712));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__6_ (.o(regtop_dchdi_w1_hdi00[1478]),
	.ck(clk),
	.d(n185711));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__7_ (.o(regtop_dchdi_w1_hdi00[1479]),
	.ck(clk),
	.d(n185710));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__8_ (.o(regtop_dchdi_w1_hdi00[1480]),
	.ck(clk),
	.d(n185709));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__9_ (.o(regtop_dchdi_w1_hdi00[1481]),
	.ck(clk),
	.d(n185708));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__10_ (.o(regtop_dchdi_w1_hdi00[1482]),
	.ck(clk),
	.d(n185707));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__11_ (.o(regtop_dchdi_w1_hdi00[1483]),
	.ck(clk),
	.d(n185706));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__12_ (.o(regtop_dchdi_w1_hdi00[1484]),
	.ck(clk),
	.d(n185705));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__13_ (.o(regtop_dchdi_w1_hdi00[1485]),
	.ck(clk),
	.d(n185704));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__14_ (.o(regtop_dchdi_w1_hdi00[1486]),
	.ck(clk),
	.d(n185703));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__15_ (.o(regtop_dchdi_w1_hdi00[1487]),
	.ck(clk),
	.d(n185702));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__16_ (.o(regtop_dchdi_w1_hdi00[1488]),
	.ck(clk),
	.d(n185701));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__17_ (.o(regtop_dchdi_w1_hdi00[1489]),
	.ck(clk),
	.d(n185700));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__18_ (.o(regtop_dchdi_w1_hdi00[1490]),
	.ck(clk),
	.d(n185699));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__19_ (.o(regtop_dchdi_w1_hdi00[1491]),
	.ck(clk),
	.d(n185698));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__20_ (.o(regtop_dchdi_w1_hdi00[1492]),
	.ck(clk),
	.d(n185697));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__21_ (.o(regtop_dchdi_w1_hdi00[1493]),
	.ck(clk),
	.d(n185696));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__22_ (.o(regtop_dchdi_w1_hdi00[1494]),
	.ck(clk),
	.d(n185695));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__23_ (.o(regtop_dchdi_w1_hdi00[1495]),
	.ck(clk),
	.d(n185694));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__24_ (.o(regtop_dchdi_w1_hdi00[1496]),
	.ck(clk),
	.d(n185693));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__25_ (.o(regtop_dchdi_w1_hdi00[1497]),
	.ck(clk),
	.d(n185692));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__26_ (.o(regtop_dchdi_w1_hdi00[1498]),
	.ck(clk),
	.d(n185691));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__27_ (.o(regtop_dchdi_w1_hdi00[1499]),
	.ck(clk),
	.d(n185690));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__28_ (.o(regtop_dchdi_w1_hdi00[1500]),
	.ck(clk),
	.d(n185689));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__29_ (.o(regtop_dchdi_w1_hdi00[1501]),
	.ck(clk),
	.d(n185688));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__30_ (.o(regtop_dchdi_w1_hdi00[1502]),
	.ck(clk),
	.d(n185687));
   ms00f80 regtop_dchdi_w1_hdi00_reg_30__31_ (.o(regtop_dchdi_w1_hdi00[1503]),
	.ck(clk),
	.d(n185686));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__0_ (.o(regtop_dchdi_w1_hdi00[1504]),
	.ck(clk),
	.d(n185685));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__1_ (.o(regtop_dchdi_w1_hdi00[1505]),
	.ck(clk),
	.d(n185684));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__2_ (.o(regtop_dchdi_w1_hdi00[1506]),
	.ck(clk),
	.d(n185683));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__3_ (.o(regtop_dchdi_w1_hdi00[1507]),
	.ck(clk),
	.d(n185682));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__4_ (.o(regtop_dchdi_w1_hdi00[1508]),
	.ck(clk),
	.d(n185681));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__5_ (.o(regtop_dchdi_w1_hdi00[1509]),
	.ck(clk),
	.d(n185680));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__6_ (.o(regtop_dchdi_w1_hdi00[1510]),
	.ck(clk),
	.d(n185679));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__7_ (.o(regtop_dchdi_w1_hdi00[1511]),
	.ck(clk),
	.d(n185678));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__8_ (.o(regtop_dchdi_w1_hdi00[1512]),
	.ck(clk),
	.d(n185677));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__9_ (.o(regtop_dchdi_w1_hdi00[1513]),
	.ck(clk),
	.d(n185676));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__10_ (.o(regtop_dchdi_w1_hdi00[1514]),
	.ck(clk),
	.d(n185675));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__11_ (.o(regtop_dchdi_w1_hdi00[1515]),
	.ck(clk),
	.d(n185674));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__12_ (.o(regtop_dchdi_w1_hdi00[1516]),
	.ck(clk),
	.d(n185673));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__13_ (.o(regtop_dchdi_w1_hdi00[1517]),
	.ck(clk),
	.d(n185672));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__14_ (.o(regtop_dchdi_w1_hdi00[1518]),
	.ck(clk),
	.d(n185671));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__15_ (.o(regtop_dchdi_w1_hdi00[1519]),
	.ck(clk),
	.d(n185670));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__16_ (.o(regtop_dchdi_w1_hdi00[1520]),
	.ck(clk),
	.d(n185669));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__17_ (.o(regtop_dchdi_w1_hdi00[1521]),
	.ck(clk),
	.d(n185668));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__18_ (.o(regtop_dchdi_w1_hdi00[1522]),
	.ck(clk),
	.d(n185667));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__19_ (.o(regtop_dchdi_w1_hdi00[1523]),
	.ck(clk),
	.d(n185666));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__20_ (.o(regtop_dchdi_w1_hdi00[1524]),
	.ck(clk),
	.d(n185665));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__21_ (.o(regtop_dchdi_w1_hdi00[1525]),
	.ck(clk),
	.d(n185664));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__22_ (.o(regtop_dchdi_w1_hdi00[1526]),
	.ck(clk),
	.d(n185663));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__23_ (.o(regtop_dchdi_w1_hdi00[1527]),
	.ck(clk),
	.d(n185662));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__24_ (.o(regtop_dchdi_w1_hdi00[1528]),
	.ck(clk),
	.d(n185661));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__25_ (.o(regtop_dchdi_w1_hdi00[1529]),
	.ck(clk),
	.d(n185660));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__26_ (.o(regtop_dchdi_w1_hdi00[1530]),
	.ck(clk),
	.d(n185659));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__27_ (.o(regtop_dchdi_w1_hdi00[1531]),
	.ck(clk),
	.d(n185658));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__28_ (.o(regtop_dchdi_w1_hdi00[1532]),
	.ck(clk),
	.d(n185657));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__29_ (.o(regtop_dchdi_w1_hdi00[1533]),
	.ck(clk),
	.d(n185656));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__30_ (.o(regtop_dchdi_w1_hdi00[1534]),
	.ck(clk),
	.d(n185655));
   ms00f80 regtop_dchdi_w1_hdi00_reg_31__31_ (.o(regtop_dchdi_w1_hdi00[1535]),
	.ck(clk),
	.d(n185654));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__0_ (.o(regtop_dchdi_w1_hdi00[512]),
	.ck(clk),
	.d(n185653));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__1_ (.o(regtop_dchdi_w1_hdi00[513]),
	.ck(clk),
	.d(n185652));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__2_ (.o(regtop_dchdi_w1_hdi00[514]),
	.ck(clk),
	.d(n185651));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__3_ (.o(regtop_dchdi_w1_hdi00[515]),
	.ck(clk),
	.d(n185650));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__4_ (.o(regtop_dchdi_w1_hdi00[516]),
	.ck(clk),
	.d(n185649));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__5_ (.o(regtop_dchdi_w1_hdi00[517]),
	.ck(clk),
	.d(n185648));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__6_ (.o(regtop_dchdi_w1_hdi00[518]),
	.ck(clk),
	.d(n185647));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__7_ (.o(regtop_dchdi_w1_hdi00[519]),
	.ck(clk),
	.d(n185646));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__8_ (.o(regtop_dchdi_w1_hdi00[520]),
	.ck(clk),
	.d(n185645));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__9_ (.o(regtop_dchdi_w1_hdi00[521]),
	.ck(clk),
	.d(n185644));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__10_ (.o(regtop_dchdi_w1_hdi00[522]),
	.ck(clk),
	.d(n185643));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__11_ (.o(regtop_dchdi_w1_hdi00[523]),
	.ck(clk),
	.d(n185642));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__12_ (.o(regtop_dchdi_w1_hdi00[524]),
	.ck(clk),
	.d(n185641));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__13_ (.o(regtop_dchdi_w1_hdi00[525]),
	.ck(clk),
	.d(n185640));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__14_ (.o(regtop_dchdi_w1_hdi00[526]),
	.ck(clk),
	.d(n185639));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__15_ (.o(regtop_dchdi_w1_hdi00[527]),
	.ck(clk),
	.d(n185638));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__16_ (.o(regtop_dchdi_w1_hdi00[528]),
	.ck(clk),
	.d(n185637));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__17_ (.o(regtop_dchdi_w1_hdi00[529]),
	.ck(clk),
	.d(n185636));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__18_ (.o(regtop_dchdi_w1_hdi00[530]),
	.ck(clk),
	.d(n185635));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__19_ (.o(regtop_dchdi_w1_hdi00[531]),
	.ck(clk),
	.d(n185634));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__20_ (.o(regtop_dchdi_w1_hdi00[532]),
	.ck(clk),
	.d(n185633));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__21_ (.o(regtop_dchdi_w1_hdi00[533]),
	.ck(clk),
	.d(n185632));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__22_ (.o(regtop_dchdi_w1_hdi00[534]),
	.ck(clk),
	.d(n185631));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__23_ (.o(regtop_dchdi_w1_hdi00[535]),
	.ck(clk),
	.d(n185630));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__24_ (.o(regtop_dchdi_w1_hdi00[536]),
	.ck(clk),
	.d(n185629));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__25_ (.o(regtop_dchdi_w1_hdi00[537]),
	.ck(clk),
	.d(n185628));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__26_ (.o(regtop_dchdi_w1_hdi00[538]),
	.ck(clk),
	.d(n185627));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__27_ (.o(regtop_dchdi_w1_hdi00[539]),
	.ck(clk),
	.d(n185626));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__28_ (.o(regtop_dchdi_w1_hdi00[540]),
	.ck(clk),
	.d(n185625));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__29_ (.o(regtop_dchdi_w1_hdi00[541]),
	.ck(clk),
	.d(n185624));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__30_ (.o(regtop_dchdi_w1_hdi00[542]),
	.ck(clk),
	.d(n185623));
   ms00f80 regtop_dchdi_w1_hdi00_reg_32__31_ (.o(regtop_dchdi_w1_hdi00[543]),
	.ck(clk),
	.d(n185622));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__0_ (.o(regtop_dchdi_w1_hdi00[544]),
	.ck(clk),
	.d(n185621));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__1_ (.o(regtop_dchdi_w1_hdi00[545]),
	.ck(clk),
	.d(n185620));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__2_ (.o(regtop_dchdi_w1_hdi00[546]),
	.ck(clk),
	.d(n185619));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__3_ (.o(regtop_dchdi_w1_hdi00[547]),
	.ck(clk),
	.d(n185618));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__4_ (.o(regtop_dchdi_w1_hdi00[548]),
	.ck(clk),
	.d(n185617));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__5_ (.o(regtop_dchdi_w1_hdi00[549]),
	.ck(clk),
	.d(n185616));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__6_ (.o(regtop_dchdi_w1_hdi00[550]),
	.ck(clk),
	.d(n185615));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__7_ (.o(regtop_dchdi_w1_hdi00[551]),
	.ck(clk),
	.d(n185614));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__8_ (.o(regtop_dchdi_w1_hdi00[552]),
	.ck(clk),
	.d(n185613));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__9_ (.o(regtop_dchdi_w1_hdi00[553]),
	.ck(clk),
	.d(n185612));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__10_ (.o(regtop_dchdi_w1_hdi00[554]),
	.ck(clk),
	.d(n185611));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__11_ (.o(regtop_dchdi_w1_hdi00[555]),
	.ck(clk),
	.d(n185610));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__12_ (.o(regtop_dchdi_w1_hdi00[556]),
	.ck(clk),
	.d(n185609));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__13_ (.o(regtop_dchdi_w1_hdi00[557]),
	.ck(clk),
	.d(n185608));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__14_ (.o(regtop_dchdi_w1_hdi00[558]),
	.ck(clk),
	.d(n185607));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__15_ (.o(regtop_dchdi_w1_hdi00[559]),
	.ck(clk),
	.d(n185606));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__16_ (.o(regtop_dchdi_w1_hdi00[560]),
	.ck(clk),
	.d(n185605));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__17_ (.o(regtop_dchdi_w1_hdi00[561]),
	.ck(clk),
	.d(n185604));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__18_ (.o(regtop_dchdi_w1_hdi00[562]),
	.ck(clk),
	.d(n185603));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__19_ (.o(regtop_dchdi_w1_hdi00[563]),
	.ck(clk),
	.d(n185602));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__20_ (.o(regtop_dchdi_w1_hdi00[564]),
	.ck(clk),
	.d(n185601));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__21_ (.o(regtop_dchdi_w1_hdi00[565]),
	.ck(clk),
	.d(n185600));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__22_ (.o(regtop_dchdi_w1_hdi00[566]),
	.ck(clk),
	.d(n185599));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__23_ (.o(regtop_dchdi_w1_hdi00[567]),
	.ck(clk),
	.d(n185598));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__24_ (.o(regtop_dchdi_w1_hdi00[568]),
	.ck(clk),
	.d(n185597));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__25_ (.o(regtop_dchdi_w1_hdi00[569]),
	.ck(clk),
	.d(n185596));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__26_ (.o(regtop_dchdi_w1_hdi00[570]),
	.ck(clk),
	.d(n185595));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__27_ (.o(regtop_dchdi_w1_hdi00[571]),
	.ck(clk),
	.d(n185594));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__28_ (.o(regtop_dchdi_w1_hdi00[572]),
	.ck(clk),
	.d(n185593));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__29_ (.o(regtop_dchdi_w1_hdi00[573]),
	.ck(clk),
	.d(n185592));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__30_ (.o(regtop_dchdi_w1_hdi00[574]),
	.ck(clk),
	.d(n185591));
   ms00f80 regtop_dchdi_w1_hdi00_reg_33__31_ (.o(regtop_dchdi_w1_hdi00[575]),
	.ck(clk),
	.d(n185590));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__0_ (.o(regtop_dchdi_w1_hdi00[576]),
	.ck(clk),
	.d(n185589));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__1_ (.o(regtop_dchdi_w1_hdi00[577]),
	.ck(clk),
	.d(n185588));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__2_ (.o(regtop_dchdi_w1_hdi00[578]),
	.ck(clk),
	.d(n185587));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__3_ (.o(regtop_dchdi_w1_hdi00[579]),
	.ck(clk),
	.d(n185586));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__4_ (.o(regtop_dchdi_w1_hdi00[580]),
	.ck(clk),
	.d(n185585));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__5_ (.o(regtop_dchdi_w1_hdi00[581]),
	.ck(clk),
	.d(n185584));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__6_ (.o(regtop_dchdi_w1_hdi00[582]),
	.ck(clk),
	.d(n185583));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__7_ (.o(regtop_dchdi_w1_hdi00[583]),
	.ck(clk),
	.d(n185582));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__8_ (.o(regtop_dchdi_w1_hdi00[584]),
	.ck(clk),
	.d(n185581));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__9_ (.o(regtop_dchdi_w1_hdi00[585]),
	.ck(clk),
	.d(n185580));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__10_ (.o(regtop_dchdi_w1_hdi00[586]),
	.ck(clk),
	.d(n185579));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__11_ (.o(regtop_dchdi_w1_hdi00[587]),
	.ck(clk),
	.d(n185578));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__12_ (.o(regtop_dchdi_w1_hdi00[588]),
	.ck(clk),
	.d(n185577));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__13_ (.o(regtop_dchdi_w1_hdi00[589]),
	.ck(clk),
	.d(n185576));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__14_ (.o(regtop_dchdi_w1_hdi00[590]),
	.ck(clk),
	.d(n185575));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__15_ (.o(regtop_dchdi_w1_hdi00[591]),
	.ck(clk),
	.d(n185574));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__16_ (.o(regtop_dchdi_w1_hdi00[592]),
	.ck(clk),
	.d(n185573));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__17_ (.o(regtop_dchdi_w1_hdi00[593]),
	.ck(clk),
	.d(n185572));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__18_ (.o(regtop_dchdi_w1_hdi00[594]),
	.ck(clk),
	.d(n185571));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__19_ (.o(regtop_dchdi_w1_hdi00[595]),
	.ck(clk),
	.d(n185570));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__20_ (.o(regtop_dchdi_w1_hdi00[596]),
	.ck(clk),
	.d(n185569));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__21_ (.o(regtop_dchdi_w1_hdi00[597]),
	.ck(clk),
	.d(n185568));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__22_ (.o(regtop_dchdi_w1_hdi00[598]),
	.ck(clk),
	.d(n185567));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__23_ (.o(regtop_dchdi_w1_hdi00[599]),
	.ck(clk),
	.d(n185566));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__24_ (.o(regtop_dchdi_w1_hdi00[600]),
	.ck(clk),
	.d(n185565));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__25_ (.o(regtop_dchdi_w1_hdi00[601]),
	.ck(clk),
	.d(n185564));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__26_ (.o(regtop_dchdi_w1_hdi00[602]),
	.ck(clk),
	.d(n185563));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__27_ (.o(regtop_dchdi_w1_hdi00[603]),
	.ck(clk),
	.d(n185562));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__28_ (.o(regtop_dchdi_w1_hdi00[604]),
	.ck(clk),
	.d(n185561));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__29_ (.o(regtop_dchdi_w1_hdi00[605]),
	.ck(clk),
	.d(n185560));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__30_ (.o(regtop_dchdi_w1_hdi00[606]),
	.ck(clk),
	.d(n185559));
   ms00f80 regtop_dchdi_w1_hdi00_reg_34__31_ (.o(regtop_dchdi_w1_hdi00[607]),
	.ck(clk),
	.d(n185558));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__0_ (.o(regtop_dchdi_w1_hdi00[608]),
	.ck(clk),
	.d(n185557));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__1_ (.o(regtop_dchdi_w1_hdi00[609]),
	.ck(clk),
	.d(n185556));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__2_ (.o(regtop_dchdi_w1_hdi00[610]),
	.ck(clk),
	.d(n185555));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__3_ (.o(regtop_dchdi_w1_hdi00[611]),
	.ck(clk),
	.d(n185554));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__4_ (.o(regtop_dchdi_w1_hdi00[612]),
	.ck(clk),
	.d(n185553));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__5_ (.o(regtop_dchdi_w1_hdi00[613]),
	.ck(clk),
	.d(n185552));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__6_ (.o(regtop_dchdi_w1_hdi00[614]),
	.ck(clk),
	.d(n185551));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__7_ (.o(regtop_dchdi_w1_hdi00[615]),
	.ck(clk),
	.d(n185550));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__8_ (.o(regtop_dchdi_w1_hdi00[616]),
	.ck(clk),
	.d(n185549));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__9_ (.o(regtop_dchdi_w1_hdi00[617]),
	.ck(clk),
	.d(n185548));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__10_ (.o(regtop_dchdi_w1_hdi00[618]),
	.ck(clk),
	.d(n185547));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__11_ (.o(regtop_dchdi_w1_hdi00[619]),
	.ck(clk),
	.d(n185546));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__12_ (.o(regtop_dchdi_w1_hdi00[620]),
	.ck(clk),
	.d(n185545));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__13_ (.o(regtop_dchdi_w1_hdi00[621]),
	.ck(clk),
	.d(n185544));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__14_ (.o(regtop_dchdi_w1_hdi00[622]),
	.ck(clk),
	.d(n185543));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__15_ (.o(regtop_dchdi_w1_hdi00[623]),
	.ck(clk),
	.d(n185542));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__16_ (.o(regtop_dchdi_w1_hdi00[624]),
	.ck(clk),
	.d(n185541));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__17_ (.o(regtop_dchdi_w1_hdi00[625]),
	.ck(clk),
	.d(n185540));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__18_ (.o(regtop_dchdi_w1_hdi00[626]),
	.ck(clk),
	.d(n185539));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__19_ (.o(regtop_dchdi_w1_hdi00[627]),
	.ck(clk),
	.d(n185538));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__20_ (.o(regtop_dchdi_w1_hdi00[628]),
	.ck(clk),
	.d(n185537));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__21_ (.o(regtop_dchdi_w1_hdi00[629]),
	.ck(clk),
	.d(n185536));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__22_ (.o(regtop_dchdi_w1_hdi00[630]),
	.ck(clk),
	.d(n185535));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__23_ (.o(regtop_dchdi_w1_hdi00[631]),
	.ck(clk),
	.d(n185534));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__24_ (.o(regtop_dchdi_w1_hdi00[632]),
	.ck(clk),
	.d(n185533));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__25_ (.o(regtop_dchdi_w1_hdi00[633]),
	.ck(clk),
	.d(n185532));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__26_ (.o(regtop_dchdi_w1_hdi00[634]),
	.ck(clk),
	.d(n185531));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__27_ (.o(regtop_dchdi_w1_hdi00[635]),
	.ck(clk),
	.d(n185530));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__28_ (.o(regtop_dchdi_w1_hdi00[636]),
	.ck(clk),
	.d(n185529));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__29_ (.o(regtop_dchdi_w1_hdi00[637]),
	.ck(clk),
	.d(n185528));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__30_ (.o(regtop_dchdi_w1_hdi00[638]),
	.ck(clk),
	.d(n185527));
   ms00f80 regtop_dchdi_w1_hdi00_reg_35__31_ (.o(regtop_dchdi_w1_hdi00[639]),
	.ck(clk),
	.d(n185526));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__0_ (.o(regtop_dchdi_w1_hdi00[640]),
	.ck(clk),
	.d(n185525));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__1_ (.o(regtop_dchdi_w1_hdi00[641]),
	.ck(clk),
	.d(n185524));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__2_ (.o(regtop_dchdi_w1_hdi00[642]),
	.ck(clk),
	.d(n185523));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__3_ (.o(regtop_dchdi_w1_hdi00[643]),
	.ck(clk),
	.d(n185522));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__4_ (.o(regtop_dchdi_w1_hdi00[644]),
	.ck(clk),
	.d(n185521));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__5_ (.o(regtop_dchdi_w1_hdi00[645]),
	.ck(clk),
	.d(n185520));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__6_ (.o(regtop_dchdi_w1_hdi00[646]),
	.ck(clk),
	.d(n185519));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__7_ (.o(regtop_dchdi_w1_hdi00[647]),
	.ck(clk),
	.d(n185518));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__8_ (.o(regtop_dchdi_w1_hdi00[648]),
	.ck(clk),
	.d(n185517));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__9_ (.o(regtop_dchdi_w1_hdi00[649]),
	.ck(clk),
	.d(n185516));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__10_ (.o(regtop_dchdi_w1_hdi00[650]),
	.ck(clk),
	.d(n185515));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__11_ (.o(regtop_dchdi_w1_hdi00[651]),
	.ck(clk),
	.d(n185514));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__12_ (.o(regtop_dchdi_w1_hdi00[652]),
	.ck(clk),
	.d(n185513));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__13_ (.o(regtop_dchdi_w1_hdi00[653]),
	.ck(clk),
	.d(n185512));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__14_ (.o(regtop_dchdi_w1_hdi00[654]),
	.ck(clk),
	.d(n185511));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__15_ (.o(regtop_dchdi_w1_hdi00[655]),
	.ck(clk),
	.d(n185510));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__16_ (.o(regtop_dchdi_w1_hdi00[656]),
	.ck(clk),
	.d(n185509));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__17_ (.o(regtop_dchdi_w1_hdi00[657]),
	.ck(clk),
	.d(n185508));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__18_ (.o(regtop_dchdi_w1_hdi00[658]),
	.ck(clk),
	.d(n185507));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__19_ (.o(regtop_dchdi_w1_hdi00[659]),
	.ck(clk),
	.d(n185506));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__20_ (.o(regtop_dchdi_w1_hdi00[660]),
	.ck(clk),
	.d(n185505));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__21_ (.o(regtop_dchdi_w1_hdi00[661]),
	.ck(clk),
	.d(n185504));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__22_ (.o(regtop_dchdi_w1_hdi00[662]),
	.ck(clk),
	.d(n185503));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__23_ (.o(regtop_dchdi_w1_hdi00[663]),
	.ck(clk),
	.d(n185502));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__24_ (.o(regtop_dchdi_w1_hdi00[664]),
	.ck(clk),
	.d(n185501));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__25_ (.o(regtop_dchdi_w1_hdi00[665]),
	.ck(clk),
	.d(n185500));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__26_ (.o(regtop_dchdi_w1_hdi00[666]),
	.ck(clk),
	.d(n185499));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__27_ (.o(regtop_dchdi_w1_hdi00[667]),
	.ck(clk),
	.d(n185498));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__28_ (.o(regtop_dchdi_w1_hdi00[668]),
	.ck(clk),
	.d(n185497));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__29_ (.o(regtop_dchdi_w1_hdi00[669]),
	.ck(clk),
	.d(n185496));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__30_ (.o(regtop_dchdi_w1_hdi00[670]),
	.ck(clk),
	.d(n185495));
   ms00f80 regtop_dchdi_w1_hdi00_reg_36__31_ (.o(regtop_dchdi_w1_hdi00[671]),
	.ck(clk),
	.d(n185494));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__0_ (.o(regtop_dchdi_w1_hdi00[672]),
	.ck(clk),
	.d(n185493));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__1_ (.o(regtop_dchdi_w1_hdi00[673]),
	.ck(clk),
	.d(n185492));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__2_ (.o(regtop_dchdi_w1_hdi00[674]),
	.ck(clk),
	.d(n185491));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__3_ (.o(regtop_dchdi_w1_hdi00[675]),
	.ck(clk),
	.d(n185490));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__4_ (.o(regtop_dchdi_w1_hdi00[676]),
	.ck(clk),
	.d(n185489));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__5_ (.o(regtop_dchdi_w1_hdi00[677]),
	.ck(clk),
	.d(n185488));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__6_ (.o(regtop_dchdi_w1_hdi00[678]),
	.ck(clk),
	.d(n185487));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__7_ (.o(regtop_dchdi_w1_hdi00[679]),
	.ck(clk),
	.d(n185486));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__8_ (.o(regtop_dchdi_w1_hdi00[680]),
	.ck(clk),
	.d(n185485));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__9_ (.o(regtop_dchdi_w1_hdi00[681]),
	.ck(clk),
	.d(n185484));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__10_ (.o(regtop_dchdi_w1_hdi00[682]),
	.ck(clk),
	.d(n185483));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__11_ (.o(regtop_dchdi_w1_hdi00[683]),
	.ck(clk),
	.d(n185482));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__12_ (.o(regtop_dchdi_w1_hdi00[684]),
	.ck(clk),
	.d(n185481));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__13_ (.o(regtop_dchdi_w1_hdi00[685]),
	.ck(clk),
	.d(n185480));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__14_ (.o(regtop_dchdi_w1_hdi00[686]),
	.ck(clk),
	.d(n185479));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__15_ (.o(regtop_dchdi_w1_hdi00[687]),
	.ck(clk),
	.d(n185478));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__16_ (.o(regtop_dchdi_w1_hdi00[688]),
	.ck(clk),
	.d(n185477));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__17_ (.o(regtop_dchdi_w1_hdi00[689]),
	.ck(clk),
	.d(n185476));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__18_ (.o(regtop_dchdi_w1_hdi00[690]),
	.ck(clk),
	.d(n185475));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__19_ (.o(regtop_dchdi_w1_hdi00[691]),
	.ck(clk),
	.d(n185474));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__20_ (.o(regtop_dchdi_w1_hdi00[692]),
	.ck(clk),
	.d(n185473));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__21_ (.o(regtop_dchdi_w1_hdi00[693]),
	.ck(clk),
	.d(n185472));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__22_ (.o(regtop_dchdi_w1_hdi00[694]),
	.ck(clk),
	.d(n185471));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__23_ (.o(regtop_dchdi_w1_hdi00[695]),
	.ck(clk),
	.d(n185470));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__24_ (.o(regtop_dchdi_w1_hdi00[696]),
	.ck(clk),
	.d(n185469));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__25_ (.o(regtop_dchdi_w1_hdi00[697]),
	.ck(clk),
	.d(n185468));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__26_ (.o(regtop_dchdi_w1_hdi00[698]),
	.ck(clk),
	.d(n185467));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__27_ (.o(regtop_dchdi_w1_hdi00[699]),
	.ck(clk),
	.d(n185466));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__28_ (.o(regtop_dchdi_w1_hdi00[700]),
	.ck(clk),
	.d(n185465));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__29_ (.o(regtop_dchdi_w1_hdi00[701]),
	.ck(clk),
	.d(n185464));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__30_ (.o(regtop_dchdi_w1_hdi00[702]),
	.ck(clk),
	.d(n185463));
   ms00f80 regtop_dchdi_w1_hdi00_reg_37__31_ (.o(regtop_dchdi_w1_hdi00[703]),
	.ck(clk),
	.d(n185462));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__0_ (.o(regtop_dchdi_w1_hdi00[704]),
	.ck(clk),
	.d(n185461));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__1_ (.o(regtop_dchdi_w1_hdi00[705]),
	.ck(clk),
	.d(n185460));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__2_ (.o(regtop_dchdi_w1_hdi00[706]),
	.ck(clk),
	.d(n185459));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__3_ (.o(regtop_dchdi_w1_hdi00[707]),
	.ck(clk),
	.d(n185458));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__4_ (.o(regtop_dchdi_w1_hdi00[708]),
	.ck(clk),
	.d(n185457));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__5_ (.o(regtop_dchdi_w1_hdi00[709]),
	.ck(clk),
	.d(n185456));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__6_ (.o(regtop_dchdi_w1_hdi00[710]),
	.ck(clk),
	.d(n185455));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__7_ (.o(regtop_dchdi_w1_hdi00[711]),
	.ck(clk),
	.d(n185454));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__8_ (.o(regtop_dchdi_w1_hdi00[712]),
	.ck(clk),
	.d(n185453));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__9_ (.o(regtop_dchdi_w1_hdi00[713]),
	.ck(clk),
	.d(n185452));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__10_ (.o(regtop_dchdi_w1_hdi00[714]),
	.ck(clk),
	.d(n185451));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__11_ (.o(regtop_dchdi_w1_hdi00[715]),
	.ck(clk),
	.d(n185450));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__12_ (.o(regtop_dchdi_w1_hdi00[716]),
	.ck(clk),
	.d(n185449));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__13_ (.o(regtop_dchdi_w1_hdi00[717]),
	.ck(clk),
	.d(n185448));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__14_ (.o(regtop_dchdi_w1_hdi00[718]),
	.ck(clk),
	.d(n185447));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__15_ (.o(regtop_dchdi_w1_hdi00[719]),
	.ck(clk),
	.d(n185446));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__16_ (.o(regtop_dchdi_w1_hdi00[720]),
	.ck(clk),
	.d(n185445));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__17_ (.o(regtop_dchdi_w1_hdi00[721]),
	.ck(clk),
	.d(n185444));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__18_ (.o(regtop_dchdi_w1_hdi00[722]),
	.ck(clk),
	.d(n185443));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__19_ (.o(regtop_dchdi_w1_hdi00[723]),
	.ck(clk),
	.d(n185442));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__20_ (.o(regtop_dchdi_w1_hdi00[724]),
	.ck(clk),
	.d(n185441));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__21_ (.o(regtop_dchdi_w1_hdi00[725]),
	.ck(clk),
	.d(n185440));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__22_ (.o(regtop_dchdi_w1_hdi00[726]),
	.ck(clk),
	.d(n185439));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__23_ (.o(regtop_dchdi_w1_hdi00[727]),
	.ck(clk),
	.d(n185438));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__24_ (.o(regtop_dchdi_w1_hdi00[728]),
	.ck(clk),
	.d(n185437));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__25_ (.o(regtop_dchdi_w1_hdi00[729]),
	.ck(clk),
	.d(n185436));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__26_ (.o(regtop_dchdi_w1_hdi00[730]),
	.ck(clk),
	.d(n185435));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__27_ (.o(regtop_dchdi_w1_hdi00[731]),
	.ck(clk),
	.d(n185434));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__28_ (.o(regtop_dchdi_w1_hdi00[732]),
	.ck(clk),
	.d(n185433));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__29_ (.o(regtop_dchdi_w1_hdi00[733]),
	.ck(clk),
	.d(n185432));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__30_ (.o(regtop_dchdi_w1_hdi00[734]),
	.ck(clk),
	.d(n185431));
   ms00f80 regtop_dchdi_w1_hdi00_reg_38__31_ (.o(regtop_dchdi_w1_hdi00[735]),
	.ck(clk),
	.d(n185430));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__0_ (.o(regtop_dchdi_w1_hdi00[736]),
	.ck(clk),
	.d(n185429));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__1_ (.o(regtop_dchdi_w1_hdi00[737]),
	.ck(clk),
	.d(n185428));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__2_ (.o(regtop_dchdi_w1_hdi00[738]),
	.ck(clk),
	.d(n185427));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__3_ (.o(regtop_dchdi_w1_hdi00[739]),
	.ck(clk),
	.d(n185426));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__4_ (.o(regtop_dchdi_w1_hdi00[740]),
	.ck(clk),
	.d(n185425));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__5_ (.o(regtop_dchdi_w1_hdi00[741]),
	.ck(clk),
	.d(n185424));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__6_ (.o(regtop_dchdi_w1_hdi00[742]),
	.ck(clk),
	.d(n185423));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__7_ (.o(regtop_dchdi_w1_hdi00[743]),
	.ck(clk),
	.d(n185422));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__8_ (.o(regtop_dchdi_w1_hdi00[744]),
	.ck(clk),
	.d(n185421));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__9_ (.o(regtop_dchdi_w1_hdi00[745]),
	.ck(clk),
	.d(n185420));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__10_ (.o(regtop_dchdi_w1_hdi00[746]),
	.ck(clk),
	.d(n185419));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__11_ (.o(regtop_dchdi_w1_hdi00[747]),
	.ck(clk),
	.d(n185418));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__12_ (.o(regtop_dchdi_w1_hdi00[748]),
	.ck(clk),
	.d(n185417));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__13_ (.o(regtop_dchdi_w1_hdi00[749]),
	.ck(clk),
	.d(n185416));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__14_ (.o(regtop_dchdi_w1_hdi00[750]),
	.ck(clk),
	.d(n185415));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__15_ (.o(regtop_dchdi_w1_hdi00[751]),
	.ck(clk),
	.d(n185414));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__16_ (.o(regtop_dchdi_w1_hdi00[752]),
	.ck(clk),
	.d(n185413));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__17_ (.o(regtop_dchdi_w1_hdi00[753]),
	.ck(clk),
	.d(n185412));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__18_ (.o(regtop_dchdi_w1_hdi00[754]),
	.ck(clk),
	.d(n185411));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__19_ (.o(regtop_dchdi_w1_hdi00[755]),
	.ck(clk),
	.d(n185410));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__20_ (.o(regtop_dchdi_w1_hdi00[756]),
	.ck(clk),
	.d(n185409));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__21_ (.o(regtop_dchdi_w1_hdi00[757]),
	.ck(clk),
	.d(n185408));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__22_ (.o(regtop_dchdi_w1_hdi00[758]),
	.ck(clk),
	.d(n185407));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__23_ (.o(regtop_dchdi_w1_hdi00[759]),
	.ck(clk),
	.d(n185406));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__24_ (.o(regtop_dchdi_w1_hdi00[760]),
	.ck(clk),
	.d(n185405));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__25_ (.o(regtop_dchdi_w1_hdi00[761]),
	.ck(clk),
	.d(n185404));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__26_ (.o(regtop_dchdi_w1_hdi00[762]),
	.ck(clk),
	.d(n185403));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__27_ (.o(regtop_dchdi_w1_hdi00[763]),
	.ck(clk),
	.d(n185402));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__28_ (.o(regtop_dchdi_w1_hdi00[764]),
	.ck(clk),
	.d(n185401));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__29_ (.o(regtop_dchdi_w1_hdi00[765]),
	.ck(clk),
	.d(n185400));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__30_ (.o(regtop_dchdi_w1_hdi00[766]),
	.ck(clk),
	.d(n185399));
   ms00f80 regtop_dchdi_w1_hdi00_reg_39__31_ (.o(regtop_dchdi_w1_hdi00[767]),
	.ck(clk),
	.d(n185398));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__0_ (.o(regtop_dchdi_w1_hdi00[768]),
	.ck(clk),
	.d(n185397));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__1_ (.o(regtop_dchdi_w1_hdi00[769]),
	.ck(clk),
	.d(n185396));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__2_ (.o(regtop_dchdi_w1_hdi00[770]),
	.ck(clk),
	.d(n185395));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__3_ (.o(regtop_dchdi_w1_hdi00[771]),
	.ck(clk),
	.d(n185394));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__4_ (.o(regtop_dchdi_w1_hdi00[772]),
	.ck(clk),
	.d(n185393));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__5_ (.o(regtop_dchdi_w1_hdi00[773]),
	.ck(clk),
	.d(n185392));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__6_ (.o(regtop_dchdi_w1_hdi00[774]),
	.ck(clk),
	.d(n185391));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__7_ (.o(regtop_dchdi_w1_hdi00[775]),
	.ck(clk),
	.d(n185390));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__8_ (.o(regtop_dchdi_w1_hdi00[776]),
	.ck(clk),
	.d(n185389));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__9_ (.o(regtop_dchdi_w1_hdi00[777]),
	.ck(clk),
	.d(n185388));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__10_ (.o(regtop_dchdi_w1_hdi00[778]),
	.ck(clk),
	.d(n185387));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__11_ (.o(regtop_dchdi_w1_hdi00[779]),
	.ck(clk),
	.d(n185386));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__12_ (.o(regtop_dchdi_w1_hdi00[780]),
	.ck(clk),
	.d(n185385));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__13_ (.o(regtop_dchdi_w1_hdi00[781]),
	.ck(clk),
	.d(n185384));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__14_ (.o(regtop_dchdi_w1_hdi00[782]),
	.ck(clk),
	.d(n185383));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__15_ (.o(regtop_dchdi_w1_hdi00[783]),
	.ck(clk),
	.d(n185382));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__16_ (.o(regtop_dchdi_w1_hdi00[784]),
	.ck(clk),
	.d(n185381));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__17_ (.o(regtop_dchdi_w1_hdi00[785]),
	.ck(clk),
	.d(n185380));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__18_ (.o(regtop_dchdi_w1_hdi00[786]),
	.ck(clk),
	.d(n185379));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__19_ (.o(regtop_dchdi_w1_hdi00[787]),
	.ck(clk),
	.d(n185378));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__20_ (.o(regtop_dchdi_w1_hdi00[788]),
	.ck(clk),
	.d(n185377));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__21_ (.o(regtop_dchdi_w1_hdi00[789]),
	.ck(clk),
	.d(n185376));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__22_ (.o(regtop_dchdi_w1_hdi00[790]),
	.ck(clk),
	.d(n185375));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__23_ (.o(regtop_dchdi_w1_hdi00[791]),
	.ck(clk),
	.d(n185374));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__24_ (.o(regtop_dchdi_w1_hdi00[792]),
	.ck(clk),
	.d(n185373));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__25_ (.o(regtop_dchdi_w1_hdi00[793]),
	.ck(clk),
	.d(n185372));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__26_ (.o(regtop_dchdi_w1_hdi00[794]),
	.ck(clk),
	.d(n185371));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__27_ (.o(regtop_dchdi_w1_hdi00[795]),
	.ck(clk),
	.d(n185370));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__28_ (.o(regtop_dchdi_w1_hdi00[796]),
	.ck(clk),
	.d(n185369));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__29_ (.o(regtop_dchdi_w1_hdi00[797]),
	.ck(clk),
	.d(n185368));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__30_ (.o(regtop_dchdi_w1_hdi00[798]),
	.ck(clk),
	.d(n185367));
   ms00f80 regtop_dchdi_w1_hdi00_reg_40__31_ (.o(regtop_dchdi_w1_hdi00[799]),
	.ck(clk),
	.d(n185366));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__0_ (.o(regtop_dchdi_w1_hdi00[800]),
	.ck(clk),
	.d(n185365));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__1_ (.o(regtop_dchdi_w1_hdi00[801]),
	.ck(clk),
	.d(n185364));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__2_ (.o(regtop_dchdi_w1_hdi00[802]),
	.ck(clk),
	.d(n185363));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__3_ (.o(regtop_dchdi_w1_hdi00[803]),
	.ck(clk),
	.d(n185362));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__4_ (.o(regtop_dchdi_w1_hdi00[804]),
	.ck(clk),
	.d(n185361));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__5_ (.o(regtop_dchdi_w1_hdi00[805]),
	.ck(clk),
	.d(n185360));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__6_ (.o(regtop_dchdi_w1_hdi00[806]),
	.ck(clk),
	.d(n185359));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__7_ (.o(regtop_dchdi_w1_hdi00[807]),
	.ck(clk),
	.d(n185358));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__8_ (.o(regtop_dchdi_w1_hdi00[808]),
	.ck(clk),
	.d(n185357));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__9_ (.o(regtop_dchdi_w1_hdi00[809]),
	.ck(clk),
	.d(n185356));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__10_ (.o(regtop_dchdi_w1_hdi00[810]),
	.ck(clk),
	.d(n185355));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__11_ (.o(regtop_dchdi_w1_hdi00[811]),
	.ck(clk),
	.d(n185354));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__12_ (.o(regtop_dchdi_w1_hdi00[812]),
	.ck(clk),
	.d(n185353));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__13_ (.o(regtop_dchdi_w1_hdi00[813]),
	.ck(clk),
	.d(n185352));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__14_ (.o(regtop_dchdi_w1_hdi00[814]),
	.ck(clk),
	.d(n185351));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__15_ (.o(regtop_dchdi_w1_hdi00[815]),
	.ck(clk),
	.d(n185350));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__16_ (.o(regtop_dchdi_w1_hdi00[816]),
	.ck(clk),
	.d(n185349));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__17_ (.o(regtop_dchdi_w1_hdi00[817]),
	.ck(clk),
	.d(n185348));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__18_ (.o(regtop_dchdi_w1_hdi00[818]),
	.ck(clk),
	.d(n185347));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__19_ (.o(regtop_dchdi_w1_hdi00[819]),
	.ck(clk),
	.d(n185346));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__20_ (.o(regtop_dchdi_w1_hdi00[820]),
	.ck(clk),
	.d(n185345));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__21_ (.o(regtop_dchdi_w1_hdi00[821]),
	.ck(clk),
	.d(n185344));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__22_ (.o(regtop_dchdi_w1_hdi00[822]),
	.ck(clk),
	.d(n185343));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__23_ (.o(regtop_dchdi_w1_hdi00[823]),
	.ck(clk),
	.d(n185342));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__24_ (.o(regtop_dchdi_w1_hdi00[824]),
	.ck(clk),
	.d(n185341));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__25_ (.o(regtop_dchdi_w1_hdi00[825]),
	.ck(clk),
	.d(n185340));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__26_ (.o(regtop_dchdi_w1_hdi00[826]),
	.ck(clk),
	.d(n185339));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__27_ (.o(regtop_dchdi_w1_hdi00[827]),
	.ck(clk),
	.d(n185338));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__28_ (.o(regtop_dchdi_w1_hdi00[828]),
	.ck(clk),
	.d(n185337));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__29_ (.o(regtop_dchdi_w1_hdi00[829]),
	.ck(clk),
	.d(n185336));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__30_ (.o(regtop_dchdi_w1_hdi00[830]),
	.ck(clk),
	.d(n185335));
   ms00f80 regtop_dchdi_w1_hdi00_reg_41__31_ (.o(regtop_dchdi_w1_hdi00[831]),
	.ck(clk),
	.d(n185334));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__0_ (.o(regtop_dchdi_w1_hdi00[832]),
	.ck(clk),
	.d(n185333));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__1_ (.o(regtop_dchdi_w1_hdi00[833]),
	.ck(clk),
	.d(n185332));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__2_ (.o(regtop_dchdi_w1_hdi00[834]),
	.ck(clk),
	.d(n185331));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__3_ (.o(regtop_dchdi_w1_hdi00[835]),
	.ck(clk),
	.d(n185330));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__4_ (.o(regtop_dchdi_w1_hdi00[836]),
	.ck(clk),
	.d(n185329));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__5_ (.o(regtop_dchdi_w1_hdi00[837]),
	.ck(clk),
	.d(n185328));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__6_ (.o(regtop_dchdi_w1_hdi00[838]),
	.ck(clk),
	.d(n185327));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__7_ (.o(regtop_dchdi_w1_hdi00[839]),
	.ck(clk),
	.d(n185326));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__8_ (.o(regtop_dchdi_w1_hdi00[840]),
	.ck(clk),
	.d(n185325));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__9_ (.o(regtop_dchdi_w1_hdi00[841]),
	.ck(clk),
	.d(n185324));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__10_ (.o(regtop_dchdi_w1_hdi00[842]),
	.ck(clk),
	.d(n185323));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__11_ (.o(regtop_dchdi_w1_hdi00[843]),
	.ck(clk),
	.d(n185322));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__12_ (.o(regtop_dchdi_w1_hdi00[844]),
	.ck(clk),
	.d(n185321));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__13_ (.o(regtop_dchdi_w1_hdi00[845]),
	.ck(clk),
	.d(n185320));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__14_ (.o(regtop_dchdi_w1_hdi00[846]),
	.ck(clk),
	.d(n185319));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__15_ (.o(regtop_dchdi_w1_hdi00[847]),
	.ck(clk),
	.d(n185318));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__16_ (.o(regtop_dchdi_w1_hdi00[848]),
	.ck(clk),
	.d(n185317));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__17_ (.o(regtop_dchdi_w1_hdi00[849]),
	.ck(clk),
	.d(n185316));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__18_ (.o(regtop_dchdi_w1_hdi00[850]),
	.ck(clk),
	.d(n185315));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__19_ (.o(regtop_dchdi_w1_hdi00[851]),
	.ck(clk),
	.d(n185314));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__20_ (.o(regtop_dchdi_w1_hdi00[852]),
	.ck(clk),
	.d(n185313));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__21_ (.o(regtop_dchdi_w1_hdi00[853]),
	.ck(clk),
	.d(n185312));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__22_ (.o(regtop_dchdi_w1_hdi00[854]),
	.ck(clk),
	.d(n185311));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__23_ (.o(regtop_dchdi_w1_hdi00[855]),
	.ck(clk),
	.d(n185310));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__24_ (.o(regtop_dchdi_w1_hdi00[856]),
	.ck(clk),
	.d(n185309));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__25_ (.o(regtop_dchdi_w1_hdi00[857]),
	.ck(clk),
	.d(n185308));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__26_ (.o(regtop_dchdi_w1_hdi00[858]),
	.ck(clk),
	.d(n185307));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__27_ (.o(regtop_dchdi_w1_hdi00[859]),
	.ck(clk),
	.d(n185306));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__28_ (.o(regtop_dchdi_w1_hdi00[860]),
	.ck(clk),
	.d(n185305));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__29_ (.o(regtop_dchdi_w1_hdi00[861]),
	.ck(clk),
	.d(n185304));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__30_ (.o(regtop_dchdi_w1_hdi00[862]),
	.ck(clk),
	.d(n185303));
   ms00f80 regtop_dchdi_w1_hdi00_reg_42__31_ (.o(regtop_dchdi_w1_hdi00[863]),
	.ck(clk),
	.d(n185302));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__0_ (.o(regtop_dchdi_w1_hdi00[864]),
	.ck(clk),
	.d(n185301));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__1_ (.o(regtop_dchdi_w1_hdi00[865]),
	.ck(clk),
	.d(n185300));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__2_ (.o(regtop_dchdi_w1_hdi00[866]),
	.ck(clk),
	.d(n185299));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__3_ (.o(regtop_dchdi_w1_hdi00[867]),
	.ck(clk),
	.d(n185298));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__4_ (.o(regtop_dchdi_w1_hdi00[868]),
	.ck(clk),
	.d(n185297));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__5_ (.o(regtop_dchdi_w1_hdi00[869]),
	.ck(clk),
	.d(n185296));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__6_ (.o(regtop_dchdi_w1_hdi00[870]),
	.ck(clk),
	.d(n185295));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__7_ (.o(regtop_dchdi_w1_hdi00[871]),
	.ck(clk),
	.d(n185294));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__8_ (.o(regtop_dchdi_w1_hdi00[872]),
	.ck(clk),
	.d(n185293));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__9_ (.o(regtop_dchdi_w1_hdi00[873]),
	.ck(clk),
	.d(n185292));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__10_ (.o(regtop_dchdi_w1_hdi00[874]),
	.ck(clk),
	.d(n185291));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__11_ (.o(regtop_dchdi_w1_hdi00[875]),
	.ck(clk),
	.d(n185290));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__12_ (.o(regtop_dchdi_w1_hdi00[876]),
	.ck(clk),
	.d(n185289));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__13_ (.o(regtop_dchdi_w1_hdi00[877]),
	.ck(clk),
	.d(n185288));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__14_ (.o(regtop_dchdi_w1_hdi00[878]),
	.ck(clk),
	.d(n185287));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__15_ (.o(regtop_dchdi_w1_hdi00[879]),
	.ck(clk),
	.d(n185286));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__16_ (.o(regtop_dchdi_w1_hdi00[880]),
	.ck(clk),
	.d(n185285));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__17_ (.o(regtop_dchdi_w1_hdi00[881]),
	.ck(clk),
	.d(n185284));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__18_ (.o(regtop_dchdi_w1_hdi00[882]),
	.ck(clk),
	.d(n185283));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__19_ (.o(regtop_dchdi_w1_hdi00[883]),
	.ck(clk),
	.d(n185282));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__20_ (.o(regtop_dchdi_w1_hdi00[884]),
	.ck(clk),
	.d(n185281));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__21_ (.o(regtop_dchdi_w1_hdi00[885]),
	.ck(clk),
	.d(n185280));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__22_ (.o(regtop_dchdi_w1_hdi00[886]),
	.ck(clk),
	.d(n185279));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__23_ (.o(regtop_dchdi_w1_hdi00[887]),
	.ck(clk),
	.d(n185278));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__24_ (.o(regtop_dchdi_w1_hdi00[888]),
	.ck(clk),
	.d(n185277));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__25_ (.o(regtop_dchdi_w1_hdi00[889]),
	.ck(clk),
	.d(n185276));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__26_ (.o(regtop_dchdi_w1_hdi00[890]),
	.ck(clk),
	.d(n185275));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__27_ (.o(regtop_dchdi_w1_hdi00[891]),
	.ck(clk),
	.d(n185274));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__28_ (.o(regtop_dchdi_w1_hdi00[892]),
	.ck(clk),
	.d(n185273));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__29_ (.o(regtop_dchdi_w1_hdi00[893]),
	.ck(clk),
	.d(n185272));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__30_ (.o(regtop_dchdi_w1_hdi00[894]),
	.ck(clk),
	.d(n185271));
   ms00f80 regtop_dchdi_w1_hdi00_reg_43__31_ (.o(regtop_dchdi_w1_hdi00[895]),
	.ck(clk),
	.d(n185270));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__0_ (.o(regtop_dchdi_w1_hdi00[896]),
	.ck(clk),
	.d(n185269));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__1_ (.o(regtop_dchdi_w1_hdi00[897]),
	.ck(clk),
	.d(n185268));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__2_ (.o(regtop_dchdi_w1_hdi00[898]),
	.ck(clk),
	.d(n185267));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__3_ (.o(regtop_dchdi_w1_hdi00[899]),
	.ck(clk),
	.d(n185266));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__4_ (.o(regtop_dchdi_w1_hdi00[900]),
	.ck(clk),
	.d(n185265));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__5_ (.o(regtop_dchdi_w1_hdi00[901]),
	.ck(clk),
	.d(n185264));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__6_ (.o(regtop_dchdi_w1_hdi00[902]),
	.ck(clk),
	.d(n185263));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__7_ (.o(regtop_dchdi_w1_hdi00[903]),
	.ck(clk),
	.d(n185262));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__8_ (.o(regtop_dchdi_w1_hdi00[904]),
	.ck(clk),
	.d(n185261));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__9_ (.o(regtop_dchdi_w1_hdi00[905]),
	.ck(clk),
	.d(n185260));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__10_ (.o(regtop_dchdi_w1_hdi00[906]),
	.ck(clk),
	.d(n185259));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__11_ (.o(regtop_dchdi_w1_hdi00[907]),
	.ck(clk),
	.d(n185258));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__12_ (.o(regtop_dchdi_w1_hdi00[908]),
	.ck(clk),
	.d(n185257));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__13_ (.o(regtop_dchdi_w1_hdi00[909]),
	.ck(clk),
	.d(n185256));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__14_ (.o(regtop_dchdi_w1_hdi00[910]),
	.ck(clk),
	.d(n185255));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__15_ (.o(regtop_dchdi_w1_hdi00[911]),
	.ck(clk),
	.d(n185254));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__16_ (.o(regtop_dchdi_w1_hdi00[912]),
	.ck(clk),
	.d(n185253));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__17_ (.o(regtop_dchdi_w1_hdi00[913]),
	.ck(clk),
	.d(n185252));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__18_ (.o(regtop_dchdi_w1_hdi00[914]),
	.ck(clk),
	.d(n185251));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__19_ (.o(regtop_dchdi_w1_hdi00[915]),
	.ck(clk),
	.d(n185250));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__20_ (.o(regtop_dchdi_w1_hdi00[916]),
	.ck(clk),
	.d(n185249));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__21_ (.o(regtop_dchdi_w1_hdi00[917]),
	.ck(clk),
	.d(n185248));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__22_ (.o(regtop_dchdi_w1_hdi00[918]),
	.ck(clk),
	.d(n185247));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__23_ (.o(regtop_dchdi_w1_hdi00[919]),
	.ck(clk),
	.d(n185246));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__24_ (.o(regtop_dchdi_w1_hdi00[920]),
	.ck(clk),
	.d(n185245));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__25_ (.o(regtop_dchdi_w1_hdi00[921]),
	.ck(clk),
	.d(n185244));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__26_ (.o(regtop_dchdi_w1_hdi00[922]),
	.ck(clk),
	.d(n185243));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__27_ (.o(regtop_dchdi_w1_hdi00[923]),
	.ck(clk),
	.d(n185242));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__28_ (.o(regtop_dchdi_w1_hdi00[924]),
	.ck(clk),
	.d(n185241));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__29_ (.o(regtop_dchdi_w1_hdi00[925]),
	.ck(clk),
	.d(n185240));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__30_ (.o(regtop_dchdi_w1_hdi00[926]),
	.ck(clk),
	.d(n185239));
   ms00f80 regtop_dchdi_w1_hdi00_reg_44__31_ (.o(regtop_dchdi_w1_hdi00[927]),
	.ck(clk),
	.d(n185238));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__0_ (.o(regtop_dchdi_w1_hdi00[928]),
	.ck(clk),
	.d(n185237));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__1_ (.o(regtop_dchdi_w1_hdi00[929]),
	.ck(clk),
	.d(n185236));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__2_ (.o(regtop_dchdi_w1_hdi00[930]),
	.ck(clk),
	.d(n185235));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__3_ (.o(regtop_dchdi_w1_hdi00[931]),
	.ck(clk),
	.d(n185234));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__4_ (.o(regtop_dchdi_w1_hdi00[932]),
	.ck(clk),
	.d(n185233));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__5_ (.o(regtop_dchdi_w1_hdi00[933]),
	.ck(clk),
	.d(n185232));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__6_ (.o(regtop_dchdi_w1_hdi00[934]),
	.ck(clk),
	.d(n185231));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__7_ (.o(regtop_dchdi_w1_hdi00[935]),
	.ck(clk),
	.d(n185230));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__8_ (.o(regtop_dchdi_w1_hdi00[936]),
	.ck(clk),
	.d(n185229));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__9_ (.o(regtop_dchdi_w1_hdi00[937]),
	.ck(clk),
	.d(n185228));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__10_ (.o(regtop_dchdi_w1_hdi00[938]),
	.ck(clk),
	.d(n185227));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__11_ (.o(regtop_dchdi_w1_hdi00[939]),
	.ck(clk),
	.d(n185226));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__12_ (.o(regtop_dchdi_w1_hdi00[940]),
	.ck(clk),
	.d(n185225));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__13_ (.o(regtop_dchdi_w1_hdi00[941]),
	.ck(clk),
	.d(n185224));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__14_ (.o(regtop_dchdi_w1_hdi00[942]),
	.ck(clk),
	.d(n185223));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__15_ (.o(regtop_dchdi_w1_hdi00[943]),
	.ck(clk),
	.d(n185222));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__16_ (.o(regtop_dchdi_w1_hdi00[944]),
	.ck(clk),
	.d(n185221));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__17_ (.o(regtop_dchdi_w1_hdi00[945]),
	.ck(clk),
	.d(n185220));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__18_ (.o(regtop_dchdi_w1_hdi00[946]),
	.ck(clk),
	.d(n185219));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__19_ (.o(regtop_dchdi_w1_hdi00[947]),
	.ck(clk),
	.d(n185218));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__20_ (.o(regtop_dchdi_w1_hdi00[948]),
	.ck(clk),
	.d(n185217));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__21_ (.o(regtop_dchdi_w1_hdi00[949]),
	.ck(clk),
	.d(n185216));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__22_ (.o(regtop_dchdi_w1_hdi00[950]),
	.ck(clk),
	.d(n185215));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__23_ (.o(regtop_dchdi_w1_hdi00[951]),
	.ck(clk),
	.d(n185214));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__24_ (.o(regtop_dchdi_w1_hdi00[952]),
	.ck(clk),
	.d(n185213));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__25_ (.o(regtop_dchdi_w1_hdi00[953]),
	.ck(clk),
	.d(n185212));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__26_ (.o(regtop_dchdi_w1_hdi00[954]),
	.ck(clk),
	.d(n185211));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__27_ (.o(regtop_dchdi_w1_hdi00[955]),
	.ck(clk),
	.d(n185210));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__28_ (.o(regtop_dchdi_w1_hdi00[956]),
	.ck(clk),
	.d(n185209));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__29_ (.o(regtop_dchdi_w1_hdi00[957]),
	.ck(clk),
	.d(n185208));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__30_ (.o(regtop_dchdi_w1_hdi00[958]),
	.ck(clk),
	.d(n185207));
   ms00f80 regtop_dchdi_w1_hdi00_reg_45__31_ (.o(regtop_dchdi_w1_hdi00[959]),
	.ck(clk),
	.d(n185206));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__0_ (.o(regtop_dchdi_w1_hdi00[960]),
	.ck(clk),
	.d(n185205));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__1_ (.o(regtop_dchdi_w1_hdi00[961]),
	.ck(clk),
	.d(n185204));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__2_ (.o(regtop_dchdi_w1_hdi00[962]),
	.ck(clk),
	.d(n185203));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__3_ (.o(regtop_dchdi_w1_hdi00[963]),
	.ck(clk),
	.d(n185202));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__4_ (.o(regtop_dchdi_w1_hdi00[964]),
	.ck(clk),
	.d(n185201));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__5_ (.o(regtop_dchdi_w1_hdi00[965]),
	.ck(clk),
	.d(n185200));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__6_ (.o(regtop_dchdi_w1_hdi00[966]),
	.ck(clk),
	.d(n185199));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__7_ (.o(regtop_dchdi_w1_hdi00[967]),
	.ck(clk),
	.d(n185198));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__8_ (.o(regtop_dchdi_w1_hdi00[968]),
	.ck(clk),
	.d(n185197));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__9_ (.o(regtop_dchdi_w1_hdi00[969]),
	.ck(clk),
	.d(n185196));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__10_ (.o(regtop_dchdi_w1_hdi00[970]),
	.ck(clk),
	.d(n185195));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__11_ (.o(regtop_dchdi_w1_hdi00[971]),
	.ck(clk),
	.d(n185194));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__12_ (.o(regtop_dchdi_w1_hdi00[972]),
	.ck(clk),
	.d(n185193));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__13_ (.o(regtop_dchdi_w1_hdi00[973]),
	.ck(clk),
	.d(n185192));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__14_ (.o(regtop_dchdi_w1_hdi00[974]),
	.ck(clk),
	.d(n185191));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__15_ (.o(regtop_dchdi_w1_hdi00[975]),
	.ck(clk),
	.d(n185190));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__16_ (.o(regtop_dchdi_w1_hdi00[976]),
	.ck(clk),
	.d(n185189));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__17_ (.o(regtop_dchdi_w1_hdi00[977]),
	.ck(clk),
	.d(n185188));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__18_ (.o(regtop_dchdi_w1_hdi00[978]),
	.ck(clk),
	.d(n185187));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__19_ (.o(regtop_dchdi_w1_hdi00[979]),
	.ck(clk),
	.d(n185186));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__20_ (.o(regtop_dchdi_w1_hdi00[980]),
	.ck(clk),
	.d(n185185));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__21_ (.o(regtop_dchdi_w1_hdi00[981]),
	.ck(clk),
	.d(n185184));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__22_ (.o(regtop_dchdi_w1_hdi00[982]),
	.ck(clk),
	.d(n185183));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__23_ (.o(regtop_dchdi_w1_hdi00[983]),
	.ck(clk),
	.d(n185182));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__24_ (.o(regtop_dchdi_w1_hdi00[984]),
	.ck(clk),
	.d(n185181));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__25_ (.o(regtop_dchdi_w1_hdi00[985]),
	.ck(clk),
	.d(n185180));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__26_ (.o(regtop_dchdi_w1_hdi00[986]),
	.ck(clk),
	.d(n185179));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__27_ (.o(regtop_dchdi_w1_hdi00[987]),
	.ck(clk),
	.d(n185178));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__28_ (.o(regtop_dchdi_w1_hdi00[988]),
	.ck(clk),
	.d(n185177));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__29_ (.o(regtop_dchdi_w1_hdi00[989]),
	.ck(clk),
	.d(n185176));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__30_ (.o(regtop_dchdi_w1_hdi00[990]),
	.ck(clk),
	.d(n185175));
   ms00f80 regtop_dchdi_w1_hdi00_reg_46__31_ (.o(regtop_dchdi_w1_hdi00[991]),
	.ck(clk),
	.d(n185174));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__0_ (.o(regtop_dchdi_w1_hdi00[992]),
	.ck(clk),
	.d(n185173));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__1_ (.o(regtop_dchdi_w1_hdi00[993]),
	.ck(clk),
	.d(n185172));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__2_ (.o(regtop_dchdi_w1_hdi00[994]),
	.ck(clk),
	.d(n185171));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__3_ (.o(regtop_dchdi_w1_hdi00[995]),
	.ck(clk),
	.d(n185170));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__4_ (.o(regtop_dchdi_w1_hdi00[996]),
	.ck(clk),
	.d(n185169));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__5_ (.o(regtop_dchdi_w1_hdi00[997]),
	.ck(clk),
	.d(n185168));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__6_ (.o(regtop_dchdi_w1_hdi00[998]),
	.ck(clk),
	.d(n185167));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__7_ (.o(regtop_dchdi_w1_hdi00[999]),
	.ck(clk),
	.d(n185166));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__8_ (.o(regtop_dchdi_w1_hdi00[1000]),
	.ck(clk),
	.d(n185165));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__9_ (.o(regtop_dchdi_w1_hdi00[1001]),
	.ck(clk),
	.d(n185164));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__10_ (.o(regtop_dchdi_w1_hdi00[1002]),
	.ck(clk),
	.d(n185163));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__11_ (.o(regtop_dchdi_w1_hdi00[1003]),
	.ck(clk),
	.d(n185162));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__12_ (.o(regtop_dchdi_w1_hdi00[1004]),
	.ck(clk),
	.d(n185161));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__13_ (.o(regtop_dchdi_w1_hdi00[1005]),
	.ck(clk),
	.d(n185160));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__14_ (.o(regtop_dchdi_w1_hdi00[1006]),
	.ck(clk),
	.d(n185159));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__15_ (.o(regtop_dchdi_w1_hdi00[1007]),
	.ck(clk),
	.d(n185158));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__16_ (.o(regtop_dchdi_w1_hdi00[1008]),
	.ck(clk),
	.d(n185157));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__17_ (.o(regtop_dchdi_w1_hdi00[1009]),
	.ck(clk),
	.d(n185156));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__18_ (.o(regtop_dchdi_w1_hdi00[1010]),
	.ck(clk),
	.d(n185155));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__19_ (.o(regtop_dchdi_w1_hdi00[1011]),
	.ck(clk),
	.d(n185154));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__20_ (.o(regtop_dchdi_w1_hdi00[1012]),
	.ck(clk),
	.d(n185153));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__21_ (.o(regtop_dchdi_w1_hdi00[1013]),
	.ck(clk),
	.d(n185152));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__22_ (.o(regtop_dchdi_w1_hdi00[1014]),
	.ck(clk),
	.d(n185151));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__23_ (.o(regtop_dchdi_w1_hdi00[1015]),
	.ck(clk),
	.d(n185150));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__24_ (.o(regtop_dchdi_w1_hdi00[1016]),
	.ck(clk),
	.d(n185149));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__25_ (.o(regtop_dchdi_w1_hdi00[1017]),
	.ck(clk),
	.d(n185148));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__26_ (.o(regtop_dchdi_w1_hdi00[1018]),
	.ck(clk),
	.d(n185147));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__27_ (.o(regtop_dchdi_w1_hdi00[1019]),
	.ck(clk),
	.d(n185146));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__28_ (.o(regtop_dchdi_w1_hdi00[1020]),
	.ck(clk),
	.d(n185145));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__29_ (.o(regtop_dchdi_w1_hdi00[1021]),
	.ck(clk),
	.d(n185144));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__30_ (.o(regtop_dchdi_w1_hdi00[1022]),
	.ck(clk),
	.d(n185143));
   ms00f80 regtop_dchdi_w1_hdi00_reg_47__31_ (.o(regtop_dchdi_w1_hdi00[1023]),
	.ck(clk),
	.d(n185142));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__0_ (.o(regtop_dchdi_w1_hdi00[0]),
	.ck(clk),
	.d(n185141));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__1_ (.o(regtop_dchdi_w1_hdi00[1]),
	.ck(clk),
	.d(n185140));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__2_ (.o(regtop_dchdi_w1_hdi00[2]),
	.ck(clk),
	.d(n185139));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__3_ (.o(regtop_dchdi_w1_hdi00[3]),
	.ck(clk),
	.d(n185138));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__4_ (.o(regtop_dchdi_w1_hdi00[4]),
	.ck(clk),
	.d(n185137));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__5_ (.o(regtop_dchdi_w1_hdi00[5]),
	.ck(clk),
	.d(n185136));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__6_ (.o(regtop_dchdi_w1_hdi00[6]),
	.ck(clk),
	.d(n185135));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__7_ (.o(regtop_dchdi_w1_hdi00[7]),
	.ck(clk),
	.d(n185134));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__8_ (.o(regtop_dchdi_w1_hdi00[8]),
	.ck(clk),
	.d(n185133));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__9_ (.o(regtop_dchdi_w1_hdi00[9]),
	.ck(clk),
	.d(n185132));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__10_ (.o(regtop_dchdi_w1_hdi00[10]),
	.ck(clk),
	.d(n185131));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__11_ (.o(regtop_dchdi_w1_hdi00[11]),
	.ck(clk),
	.d(n185130));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__12_ (.o(regtop_dchdi_w1_hdi00[12]),
	.ck(clk),
	.d(n185129));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__13_ (.o(regtop_dchdi_w1_hdi00[13]),
	.ck(clk),
	.d(n185128));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__14_ (.o(regtop_dchdi_w1_hdi00[14]),
	.ck(clk),
	.d(n185127));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__15_ (.o(regtop_dchdi_w1_hdi00[15]),
	.ck(clk),
	.d(n185126));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__16_ (.o(regtop_dchdi_w1_hdi00[16]),
	.ck(clk),
	.d(n185125));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__17_ (.o(regtop_dchdi_w1_hdi00[17]),
	.ck(clk),
	.d(n185124));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__18_ (.o(regtop_dchdi_w1_hdi00[18]),
	.ck(clk),
	.d(n185123));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__19_ (.o(regtop_dchdi_w1_hdi00[19]),
	.ck(clk),
	.d(n185122));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__20_ (.o(regtop_dchdi_w1_hdi00[20]),
	.ck(clk),
	.d(n185121));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__21_ (.o(regtop_dchdi_w1_hdi00[21]),
	.ck(clk),
	.d(n185120));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__22_ (.o(regtop_dchdi_w1_hdi00[22]),
	.ck(clk),
	.d(n185119));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__23_ (.o(regtop_dchdi_w1_hdi00[23]),
	.ck(clk),
	.d(n185118));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__24_ (.o(regtop_dchdi_w1_hdi00[24]),
	.ck(clk),
	.d(n185117));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__25_ (.o(regtop_dchdi_w1_hdi00[25]),
	.ck(clk),
	.d(n185116));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__26_ (.o(regtop_dchdi_w1_hdi00[26]),
	.ck(clk),
	.d(n185115));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__27_ (.o(regtop_dchdi_w1_hdi00[27]),
	.ck(clk),
	.d(n185114));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__28_ (.o(regtop_dchdi_w1_hdi00[28]),
	.ck(clk),
	.d(n185113));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__29_ (.o(regtop_dchdi_w1_hdi00[29]),
	.ck(clk),
	.d(n185112));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__30_ (.o(regtop_dchdi_w1_hdi00[30]),
	.ck(clk),
	.d(n185111));
   ms00f80 regtop_dchdi_w1_hdi00_reg_48__31_ (.o(regtop_dchdi_w1_hdi00[31]),
	.ck(clk),
	.d(n185110));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__0_ (.o(regtop_dchdi_w1_hdi00[32]),
	.ck(clk),
	.d(n185109));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__1_ (.o(regtop_dchdi_w1_hdi00[33]),
	.ck(clk),
	.d(n185108));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__2_ (.o(regtop_dchdi_w1_hdi00[34]),
	.ck(clk),
	.d(n185107));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__3_ (.o(regtop_dchdi_w1_hdi00[35]),
	.ck(clk),
	.d(n185106));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__4_ (.o(regtop_dchdi_w1_hdi00[36]),
	.ck(clk),
	.d(n185105));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__5_ (.o(regtop_dchdi_w1_hdi00[37]),
	.ck(clk),
	.d(n185104));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__6_ (.o(regtop_dchdi_w1_hdi00[38]),
	.ck(clk),
	.d(n185103));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__7_ (.o(regtop_dchdi_w1_hdi00[39]),
	.ck(clk),
	.d(n185102));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__8_ (.o(regtop_dchdi_w1_hdi00[40]),
	.ck(clk),
	.d(n185101));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__9_ (.o(regtop_dchdi_w1_hdi00[41]),
	.ck(clk),
	.d(n185100));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__10_ (.o(regtop_dchdi_w1_hdi00[42]),
	.ck(clk),
	.d(n185099));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__11_ (.o(regtop_dchdi_w1_hdi00[43]),
	.ck(clk),
	.d(n185098));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__12_ (.o(regtop_dchdi_w1_hdi00[44]),
	.ck(clk),
	.d(n185097));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__13_ (.o(regtop_dchdi_w1_hdi00[45]),
	.ck(clk),
	.d(n185096));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__14_ (.o(regtop_dchdi_w1_hdi00[46]),
	.ck(clk),
	.d(n185095));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__15_ (.o(regtop_dchdi_w1_hdi00[47]),
	.ck(clk),
	.d(n185094));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__16_ (.o(regtop_dchdi_w1_hdi00[48]),
	.ck(clk),
	.d(n185093));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__17_ (.o(regtop_dchdi_w1_hdi00[49]),
	.ck(clk),
	.d(n185092));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__18_ (.o(regtop_dchdi_w1_hdi00[50]),
	.ck(clk),
	.d(n185091));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__19_ (.o(regtop_dchdi_w1_hdi00[51]),
	.ck(clk),
	.d(n185090));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__20_ (.o(regtop_dchdi_w1_hdi00[52]),
	.ck(clk),
	.d(n185089));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__21_ (.o(regtop_dchdi_w1_hdi00[53]),
	.ck(clk),
	.d(n185088));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__22_ (.o(regtop_dchdi_w1_hdi00[54]),
	.ck(clk),
	.d(n185087));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__23_ (.o(regtop_dchdi_w1_hdi00[55]),
	.ck(clk),
	.d(n185086));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__24_ (.o(regtop_dchdi_w1_hdi00[56]),
	.ck(clk),
	.d(n185085));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__25_ (.o(regtop_dchdi_w1_hdi00[57]),
	.ck(clk),
	.d(n185084));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__26_ (.o(regtop_dchdi_w1_hdi00[58]),
	.ck(clk),
	.d(n185083));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__27_ (.o(regtop_dchdi_w1_hdi00[59]),
	.ck(clk),
	.d(n185082));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__28_ (.o(regtop_dchdi_w1_hdi00[60]),
	.ck(clk),
	.d(n185081));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__29_ (.o(regtop_dchdi_w1_hdi00[61]),
	.ck(clk),
	.d(n185080));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__30_ (.o(regtop_dchdi_w1_hdi00[62]),
	.ck(clk),
	.d(n185079));
   ms00f80 regtop_dchdi_w1_hdi00_reg_49__31_ (.o(regtop_dchdi_w1_hdi00[63]),
	.ck(clk),
	.d(n185078));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__0_ (.o(regtop_dchdi_w1_hdi00[64]),
	.ck(clk),
	.d(n185077));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__1_ (.o(regtop_dchdi_w1_hdi00[65]),
	.ck(clk),
	.d(n185076));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__2_ (.o(regtop_dchdi_w1_hdi00[66]),
	.ck(clk),
	.d(n185075));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__3_ (.o(regtop_dchdi_w1_hdi00[67]),
	.ck(clk),
	.d(n185074));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__4_ (.o(regtop_dchdi_w1_hdi00[68]),
	.ck(clk),
	.d(n185073));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__5_ (.o(regtop_dchdi_w1_hdi00[69]),
	.ck(clk),
	.d(n185072));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__6_ (.o(regtop_dchdi_w1_hdi00[70]),
	.ck(clk),
	.d(n185071));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__7_ (.o(regtop_dchdi_w1_hdi00[71]),
	.ck(clk),
	.d(n185070));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__8_ (.o(regtop_dchdi_w1_hdi00[72]),
	.ck(clk),
	.d(n185069));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__9_ (.o(regtop_dchdi_w1_hdi00[73]),
	.ck(clk),
	.d(n185068));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__10_ (.o(regtop_dchdi_w1_hdi00[74]),
	.ck(clk),
	.d(n185067));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__11_ (.o(regtop_dchdi_w1_hdi00[75]),
	.ck(clk),
	.d(n185066));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__12_ (.o(regtop_dchdi_w1_hdi00[76]),
	.ck(clk),
	.d(n185065));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__13_ (.o(regtop_dchdi_w1_hdi00[77]),
	.ck(clk),
	.d(n185064));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__14_ (.o(regtop_dchdi_w1_hdi00[78]),
	.ck(clk),
	.d(n185063));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__15_ (.o(regtop_dchdi_w1_hdi00[79]),
	.ck(clk),
	.d(n185062));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__16_ (.o(regtop_dchdi_w1_hdi00[80]),
	.ck(clk),
	.d(n185061));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__17_ (.o(regtop_dchdi_w1_hdi00[81]),
	.ck(clk),
	.d(n185060));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__18_ (.o(regtop_dchdi_w1_hdi00[82]),
	.ck(clk),
	.d(n185059));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__19_ (.o(regtop_dchdi_w1_hdi00[83]),
	.ck(clk),
	.d(n185058));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__20_ (.o(regtop_dchdi_w1_hdi00[84]),
	.ck(clk),
	.d(n185057));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__21_ (.o(regtop_dchdi_w1_hdi00[85]),
	.ck(clk),
	.d(n185056));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__22_ (.o(regtop_dchdi_w1_hdi00[86]),
	.ck(clk),
	.d(n185055));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__23_ (.o(regtop_dchdi_w1_hdi00[87]),
	.ck(clk),
	.d(n185054));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__24_ (.o(regtop_dchdi_w1_hdi00[88]),
	.ck(clk),
	.d(n185053));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__25_ (.o(regtop_dchdi_w1_hdi00[89]),
	.ck(clk),
	.d(n185052));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__26_ (.o(regtop_dchdi_w1_hdi00[90]),
	.ck(clk),
	.d(n185051));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__27_ (.o(regtop_dchdi_w1_hdi00[91]),
	.ck(clk),
	.d(n185050));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__28_ (.o(regtop_dchdi_w1_hdi00[92]),
	.ck(clk),
	.d(n185049));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__29_ (.o(regtop_dchdi_w1_hdi00[93]),
	.ck(clk),
	.d(n185048));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__30_ (.o(regtop_dchdi_w1_hdi00[94]),
	.ck(clk),
	.d(n185047));
   ms00f80 regtop_dchdi_w1_hdi00_reg_50__31_ (.o(regtop_dchdi_w1_hdi00[95]),
	.ck(clk),
	.d(n185046));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__0_ (.o(regtop_dchdi_w1_hdi00[96]),
	.ck(clk),
	.d(n185045));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__1_ (.o(regtop_dchdi_w1_hdi00[97]),
	.ck(clk),
	.d(n185044));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__2_ (.o(regtop_dchdi_w1_hdi00[98]),
	.ck(clk),
	.d(n185043));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__3_ (.o(regtop_dchdi_w1_hdi00[99]),
	.ck(clk),
	.d(n185042));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__4_ (.o(regtop_dchdi_w1_hdi00[100]),
	.ck(clk),
	.d(n185041));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__5_ (.o(regtop_dchdi_w1_hdi00[101]),
	.ck(clk),
	.d(n185040));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__6_ (.o(regtop_dchdi_w1_hdi00[102]),
	.ck(clk),
	.d(n185039));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__7_ (.o(regtop_dchdi_w1_hdi00[103]),
	.ck(clk),
	.d(n185038));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__8_ (.o(regtop_dchdi_w1_hdi00[104]),
	.ck(clk),
	.d(n185037));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__9_ (.o(regtop_dchdi_w1_hdi00[105]),
	.ck(clk),
	.d(n185036));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__10_ (.o(regtop_dchdi_w1_hdi00[106]),
	.ck(clk),
	.d(n185035));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__11_ (.o(regtop_dchdi_w1_hdi00[107]),
	.ck(clk),
	.d(n185034));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__12_ (.o(regtop_dchdi_w1_hdi00[108]),
	.ck(clk),
	.d(n185033));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__13_ (.o(regtop_dchdi_w1_hdi00[109]),
	.ck(clk),
	.d(n185032));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__14_ (.o(regtop_dchdi_w1_hdi00[110]),
	.ck(clk),
	.d(n185031));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__15_ (.o(regtop_dchdi_w1_hdi00[111]),
	.ck(clk),
	.d(n185030));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__16_ (.o(regtop_dchdi_w1_hdi00[112]),
	.ck(clk),
	.d(n185029));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__17_ (.o(regtop_dchdi_w1_hdi00[113]),
	.ck(clk),
	.d(n185028));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__18_ (.o(regtop_dchdi_w1_hdi00[114]),
	.ck(clk),
	.d(n185027));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__19_ (.o(regtop_dchdi_w1_hdi00[115]),
	.ck(clk),
	.d(n185026));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__20_ (.o(regtop_dchdi_w1_hdi00[116]),
	.ck(clk),
	.d(n185025));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__21_ (.o(regtop_dchdi_w1_hdi00[117]),
	.ck(clk),
	.d(n185024));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__22_ (.o(regtop_dchdi_w1_hdi00[118]),
	.ck(clk),
	.d(n185023));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__23_ (.o(regtop_dchdi_w1_hdi00[119]),
	.ck(clk),
	.d(n185022));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__24_ (.o(regtop_dchdi_w1_hdi00[120]),
	.ck(clk),
	.d(n185021));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__25_ (.o(regtop_dchdi_w1_hdi00[121]),
	.ck(clk),
	.d(n185020));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__26_ (.o(regtop_dchdi_w1_hdi00[122]),
	.ck(clk),
	.d(n185019));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__27_ (.o(regtop_dchdi_w1_hdi00[123]),
	.ck(clk),
	.d(n185018));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__28_ (.o(regtop_dchdi_w1_hdi00[124]),
	.ck(clk),
	.d(n185017));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__29_ (.o(regtop_dchdi_w1_hdi00[125]),
	.ck(clk),
	.d(n185016));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__30_ (.o(regtop_dchdi_w1_hdi00[126]),
	.ck(clk),
	.d(n185015));
   ms00f80 regtop_dchdi_w1_hdi00_reg_51__31_ (.o(regtop_dchdi_w1_hdi00[127]),
	.ck(clk),
	.d(n185014));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__0_ (.o(regtop_dchdi_w1_hdi00[128]),
	.ck(clk),
	.d(n185013));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__1_ (.o(regtop_dchdi_w1_hdi00[129]),
	.ck(clk),
	.d(n185012));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__2_ (.o(regtop_dchdi_w1_hdi00[130]),
	.ck(clk),
	.d(n185011));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__3_ (.o(regtop_dchdi_w1_hdi00[131]),
	.ck(clk),
	.d(n185010));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__4_ (.o(regtop_dchdi_w1_hdi00[132]),
	.ck(clk),
	.d(n185009));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__5_ (.o(regtop_dchdi_w1_hdi00[133]),
	.ck(clk),
	.d(n185008));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__6_ (.o(regtop_dchdi_w1_hdi00[134]),
	.ck(clk),
	.d(n185007));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__7_ (.o(regtop_dchdi_w1_hdi00[135]),
	.ck(clk),
	.d(n185006));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__8_ (.o(regtop_dchdi_w1_hdi00[136]),
	.ck(clk),
	.d(n185005));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__9_ (.o(regtop_dchdi_w1_hdi00[137]),
	.ck(clk),
	.d(n185004));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__10_ (.o(regtop_dchdi_w1_hdi00[138]),
	.ck(clk),
	.d(n185003));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__11_ (.o(regtop_dchdi_w1_hdi00[139]),
	.ck(clk),
	.d(n185002));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__12_ (.o(regtop_dchdi_w1_hdi00[140]),
	.ck(clk),
	.d(n185001));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__13_ (.o(regtop_dchdi_w1_hdi00[141]),
	.ck(clk),
	.d(n185000));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__14_ (.o(regtop_dchdi_w1_hdi00[142]),
	.ck(clk),
	.d(n184999));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__15_ (.o(regtop_dchdi_w1_hdi00[143]),
	.ck(clk),
	.d(n184998));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__16_ (.o(regtop_dchdi_w1_hdi00[144]),
	.ck(clk),
	.d(n184997));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__17_ (.o(regtop_dchdi_w1_hdi00[145]),
	.ck(clk),
	.d(n184996));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__18_ (.o(regtop_dchdi_w1_hdi00[146]),
	.ck(clk),
	.d(n184995));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__19_ (.o(regtop_dchdi_w1_hdi00[147]),
	.ck(clk),
	.d(n184994));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__20_ (.o(regtop_dchdi_w1_hdi00[148]),
	.ck(clk),
	.d(n184993));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__21_ (.o(regtop_dchdi_w1_hdi00[149]),
	.ck(clk),
	.d(n184992));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__22_ (.o(regtop_dchdi_w1_hdi00[150]),
	.ck(clk),
	.d(n184991));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__23_ (.o(regtop_dchdi_w1_hdi00[151]),
	.ck(clk),
	.d(n184990));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__24_ (.o(regtop_dchdi_w1_hdi00[152]),
	.ck(clk),
	.d(n184989));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__25_ (.o(regtop_dchdi_w1_hdi00[153]),
	.ck(clk),
	.d(n184988));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__26_ (.o(regtop_dchdi_w1_hdi00[154]),
	.ck(clk),
	.d(n184987));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__27_ (.o(regtop_dchdi_w1_hdi00[155]),
	.ck(clk),
	.d(n184986));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__28_ (.o(regtop_dchdi_w1_hdi00[156]),
	.ck(clk),
	.d(n184985));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__29_ (.o(regtop_dchdi_w1_hdi00[157]),
	.ck(clk),
	.d(n184984));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__30_ (.o(regtop_dchdi_w1_hdi00[158]),
	.ck(clk),
	.d(n184983));
   ms00f80 regtop_dchdi_w1_hdi00_reg_52__31_ (.o(regtop_dchdi_w1_hdi00[159]),
	.ck(clk),
	.d(n184982));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__0_ (.o(regtop_dchdi_w1_hdi00[160]),
	.ck(clk),
	.d(n184981));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__1_ (.o(regtop_dchdi_w1_hdi00[161]),
	.ck(clk),
	.d(n184980));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__2_ (.o(regtop_dchdi_w1_hdi00[162]),
	.ck(clk),
	.d(n184979));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__3_ (.o(regtop_dchdi_w1_hdi00[163]),
	.ck(clk),
	.d(n184978));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__4_ (.o(regtop_dchdi_w1_hdi00[164]),
	.ck(clk),
	.d(n184977));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__5_ (.o(regtop_dchdi_w1_hdi00[165]),
	.ck(clk),
	.d(n184976));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__6_ (.o(regtop_dchdi_w1_hdi00[166]),
	.ck(clk),
	.d(n184975));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__7_ (.o(regtop_dchdi_w1_hdi00[167]),
	.ck(clk),
	.d(n184974));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__8_ (.o(regtop_dchdi_w1_hdi00[168]),
	.ck(clk),
	.d(n184973));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__9_ (.o(regtop_dchdi_w1_hdi00[169]),
	.ck(clk),
	.d(n184972));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__10_ (.o(regtop_dchdi_w1_hdi00[170]),
	.ck(clk),
	.d(n184971));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__11_ (.o(regtop_dchdi_w1_hdi00[171]),
	.ck(clk),
	.d(n184970));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__12_ (.o(regtop_dchdi_w1_hdi00[172]),
	.ck(clk),
	.d(n184969));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__13_ (.o(regtop_dchdi_w1_hdi00[173]),
	.ck(clk),
	.d(n184968));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__14_ (.o(regtop_dchdi_w1_hdi00[174]),
	.ck(clk),
	.d(n184967));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__15_ (.o(regtop_dchdi_w1_hdi00[175]),
	.ck(clk),
	.d(n184966));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__16_ (.o(regtop_dchdi_w1_hdi00[176]),
	.ck(clk),
	.d(n184965));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__17_ (.o(regtop_dchdi_w1_hdi00[177]),
	.ck(clk),
	.d(n184964));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__18_ (.o(regtop_dchdi_w1_hdi00[178]),
	.ck(clk),
	.d(n184963));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__19_ (.o(regtop_dchdi_w1_hdi00[179]),
	.ck(clk),
	.d(n184962));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__20_ (.o(regtop_dchdi_w1_hdi00[180]),
	.ck(clk),
	.d(n184961));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__21_ (.o(regtop_dchdi_w1_hdi00[181]),
	.ck(clk),
	.d(n184960));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__22_ (.o(regtop_dchdi_w1_hdi00[182]),
	.ck(clk),
	.d(n184959));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__23_ (.o(regtop_dchdi_w1_hdi00[183]),
	.ck(clk),
	.d(n184958));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__24_ (.o(regtop_dchdi_w1_hdi00[184]),
	.ck(clk),
	.d(n184957));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__25_ (.o(regtop_dchdi_w1_hdi00[185]),
	.ck(clk),
	.d(n184956));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__26_ (.o(regtop_dchdi_w1_hdi00[186]),
	.ck(clk),
	.d(n184955));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__27_ (.o(regtop_dchdi_w1_hdi00[187]),
	.ck(clk),
	.d(n184954));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__28_ (.o(regtop_dchdi_w1_hdi00[188]),
	.ck(clk),
	.d(n184953));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__29_ (.o(regtop_dchdi_w1_hdi00[189]),
	.ck(clk),
	.d(n184952));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__30_ (.o(regtop_dchdi_w1_hdi00[190]),
	.ck(clk),
	.d(n184951));
   ms00f80 regtop_dchdi_w1_hdi00_reg_53__31_ (.o(regtop_dchdi_w1_hdi00[191]),
	.ck(clk),
	.d(n184950));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__0_ (.o(regtop_dchdi_w1_hdi00[192]),
	.ck(clk),
	.d(n184949));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__1_ (.o(regtop_dchdi_w1_hdi00[193]),
	.ck(clk),
	.d(n184948));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__2_ (.o(regtop_dchdi_w1_hdi00[194]),
	.ck(clk),
	.d(n184947));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__3_ (.o(regtop_dchdi_w1_hdi00[195]),
	.ck(clk),
	.d(n184946));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__4_ (.o(regtop_dchdi_w1_hdi00[196]),
	.ck(clk),
	.d(n184945));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__5_ (.o(regtop_dchdi_w1_hdi00[197]),
	.ck(clk),
	.d(n184944));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__6_ (.o(regtop_dchdi_w1_hdi00[198]),
	.ck(clk),
	.d(n184943));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__7_ (.o(regtop_dchdi_w1_hdi00[199]),
	.ck(clk),
	.d(n184942));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__8_ (.o(regtop_dchdi_w1_hdi00[200]),
	.ck(clk),
	.d(n184941));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__9_ (.o(regtop_dchdi_w1_hdi00[201]),
	.ck(clk),
	.d(n184940));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__10_ (.o(regtop_dchdi_w1_hdi00[202]),
	.ck(clk),
	.d(n184939));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__11_ (.o(regtop_dchdi_w1_hdi00[203]),
	.ck(clk),
	.d(n184938));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__12_ (.o(regtop_dchdi_w1_hdi00[204]),
	.ck(clk),
	.d(n184937));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__13_ (.o(regtop_dchdi_w1_hdi00[205]),
	.ck(clk),
	.d(n184936));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__14_ (.o(regtop_dchdi_w1_hdi00[206]),
	.ck(clk),
	.d(n184935));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__15_ (.o(regtop_dchdi_w1_hdi00[207]),
	.ck(clk),
	.d(n184934));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__16_ (.o(regtop_dchdi_w1_hdi00[208]),
	.ck(clk),
	.d(n184933));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__17_ (.o(regtop_dchdi_w1_hdi00[209]),
	.ck(clk),
	.d(n184932));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__18_ (.o(regtop_dchdi_w1_hdi00[210]),
	.ck(clk),
	.d(n184931));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__19_ (.o(regtop_dchdi_w1_hdi00[211]),
	.ck(clk),
	.d(n184930));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__20_ (.o(regtop_dchdi_w1_hdi00[212]),
	.ck(clk),
	.d(n184929));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__21_ (.o(regtop_dchdi_w1_hdi00[213]),
	.ck(clk),
	.d(n184928));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__22_ (.o(regtop_dchdi_w1_hdi00[214]),
	.ck(clk),
	.d(n184927));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__23_ (.o(regtop_dchdi_w1_hdi00[215]),
	.ck(clk),
	.d(n184926));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__24_ (.o(regtop_dchdi_w1_hdi00[216]),
	.ck(clk),
	.d(n184925));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__25_ (.o(regtop_dchdi_w1_hdi00[217]),
	.ck(clk),
	.d(n184924));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__26_ (.o(regtop_dchdi_w1_hdi00[218]),
	.ck(clk),
	.d(n184923));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__27_ (.o(regtop_dchdi_w1_hdi00[219]),
	.ck(clk),
	.d(n184922));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__28_ (.o(regtop_dchdi_w1_hdi00[220]),
	.ck(clk),
	.d(n184921));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__29_ (.o(regtop_dchdi_w1_hdi00[221]),
	.ck(clk),
	.d(n184920));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__30_ (.o(regtop_dchdi_w1_hdi00[222]),
	.ck(clk),
	.d(n184919));
   ms00f80 regtop_dchdi_w1_hdi00_reg_54__31_ (.o(regtop_dchdi_w1_hdi00[223]),
	.ck(clk),
	.d(n184918));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__0_ (.o(regtop_dchdi_w1_hdi00[224]),
	.ck(clk),
	.d(n184917));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__1_ (.o(regtop_dchdi_w1_hdi00[225]),
	.ck(clk),
	.d(n184916));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__2_ (.o(regtop_dchdi_w1_hdi00[226]),
	.ck(clk),
	.d(n184915));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__3_ (.o(regtop_dchdi_w1_hdi00[227]),
	.ck(clk),
	.d(n184914));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__4_ (.o(regtop_dchdi_w1_hdi00[228]),
	.ck(clk),
	.d(n184913));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__5_ (.o(regtop_dchdi_w1_hdi00[229]),
	.ck(clk),
	.d(n184912));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__6_ (.o(regtop_dchdi_w1_hdi00[230]),
	.ck(clk),
	.d(n184911));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__7_ (.o(regtop_dchdi_w1_hdi00[231]),
	.ck(clk),
	.d(n184910));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__8_ (.o(regtop_dchdi_w1_hdi00[232]),
	.ck(clk),
	.d(n184909));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__9_ (.o(regtop_dchdi_w1_hdi00[233]),
	.ck(clk),
	.d(n184908));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__10_ (.o(regtop_dchdi_w1_hdi00[234]),
	.ck(clk),
	.d(n184907));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__11_ (.o(regtop_dchdi_w1_hdi00[235]),
	.ck(clk),
	.d(n184906));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__12_ (.o(regtop_dchdi_w1_hdi00[236]),
	.ck(clk),
	.d(n184905));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__13_ (.o(regtop_dchdi_w1_hdi00[237]),
	.ck(clk),
	.d(n184904));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__14_ (.o(regtop_dchdi_w1_hdi00[238]),
	.ck(clk),
	.d(n184903));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__15_ (.o(regtop_dchdi_w1_hdi00[239]),
	.ck(clk),
	.d(n184902));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__16_ (.o(regtop_dchdi_w1_hdi00[240]),
	.ck(clk),
	.d(n184901));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__17_ (.o(regtop_dchdi_w1_hdi00[241]),
	.ck(clk),
	.d(n184900));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__18_ (.o(regtop_dchdi_w1_hdi00[242]),
	.ck(clk),
	.d(n184899));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__19_ (.o(regtop_dchdi_w1_hdi00[243]),
	.ck(clk),
	.d(n184898));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__20_ (.o(regtop_dchdi_w1_hdi00[244]),
	.ck(clk),
	.d(n184897));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__21_ (.o(regtop_dchdi_w1_hdi00[245]),
	.ck(clk),
	.d(n184896));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__22_ (.o(regtop_dchdi_w1_hdi00[246]),
	.ck(clk),
	.d(n184895));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__23_ (.o(regtop_dchdi_w1_hdi00[247]),
	.ck(clk),
	.d(n184894));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__24_ (.o(regtop_dchdi_w1_hdi00[248]),
	.ck(clk),
	.d(n184893));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__25_ (.o(regtop_dchdi_w1_hdi00[249]),
	.ck(clk),
	.d(n184892));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__26_ (.o(regtop_dchdi_w1_hdi00[250]),
	.ck(clk),
	.d(n184891));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__27_ (.o(regtop_dchdi_w1_hdi00[251]),
	.ck(clk),
	.d(n184890));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__28_ (.o(regtop_dchdi_w1_hdi00[252]),
	.ck(clk),
	.d(n184889));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__29_ (.o(regtop_dchdi_w1_hdi00[253]),
	.ck(clk),
	.d(n184888));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__30_ (.o(regtop_dchdi_w1_hdi00[254]),
	.ck(clk),
	.d(n184887));
   ms00f80 regtop_dchdi_w1_hdi00_reg_55__31_ (.o(regtop_dchdi_w1_hdi00[255]),
	.ck(clk),
	.d(n184886));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__0_ (.o(regtop_dchdi_w1_hdi00[256]),
	.ck(clk),
	.d(n184885));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__1_ (.o(regtop_dchdi_w1_hdi00[257]),
	.ck(clk),
	.d(n184884));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__2_ (.o(regtop_dchdi_w1_hdi00[258]),
	.ck(clk),
	.d(n184883));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__3_ (.o(regtop_dchdi_w1_hdi00[259]),
	.ck(clk),
	.d(n184882));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__4_ (.o(regtop_dchdi_w1_hdi00[260]),
	.ck(clk),
	.d(n184881));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__5_ (.o(regtop_dchdi_w1_hdi00[261]),
	.ck(clk),
	.d(n184880));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__6_ (.o(regtop_dchdi_w1_hdi00[262]),
	.ck(clk),
	.d(n184879));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__7_ (.o(regtop_dchdi_w1_hdi00[263]),
	.ck(clk),
	.d(n184878));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__8_ (.o(regtop_dchdi_w1_hdi00[264]),
	.ck(clk),
	.d(n184877));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__9_ (.o(regtop_dchdi_w1_hdi00[265]),
	.ck(clk),
	.d(n184876));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__10_ (.o(regtop_dchdi_w1_hdi00[266]),
	.ck(clk),
	.d(n184875));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__11_ (.o(regtop_dchdi_w1_hdi00[267]),
	.ck(clk),
	.d(n184874));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__12_ (.o(regtop_dchdi_w1_hdi00[268]),
	.ck(clk),
	.d(n184873));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__13_ (.o(regtop_dchdi_w1_hdi00[269]),
	.ck(clk),
	.d(n184872));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__14_ (.o(regtop_dchdi_w1_hdi00[270]),
	.ck(clk),
	.d(n184871));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__15_ (.o(regtop_dchdi_w1_hdi00[271]),
	.ck(clk),
	.d(n184870));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__16_ (.o(regtop_dchdi_w1_hdi00[272]),
	.ck(clk),
	.d(n184869));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__17_ (.o(regtop_dchdi_w1_hdi00[273]),
	.ck(clk),
	.d(n184868));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__18_ (.o(regtop_dchdi_w1_hdi00[274]),
	.ck(clk),
	.d(n184867));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__19_ (.o(regtop_dchdi_w1_hdi00[275]),
	.ck(clk),
	.d(n184866));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__20_ (.o(regtop_dchdi_w1_hdi00[276]),
	.ck(clk),
	.d(n184865));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__21_ (.o(regtop_dchdi_w1_hdi00[277]),
	.ck(clk),
	.d(n184864));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__22_ (.o(regtop_dchdi_w1_hdi00[278]),
	.ck(clk),
	.d(n184863));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__23_ (.o(regtop_dchdi_w1_hdi00[279]),
	.ck(clk),
	.d(n184862));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__24_ (.o(regtop_dchdi_w1_hdi00[280]),
	.ck(clk),
	.d(n184861));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__25_ (.o(regtop_dchdi_w1_hdi00[281]),
	.ck(clk),
	.d(n184860));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__26_ (.o(regtop_dchdi_w1_hdi00[282]),
	.ck(clk),
	.d(n184859));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__27_ (.o(regtop_dchdi_w1_hdi00[283]),
	.ck(clk),
	.d(n184858));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__28_ (.o(regtop_dchdi_w1_hdi00[284]),
	.ck(clk),
	.d(n184857));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__29_ (.o(regtop_dchdi_w1_hdi00[285]),
	.ck(clk),
	.d(n184856));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__30_ (.o(regtop_dchdi_w1_hdi00[286]),
	.ck(clk),
	.d(n184855));
   ms00f80 regtop_dchdi_w1_hdi00_reg_56__31_ (.o(regtop_dchdi_w1_hdi00[287]),
	.ck(clk),
	.d(n184854));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__0_ (.o(regtop_dchdi_w1_hdi00[288]),
	.ck(clk),
	.d(n184853));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__1_ (.o(regtop_dchdi_w1_hdi00[289]),
	.ck(clk),
	.d(n184852));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__2_ (.o(regtop_dchdi_w1_hdi00[290]),
	.ck(clk),
	.d(n184851));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__3_ (.o(regtop_dchdi_w1_hdi00[291]),
	.ck(clk),
	.d(n184850));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__4_ (.o(regtop_dchdi_w1_hdi00[292]),
	.ck(clk),
	.d(n184849));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__5_ (.o(regtop_dchdi_w1_hdi00[293]),
	.ck(clk),
	.d(n184848));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__6_ (.o(regtop_dchdi_w1_hdi00[294]),
	.ck(clk),
	.d(n184847));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__7_ (.o(regtop_dchdi_w1_hdi00[295]),
	.ck(clk),
	.d(n184846));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__8_ (.o(regtop_dchdi_w1_hdi00[296]),
	.ck(clk),
	.d(n184845));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__9_ (.o(regtop_dchdi_w1_hdi00[297]),
	.ck(clk),
	.d(n184844));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__10_ (.o(regtop_dchdi_w1_hdi00[298]),
	.ck(clk),
	.d(n184843));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__11_ (.o(regtop_dchdi_w1_hdi00[299]),
	.ck(clk),
	.d(n184842));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__12_ (.o(regtop_dchdi_w1_hdi00[300]),
	.ck(clk),
	.d(n184841));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__13_ (.o(regtop_dchdi_w1_hdi00[301]),
	.ck(clk),
	.d(n184840));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__14_ (.o(regtop_dchdi_w1_hdi00[302]),
	.ck(clk),
	.d(n184839));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__15_ (.o(regtop_dchdi_w1_hdi00[303]),
	.ck(clk),
	.d(n184838));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__16_ (.o(regtop_dchdi_w1_hdi00[304]),
	.ck(clk),
	.d(n184837));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__17_ (.o(regtop_dchdi_w1_hdi00[305]),
	.ck(clk),
	.d(n184836));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__18_ (.o(regtop_dchdi_w1_hdi00[306]),
	.ck(clk),
	.d(n184835));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__19_ (.o(regtop_dchdi_w1_hdi00[307]),
	.ck(clk),
	.d(n184834));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__20_ (.o(regtop_dchdi_w1_hdi00[308]),
	.ck(clk),
	.d(n184833));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__21_ (.o(regtop_dchdi_w1_hdi00[309]),
	.ck(clk),
	.d(n184832));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__22_ (.o(regtop_dchdi_w1_hdi00[310]),
	.ck(clk),
	.d(n184831));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__23_ (.o(regtop_dchdi_w1_hdi00[311]),
	.ck(clk),
	.d(n184830));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__24_ (.o(regtop_dchdi_w1_hdi00[312]),
	.ck(clk),
	.d(n184829));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__25_ (.o(regtop_dchdi_w1_hdi00[313]),
	.ck(clk),
	.d(n184828));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__26_ (.o(regtop_dchdi_w1_hdi00[314]),
	.ck(clk),
	.d(n184827));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__27_ (.o(regtop_dchdi_w1_hdi00[315]),
	.ck(clk),
	.d(n184826));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__28_ (.o(regtop_dchdi_w1_hdi00[316]),
	.ck(clk),
	.d(n184825));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__29_ (.o(regtop_dchdi_w1_hdi00[317]),
	.ck(clk),
	.d(n184824));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__30_ (.o(regtop_dchdi_w1_hdi00[318]),
	.ck(clk),
	.d(n184823));
   ms00f80 regtop_dchdi_w1_hdi00_reg_57__31_ (.o(regtop_dchdi_w1_hdi00[319]),
	.ck(clk),
	.d(n184822));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__0_ (.o(regtop_dchdi_w1_hdi00[320]),
	.ck(clk),
	.d(n184821));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__1_ (.o(regtop_dchdi_w1_hdi00[321]),
	.ck(clk),
	.d(n184820));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__2_ (.o(regtop_dchdi_w1_hdi00[322]),
	.ck(clk),
	.d(n184819));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__3_ (.o(regtop_dchdi_w1_hdi00[323]),
	.ck(clk),
	.d(n184818));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__4_ (.o(regtop_dchdi_w1_hdi00[324]),
	.ck(clk),
	.d(n184817));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__5_ (.o(regtop_dchdi_w1_hdi00[325]),
	.ck(clk),
	.d(n184816));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__6_ (.o(regtop_dchdi_w1_hdi00[326]),
	.ck(clk),
	.d(n184815));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__7_ (.o(regtop_dchdi_w1_hdi00[327]),
	.ck(clk),
	.d(n184814));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__8_ (.o(regtop_dchdi_w1_hdi00[328]),
	.ck(clk),
	.d(n184813));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__9_ (.o(regtop_dchdi_w1_hdi00[329]),
	.ck(clk),
	.d(n184812));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__10_ (.o(regtop_dchdi_w1_hdi00[330]),
	.ck(clk),
	.d(n184811));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__11_ (.o(regtop_dchdi_w1_hdi00[331]),
	.ck(clk),
	.d(n184810));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__12_ (.o(regtop_dchdi_w1_hdi00[332]),
	.ck(clk),
	.d(n184809));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__13_ (.o(regtop_dchdi_w1_hdi00[333]),
	.ck(clk),
	.d(n184808));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__14_ (.o(regtop_dchdi_w1_hdi00[334]),
	.ck(clk),
	.d(n184807));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__15_ (.o(regtop_dchdi_w1_hdi00[335]),
	.ck(clk),
	.d(n184806));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__16_ (.o(regtop_dchdi_w1_hdi00[336]),
	.ck(clk),
	.d(n184805));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__17_ (.o(regtop_dchdi_w1_hdi00[337]),
	.ck(clk),
	.d(n184804));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__18_ (.o(regtop_dchdi_w1_hdi00[338]),
	.ck(clk),
	.d(n184803));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__19_ (.o(regtop_dchdi_w1_hdi00[339]),
	.ck(clk),
	.d(n184802));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__20_ (.o(regtop_dchdi_w1_hdi00[340]),
	.ck(clk),
	.d(n184801));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__21_ (.o(regtop_dchdi_w1_hdi00[341]),
	.ck(clk),
	.d(n184800));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__22_ (.o(regtop_dchdi_w1_hdi00[342]),
	.ck(clk),
	.d(n184799));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__23_ (.o(regtop_dchdi_w1_hdi00[343]),
	.ck(clk),
	.d(n184798));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__24_ (.o(regtop_dchdi_w1_hdi00[344]),
	.ck(clk),
	.d(n184797));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__25_ (.o(regtop_dchdi_w1_hdi00[345]),
	.ck(clk),
	.d(n184796));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__26_ (.o(regtop_dchdi_w1_hdi00[346]),
	.ck(clk),
	.d(n184795));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__27_ (.o(regtop_dchdi_w1_hdi00[347]),
	.ck(clk),
	.d(n184794));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__28_ (.o(regtop_dchdi_w1_hdi00[348]),
	.ck(clk),
	.d(n184793));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__29_ (.o(regtop_dchdi_w1_hdi00[349]),
	.ck(clk),
	.d(n184792));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__30_ (.o(regtop_dchdi_w1_hdi00[350]),
	.ck(clk),
	.d(n184791));
   ms00f80 regtop_dchdi_w1_hdi00_reg_58__31_ (.o(regtop_dchdi_w1_hdi00[351]),
	.ck(clk),
	.d(n184790));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__0_ (.o(regtop_dchdi_w1_hdi00[352]),
	.ck(clk),
	.d(n184789));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__1_ (.o(regtop_dchdi_w1_hdi00[353]),
	.ck(clk),
	.d(n184788));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__2_ (.o(regtop_dchdi_w1_hdi00[354]),
	.ck(clk),
	.d(n184787));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__3_ (.o(regtop_dchdi_w1_hdi00[355]),
	.ck(clk),
	.d(n184786));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__4_ (.o(regtop_dchdi_w1_hdi00[356]),
	.ck(clk),
	.d(n184785));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__5_ (.o(regtop_dchdi_w1_hdi00[357]),
	.ck(clk),
	.d(n184784));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__6_ (.o(regtop_dchdi_w1_hdi00[358]),
	.ck(clk),
	.d(n184783));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__7_ (.o(regtop_dchdi_w1_hdi00[359]),
	.ck(clk),
	.d(n184782));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__8_ (.o(regtop_dchdi_w1_hdi00[360]),
	.ck(clk),
	.d(n184781));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__9_ (.o(regtop_dchdi_w1_hdi00[361]),
	.ck(clk),
	.d(n184780));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__10_ (.o(regtop_dchdi_w1_hdi00[362]),
	.ck(clk),
	.d(n184779));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__11_ (.o(regtop_dchdi_w1_hdi00[363]),
	.ck(clk),
	.d(n184778));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__12_ (.o(regtop_dchdi_w1_hdi00[364]),
	.ck(clk),
	.d(n184777));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__13_ (.o(regtop_dchdi_w1_hdi00[365]),
	.ck(clk),
	.d(n184776));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__14_ (.o(regtop_dchdi_w1_hdi00[366]),
	.ck(clk),
	.d(n184775));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__15_ (.o(regtop_dchdi_w1_hdi00[367]),
	.ck(clk),
	.d(n184774));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__16_ (.o(regtop_dchdi_w1_hdi00[368]),
	.ck(clk),
	.d(n184773));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__17_ (.o(regtop_dchdi_w1_hdi00[369]),
	.ck(clk),
	.d(n184772));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__18_ (.o(regtop_dchdi_w1_hdi00[370]),
	.ck(clk),
	.d(n184771));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__19_ (.o(regtop_dchdi_w1_hdi00[371]),
	.ck(clk),
	.d(n184770));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__20_ (.o(regtop_dchdi_w1_hdi00[372]),
	.ck(clk),
	.d(n184769));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__21_ (.o(regtop_dchdi_w1_hdi00[373]),
	.ck(clk),
	.d(n184768));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__22_ (.o(regtop_dchdi_w1_hdi00[374]),
	.ck(clk),
	.d(n184767));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__23_ (.o(regtop_dchdi_w1_hdi00[375]),
	.ck(clk),
	.d(n184766));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__24_ (.o(regtop_dchdi_w1_hdi00[376]),
	.ck(clk),
	.d(n184765));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__25_ (.o(regtop_dchdi_w1_hdi00[377]),
	.ck(clk),
	.d(n184764));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__26_ (.o(regtop_dchdi_w1_hdi00[378]),
	.ck(clk),
	.d(n184763));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__27_ (.o(regtop_dchdi_w1_hdi00[379]),
	.ck(clk),
	.d(n184762));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__28_ (.o(regtop_dchdi_w1_hdi00[380]),
	.ck(clk),
	.d(n184761));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__29_ (.o(regtop_dchdi_w1_hdi00[381]),
	.ck(clk),
	.d(n184760));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__30_ (.o(regtop_dchdi_w1_hdi00[382]),
	.ck(clk),
	.d(n184759));
   ms00f80 regtop_dchdi_w1_hdi00_reg_59__31_ (.o(regtop_dchdi_w1_hdi00[383]),
	.ck(clk),
	.d(n184758));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__0_ (.o(regtop_dchdi_w1_hdi00[384]),
	.ck(clk),
	.d(n184757));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__1_ (.o(regtop_dchdi_w1_hdi00[385]),
	.ck(clk),
	.d(n184756));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__2_ (.o(regtop_dchdi_w1_hdi00[386]),
	.ck(clk),
	.d(n184755));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__3_ (.o(regtop_dchdi_w1_hdi00[387]),
	.ck(clk),
	.d(n184754));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__4_ (.o(regtop_dchdi_w1_hdi00[388]),
	.ck(clk),
	.d(n184753));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__5_ (.o(regtop_dchdi_w1_hdi00[389]),
	.ck(clk),
	.d(n184752));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__6_ (.o(regtop_dchdi_w1_hdi00[390]),
	.ck(clk),
	.d(n184751));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__7_ (.o(regtop_dchdi_w1_hdi00[391]),
	.ck(clk),
	.d(n184750));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__8_ (.o(regtop_dchdi_w1_hdi00[392]),
	.ck(clk),
	.d(n184749));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__9_ (.o(regtop_dchdi_w1_hdi00[393]),
	.ck(clk),
	.d(n184748));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__10_ (.o(regtop_dchdi_w1_hdi00[394]),
	.ck(clk),
	.d(n184747));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__11_ (.o(regtop_dchdi_w1_hdi00[395]),
	.ck(clk),
	.d(n184746));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__12_ (.o(regtop_dchdi_w1_hdi00[396]),
	.ck(clk),
	.d(n184745));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__13_ (.o(regtop_dchdi_w1_hdi00[397]),
	.ck(clk),
	.d(n184744));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__14_ (.o(regtop_dchdi_w1_hdi00[398]),
	.ck(clk),
	.d(n184743));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__15_ (.o(regtop_dchdi_w1_hdi00[399]),
	.ck(clk),
	.d(n184742));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__16_ (.o(regtop_dchdi_w1_hdi00[400]),
	.ck(clk),
	.d(n184741));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__17_ (.o(regtop_dchdi_w1_hdi00[401]),
	.ck(clk),
	.d(n184740));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__18_ (.o(regtop_dchdi_w1_hdi00[402]),
	.ck(clk),
	.d(n184739));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__19_ (.o(regtop_dchdi_w1_hdi00[403]),
	.ck(clk),
	.d(n184738));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__20_ (.o(regtop_dchdi_w1_hdi00[404]),
	.ck(clk),
	.d(n184737));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__21_ (.o(regtop_dchdi_w1_hdi00[405]),
	.ck(clk),
	.d(n184736));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__22_ (.o(regtop_dchdi_w1_hdi00[406]),
	.ck(clk),
	.d(n184735));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__23_ (.o(regtop_dchdi_w1_hdi00[407]),
	.ck(clk),
	.d(n184734));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__24_ (.o(regtop_dchdi_w1_hdi00[408]),
	.ck(clk),
	.d(n184733));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__25_ (.o(regtop_dchdi_w1_hdi00[409]),
	.ck(clk),
	.d(n184732));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__26_ (.o(regtop_dchdi_w1_hdi00[410]),
	.ck(clk),
	.d(n184731));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__27_ (.o(regtop_dchdi_w1_hdi00[411]),
	.ck(clk),
	.d(n184730));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__28_ (.o(regtop_dchdi_w1_hdi00[412]),
	.ck(clk),
	.d(n184729));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__29_ (.o(regtop_dchdi_w1_hdi00[413]),
	.ck(clk),
	.d(n184728));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__30_ (.o(regtop_dchdi_w1_hdi00[414]),
	.ck(clk),
	.d(n184727));
   ms00f80 regtop_dchdi_w1_hdi00_reg_60__31_ (.o(regtop_dchdi_w1_hdi00[415]),
	.ck(clk),
	.d(n184726));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__0_ (.o(regtop_dchdi_w1_hdi00[416]),
	.ck(clk),
	.d(n184725));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__1_ (.o(regtop_dchdi_w1_hdi00[417]),
	.ck(clk),
	.d(n184724));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__2_ (.o(regtop_dchdi_w1_hdi00[418]),
	.ck(clk),
	.d(n184723));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__3_ (.o(regtop_dchdi_w1_hdi00[419]),
	.ck(clk),
	.d(n184722));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__4_ (.o(regtop_dchdi_w1_hdi00[420]),
	.ck(clk),
	.d(n184721));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__5_ (.o(regtop_dchdi_w1_hdi00[421]),
	.ck(clk),
	.d(n184720));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__6_ (.o(regtop_dchdi_w1_hdi00[422]),
	.ck(clk),
	.d(n184719));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__7_ (.o(regtop_dchdi_w1_hdi00[423]),
	.ck(clk),
	.d(n184718));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__8_ (.o(regtop_dchdi_w1_hdi00[424]),
	.ck(clk),
	.d(n184717));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__9_ (.o(regtop_dchdi_w1_hdi00[425]),
	.ck(clk),
	.d(n184716));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__10_ (.o(regtop_dchdi_w1_hdi00[426]),
	.ck(clk),
	.d(n184715));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__11_ (.o(regtop_dchdi_w1_hdi00[427]),
	.ck(clk),
	.d(n184714));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__12_ (.o(regtop_dchdi_w1_hdi00[428]),
	.ck(clk),
	.d(n184713));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__13_ (.o(regtop_dchdi_w1_hdi00[429]),
	.ck(clk),
	.d(n184712));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__14_ (.o(regtop_dchdi_w1_hdi00[430]),
	.ck(clk),
	.d(n184711));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__15_ (.o(regtop_dchdi_w1_hdi00[431]),
	.ck(clk),
	.d(n184710));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__16_ (.o(regtop_dchdi_w1_hdi00[432]),
	.ck(clk),
	.d(n184709));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__17_ (.o(regtop_dchdi_w1_hdi00[433]),
	.ck(clk),
	.d(n184708));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__18_ (.o(regtop_dchdi_w1_hdi00[434]),
	.ck(clk),
	.d(n184707));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__19_ (.o(regtop_dchdi_w1_hdi00[435]),
	.ck(clk),
	.d(n184706));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__20_ (.o(regtop_dchdi_w1_hdi00[436]),
	.ck(clk),
	.d(n184705));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__21_ (.o(regtop_dchdi_w1_hdi00[437]),
	.ck(clk),
	.d(n184704));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__22_ (.o(regtop_dchdi_w1_hdi00[438]),
	.ck(clk),
	.d(n184703));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__23_ (.o(regtop_dchdi_w1_hdi00[439]),
	.ck(clk),
	.d(n184702));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__24_ (.o(regtop_dchdi_w1_hdi00[440]),
	.ck(clk),
	.d(n184701));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__25_ (.o(regtop_dchdi_w1_hdi00[441]),
	.ck(clk),
	.d(n184700));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__26_ (.o(regtop_dchdi_w1_hdi00[442]),
	.ck(clk),
	.d(n184699));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__27_ (.o(regtop_dchdi_w1_hdi00[443]),
	.ck(clk),
	.d(n184698));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__28_ (.o(regtop_dchdi_w1_hdi00[444]),
	.ck(clk),
	.d(n184697));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__29_ (.o(regtop_dchdi_w1_hdi00[445]),
	.ck(clk),
	.d(n184696));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__30_ (.o(regtop_dchdi_w1_hdi00[446]),
	.ck(clk),
	.d(n184695));
   ms00f80 regtop_dchdi_w1_hdi00_reg_61__31_ (.o(regtop_dchdi_w1_hdi00[447]),
	.ck(clk),
	.d(n184694));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__0_ (.o(regtop_dchdi_w1_hdi00[448]),
	.ck(clk),
	.d(n184693));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__1_ (.o(regtop_dchdi_w1_hdi00[449]),
	.ck(clk),
	.d(n184692));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__2_ (.o(regtop_dchdi_w1_hdi00[450]),
	.ck(clk),
	.d(n184691));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__3_ (.o(regtop_dchdi_w1_hdi00[451]),
	.ck(clk),
	.d(n184690));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__4_ (.o(regtop_dchdi_w1_hdi00[452]),
	.ck(clk),
	.d(n184689));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__5_ (.o(regtop_dchdi_w1_hdi00[453]),
	.ck(clk),
	.d(n184688));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__6_ (.o(regtop_dchdi_w1_hdi00[454]),
	.ck(clk),
	.d(n184687));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__7_ (.o(regtop_dchdi_w1_hdi00[455]),
	.ck(clk),
	.d(n184686));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__8_ (.o(regtop_dchdi_w1_hdi00[456]),
	.ck(clk),
	.d(n184685));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__9_ (.o(regtop_dchdi_w1_hdi00[457]),
	.ck(clk),
	.d(n184684));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__10_ (.o(regtop_dchdi_w1_hdi00[458]),
	.ck(clk),
	.d(n184683));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__11_ (.o(regtop_dchdi_w1_hdi00[459]),
	.ck(clk),
	.d(n184682));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__12_ (.o(regtop_dchdi_w1_hdi00[460]),
	.ck(clk),
	.d(n184681));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__13_ (.o(regtop_dchdi_w1_hdi00[461]),
	.ck(clk),
	.d(n184680));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__14_ (.o(regtop_dchdi_w1_hdi00[462]),
	.ck(clk),
	.d(n184679));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__15_ (.o(regtop_dchdi_w1_hdi00[463]),
	.ck(clk),
	.d(n184678));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__16_ (.o(regtop_dchdi_w1_hdi00[464]),
	.ck(clk),
	.d(n184677));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__17_ (.o(regtop_dchdi_w1_hdi00[465]),
	.ck(clk),
	.d(n184676));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__18_ (.o(regtop_dchdi_w1_hdi00[466]),
	.ck(clk),
	.d(n184675));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__19_ (.o(regtop_dchdi_w1_hdi00[467]),
	.ck(clk),
	.d(n184674));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__20_ (.o(regtop_dchdi_w1_hdi00[468]),
	.ck(clk),
	.d(n184673));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__21_ (.o(regtop_dchdi_w1_hdi00[469]),
	.ck(clk),
	.d(n184672));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__22_ (.o(regtop_dchdi_w1_hdi00[470]),
	.ck(clk),
	.d(n184671));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__23_ (.o(regtop_dchdi_w1_hdi00[471]),
	.ck(clk),
	.d(n184670));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__24_ (.o(regtop_dchdi_w1_hdi00[472]),
	.ck(clk),
	.d(n184669));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__25_ (.o(regtop_dchdi_w1_hdi00[473]),
	.ck(clk),
	.d(n184668));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__26_ (.o(regtop_dchdi_w1_hdi00[474]),
	.ck(clk),
	.d(n184667));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__27_ (.o(regtop_dchdi_w1_hdi00[475]),
	.ck(clk),
	.d(n184666));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__28_ (.o(regtop_dchdi_w1_hdi00[476]),
	.ck(clk),
	.d(n184665));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__29_ (.o(regtop_dchdi_w1_hdi00[477]),
	.ck(clk),
	.d(n184664));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__30_ (.o(regtop_dchdi_w1_hdi00[478]),
	.ck(clk),
	.d(n184663));
   ms00f80 regtop_dchdi_w1_hdi00_reg_62__31_ (.o(regtop_dchdi_w1_hdi00[479]),
	.ck(clk),
	.d(n184662));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__0_ (.o(regtop_dchdi_w1_hdi00[480]),
	.ck(clk),
	.d(n184661));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__1_ (.o(regtop_dchdi_w1_hdi00[481]),
	.ck(clk),
	.d(n184660));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__2_ (.o(regtop_dchdi_w1_hdi00[482]),
	.ck(clk),
	.d(n184659));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__3_ (.o(regtop_dchdi_w1_hdi00[483]),
	.ck(clk),
	.d(n184658));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__4_ (.o(regtop_dchdi_w1_hdi00[484]),
	.ck(clk),
	.d(n184657));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__5_ (.o(regtop_dchdi_w1_hdi00[485]),
	.ck(clk),
	.d(n184656));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__6_ (.o(regtop_dchdi_w1_hdi00[486]),
	.ck(clk),
	.d(n184655));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__7_ (.o(regtop_dchdi_w1_hdi00[487]),
	.ck(clk),
	.d(n184654));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__8_ (.o(regtop_dchdi_w1_hdi00[488]),
	.ck(clk),
	.d(n184653));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__9_ (.o(regtop_dchdi_w1_hdi00[489]),
	.ck(clk),
	.d(n184652));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__10_ (.o(regtop_dchdi_w1_hdi00[490]),
	.ck(clk),
	.d(n184651));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__11_ (.o(regtop_dchdi_w1_hdi00[491]),
	.ck(clk),
	.d(n184650));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__12_ (.o(regtop_dchdi_w1_hdi00[492]),
	.ck(clk),
	.d(n184649));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__13_ (.o(regtop_dchdi_w1_hdi00[493]),
	.ck(clk),
	.d(n184648));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__14_ (.o(regtop_dchdi_w1_hdi00[494]),
	.ck(clk),
	.d(n184647));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__15_ (.o(regtop_dchdi_w1_hdi00[495]),
	.ck(clk),
	.d(n184646));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__16_ (.o(regtop_dchdi_w1_hdi00[496]),
	.ck(clk),
	.d(n184645));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__17_ (.o(regtop_dchdi_w1_hdi00[497]),
	.ck(clk),
	.d(n184644));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__18_ (.o(regtop_dchdi_w1_hdi00[498]),
	.ck(clk),
	.d(n184643));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__19_ (.o(regtop_dchdi_w1_hdi00[499]),
	.ck(clk),
	.d(n184642));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__20_ (.o(regtop_dchdi_w1_hdi00[500]),
	.ck(clk),
	.d(n184641));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__21_ (.o(regtop_dchdi_w1_hdi00[501]),
	.ck(clk),
	.d(n184640));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__22_ (.o(regtop_dchdi_w1_hdi00[502]),
	.ck(clk),
	.d(n184639));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__23_ (.o(regtop_dchdi_w1_hdi00[503]),
	.ck(clk),
	.d(n184638));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__24_ (.o(regtop_dchdi_w1_hdi00[504]),
	.ck(clk),
	.d(n184637));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__25_ (.o(regtop_dchdi_w1_hdi00[505]),
	.ck(clk),
	.d(n184636));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__26_ (.o(regtop_dchdi_w1_hdi00[506]),
	.ck(clk),
	.d(n184635));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__27_ (.o(regtop_dchdi_w1_hdi00[507]),
	.ck(clk),
	.d(n184634));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__28_ (.o(regtop_dchdi_w1_hdi00[508]),
	.ck(clk),
	.d(n184633));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__29_ (.o(regtop_dchdi_w1_hdi00[509]),
	.ck(clk),
	.d(n184632));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__30_ (.o(regtop_dchdi_w1_hdi00[510]),
	.ck(clk),
	.d(n184631));
   ms00f80 regtop_dchdi_w1_hdi00_reg_63__31_ (.o(regtop_dchdi_w1_hdi00[511]),
	.ck(clk),
	.d(n184630));
   ms00f80 regtop_g_issh_r_reg (.o(regtop_g_issh_r),
	.ck(clk),
	.d(n184629));
   ms00f80 regtop_v1_int23_n_reg (.o(v1_int23_n),
	.ck(clk),
	.d(n245090));
   ms00f80 regtop_v1_hpb_rd_reg_7_ (.o(wbb_dat_o[7]),
	.ck(clk),
	.d(n244969));
   ms00f80 regtop_v1_hpb_rd_reg_17_ (.o(wbb_dat_o[17]),
	.ck(clk),
	.d(FE_OFN470_n244978));
   ms00f80 regtop_v1_hpb_rd_reg_25_ (.o(wbb_dat_o[25]),
	.ck(clk),
	.d(FE_OFN472_n244982));
   ms00f80 regtop_v1_hpb_rd_reg_21_ (.o(wbb_dat_o[21]),
	.ck(clk),
	.d(n244980));
   ms00f80 regtop_v1_hpb_rd_reg_29_ (.o(wbb_dat_o[29]),
	.ck(clk),
	.d(n244984));
   ms00f80 regtop_v1_hpb_rd_reg_18_ (.o(wbb_dat_o[18]),
	.ck(clk),
	.d(n244979));
   ms00f80 regtop_v1_hpb_rd_reg_26_ (.o(wbb_dat_o[26]),
	.ck(clk),
	.d(n244983));
   ms00f80 regtop_v1_hpb_rd_reg_22_ (.o(wbb_dat_o[22]),
	.ck(clk),
	.d(n244981));
   ms00f80 regtop_v1_hpb_rd_reg_30_ (.o(wbb_dat_o[30]),
	.ck(clk),
	.d(n244985));
   ms00f80 regtop_v1_hpb_rd_reg_28_ (.o(wbb_dat_o[28]),
	.ck(clk),
	.d(n244221));
   ms00f80 regtop_v1_hpb_rd_reg_23_ (.o(wbb_dat_o[23]),
	.ck(clk),
	.d(n244216));
   ms00f80 regtop_v1_hpb_rd_reg_20_ (.o(wbb_dat_o[20]),
	.ck(clk),
	.d(n244219));
   ms00f80 regtop_v1_hpb_rd_reg_19_ (.o(wbb_dat_o[19]),
	.ck(clk),
	.d(n244217));
   ms00f80 regtop_v1_hpb_rd_reg_27_ (.o(wbb_dat_o[27]),
	.ck(clk),
	.d(n244215));
   ms00f80 regtop_v1_hpb_rd_reg_31_ (.o(wbb_dat_o[31]),
	.ck(clk),
	.d(n244214));
   ms00f80 regtop_v1_hpb_rd_reg_15_ (.o(wbb_dat_o[15]),
	.ck(clk),
	.d(n244977));
   ms00f80 regtop_g_prev_enfst_r_reg (.o(regtop_g_prev_enfst_r),
	.ck(clk),
	.d(regtop_N1279));
   ms00f80 regtop_g_embh_adr_r_reg_0_ (.o(regtop_g_embh_adr_r[0]),
	.ck(clk),
	.d(n170965));
   ms00f80 regtop_v1_hpb_rd_reg_8_ (.o(wbb_dat_o[8]),
	.ck(clk),
	.d(n244970));
   ms00f80 regtop_g_embh_adr_r_reg_1_ (.o(regtop_g_embh_adr_r[1]),
	.ck(clk),
	.d(n170964));
   ms00f80 regtop_v1_hpb_rd_reg_9_ (.o(wbb_dat_o[9]),
	.ck(clk),
	.d(n244971));
   ms00f80 regtop_g_embh_adr_r_reg_2_ (.o(regtop_g_embh_adr_r[2]),
	.ck(clk),
	.d(n170963));
   ms00f80 regtop_g_embh_adr_r_reg_3_ (.o(regtop_g_embh_adr_r[3]),
	.ck(clk),
	.d(n170962));
   ms00f80 regtop_g_embh_adr_r_reg_4_ (.o(regtop_g_embh_adr_r[4]),
	.ck(clk),
	.d(n170961));
   ms00f80 regtop_v1_hpb_rd_reg_12_ (.o(wbb_dat_o[12]),
	.ck(clk),
	.d(n244974));
   ms00f80 regtop_g_embh_adr_r_reg_5_ (.o(regtop_g_embh_adr_r[5]),
	.ck(clk),
	.d(n170960));
   ms00f80 regtop_v1_hpb_rd_reg_13_ (.o(wbb_dat_o[13]),
	.ck(clk),
	.d(n244975));
   ms00f80 regtop_g_embh_adr_r_reg_6_ (.o(regtop_g_embh_adr_r[6]),
	.ck(clk),
	.d(n170959));
   ms00f80 regtop_v1_hpb_rd_reg_14_ (.o(wbb_dat_o[14]),
	.ck(clk),
	.d(n244976));
   ms00f80 regtop_g_embv_adr_r_reg_0_ (.o(regtop_g_embv_adr_r[0]),
	.ck(clk),
	.d(n170958));
   ms00f80 regtop_v1_hpb_rd_reg_0_ (.o(wbb_dat_o[0]),
	.ck(clk),
	.d(n244222));
   ms00f80 regtop_g_embv_adr_r_reg_1_ (.o(regtop_g_embv_adr_r[1]),
	.ck(clk),
	.d(n170957));
   ms00f80 regtop_v1_hpb_rd_reg_1_ (.o(wbb_dat_o[1]),
	.ck(clk),
	.d(n244964));
   ms00f80 regtop_g_embv_adr_r_reg_2_ (.o(regtop_g_embv_adr_r[2]),
	.ck(clk),
	.d(n170956));
   ms00f80 regtop_v1_hpb_rd_reg_2_ (.o(wbb_dat_o[2]),
	.ck(clk),
	.d(n244965));
   ms00f80 regtop_g_embv_adr_r_reg_3_ (.o(regtop_g_embv_adr_r[3]),
	.ck(clk),
	.d(n170955));
   ms00f80 regtop_v1_hpb_rd_reg_3_ (.o(wbb_dat_o[3]),
	.ck(clk),
	.d(n244966));
   ms00f80 regtop_g_embv_adr_r_reg_4_ (.o(regtop_g_embv_adr_r[4]),
	.ck(clk),
	.d(n170954));
   ms00f80 regtop_v1_hpb_rd_reg_4_ (.o(wbb_dat_o[4]),
	.ck(clk),
	.d(n244213));
   ms00f80 regtop_g_embv_adr_r_reg_5_ (.o(regtop_g_embv_adr_r[5]),
	.ck(clk),
	.d(n170953));
   ms00f80 regtop_v1_hpb_rd_reg_5_ (.o(wbb_dat_o[5]),
	.ck(clk),
	.d(n244967));
   ms00f80 regtop_g_embv_adr_r_reg_6_ (.o(regtop_g_embv_adr_r[6]),
	.ck(clk),
	.d(n170952));
   ms00f80 regtop_v1_hpb_rd_reg_6_ (.o(wbb_dat_o[6]),
	.ck(clk),
	.d(n244968));
   ms00f80 regtop_v1_hpb_rd_reg_24_ (.o(wbb_dat_o[24]),
	.ck(clk),
	.d(n244220));
   ms00f80 regtop_g_isnf_r_reg (.o(regtop_g_isnf_r),
	.ck(clk),
	.d(n170951));
   ms00f80 regtop_v1_hpb_rd_reg_16_ (.o(wbb_dat_o[16]),
	.ck(clk),
	.d(FE_OFN468_n244218));
   ms00f80 busrtop_b_rreq_vrh_add1_r_reg_0_ (.o(busrtop_b_rreq_vrh_add1_r[0]),
	.ck(clk),
	.d(n253038));
   ms00f80 busrtop_b_rreq_vrh_add1_r_reg_1_ (.o(busrtop_b_rreq_vrh_add1_r[1]),
	.ck(clk),
	.d(busrtop_b_rreq_N423));
   ms00f80 busrtop_b_rreq_vrh_add1_r_reg_2_ (.o(busrtop_b_rreq_vrh_add1_r[2]),
	.ck(clk),
	.d(busrtop_b_rreq_N424));
   ms00f80 busrtop_b_rreq_vrh_add1_r_reg_3_ (.o(busrtop_b_rreq_vrh_add1_r[3]),
	.ck(clk),
	.d(busrtop_b_rreq_N425));
   ms00f80 busrtop_b_rreq_vrh_add1_r_reg_4_ (.o(busrtop_b_rreq_vrh_add1_r[4]),
	.ck(clk),
	.d(busrtop_b_rreq_N426));
   ms00f80 busrtop_b_rreq_vrh_add1_r_reg_5_ (.o(busrtop_b_rreq_vrh_add1_r[5]),
	.ck(clk),
	.d(busrtop_b_rreq_N427));
   ms00f80 busrtop_b_rreq_vrh_add1_r_reg_6_ (.o(busrtop_b_rreq_vrh_add1_r[6]),
	.ck(clk),
	.d(busrtop_b_rreq_N428));
   ms00f80 busrtop_b_rreq_vrh_add1_r_reg_7_ (.o(busrtop_b_rreq_vrh_add1_r[7]),
	.ck(clk),
	.d(busrtop_b_rreq_N429));
   ms00f80 busrtop_b_rreq_vrh_add1_r_reg_8_ (.o(busrtop_b_rreq_vrh_add1_r[8]),
	.ck(clk),
	.d(busrtop_b_rreq_N430));
   ms00f80 busrtop_b_rreq_vrh_add1_r_reg_9_ (.o(busrtop_b_rreq_vrh_add1_r[9]),
	.ck(clk),
	.d(busrtop_b_rreq_N431));
   ms00f80 busrtop_b_rreq_vrh_cnt_16byte_r_reg_0_ (.o(busrtop_b_rreq_vrh_cnt_16byte_r[0]),
	.ck(clk),
	.d(n170939));
   ms00f80 busrtop_b_rreq_vrh_cnt_16byte_r_reg_1_ (.o(busrtop_b_rreq_vrh_cnt_16byte_r[1]),
	.ck(clk),
	.d(n170938));
   ms00f80 busrtop_b_rreq_vrh_cnt_18byte_r_reg_0_ (.o(busrtop_b_rreq_vrh_cnt_18byte_r[0]),
	.ck(clk),
	.d(n170937));
   ms00f80 busrtop_b_rreq_vrh_cnt_18byte_r_reg_1_ (.o(busrtop_b_rreq_vrh_cnt_18byte_r[1]),
	.ck(clk),
	.d(n170932));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_27_ (.o(vh_1_ph_add[27]),
	.ck(clk),
	.d(busrtop_b_rreq_vrh_rrq_fldstatadd_r[27]));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_28_ (.o(vh_1_ph_add[28]),
	.ck(clk),
	.d(busrtop_b_rreq_vrh_rrq_fldstatadd_r[28]));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_29_ (.o(vh_1_ph_add[29]),
	.ck(clk),
	.d(busrtop_b_rreq_vrh_rrq_fldstatadd_r[29]));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_30_ (.o(vh_1_ph_add[30]),
	.ck(clk),
	.d(busrtop_b_rreq_vrh_rrq_fldstatadd_r[30]));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_31_ (.o(vh_1_ph_add[31]),
	.ck(clk),
	.d(busrtop_b_rreq_vrh_rrq_fldstatadd_r[31]));
   ms00f80 busiftop_status_b_current_reg_0_ (.o(busiftop_status_b_current_0_),
	.ck(clk),
	.d(n253125));
   ms00f80 regtop_g_isdc_r_reg (.o(regtop_g_isdc_r),
	.ck(clk),
	.d(n162088));
   ms00f80 regtop_v1_hpb_rd_reg_11_ (.o(wbb_dat_o[11]),
	.ck(clk),
	.d(n244973));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_0_ (.o(vh_1_ph_add[0]),
	.ck(clk),
	.d(n157840));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_1_ (.o(vh_1_ph_add[1]),
	.ck(clk),
	.d(n157839));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_2_ (.o(vh_1_ph_add[2]),
	.ck(clk),
	.d(n157838));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_3_ (.o(vh_1_ph_add[3]),
	.ck(clk),
	.d(n157837));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_4_ (.o(vh_1_ph_add[4]),
	.ck(clk),
	.d(n157836));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_5_ (.o(vh_1_ph_add[5]),
	.ck(clk),
	.d(n157835));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_6_ (.o(vh_1_ph_add[6]),
	.ck(clk),
	.d(n157834));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_7_ (.o(vh_1_ph_add[7]),
	.ck(clk),
	.d(n157833));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_8_ (.o(vh_1_ph_add[8]),
	.ck(clk),
	.d(n157832));
   ms00f80 busrtop_b_rreq_vh_1_ph_add_reg_9_ (.o(vh_1_ph_add[9]),
	.ck(clk),
	.d(n157831));
   ms00f80 regtop_g_isuc_r_reg (.o(regtop_g_isuc_r),
	.ck(clk),
	.d(n157815));
   ms00f80 regtop_v1_int18_n_reg (.o(v1_int18_n),
	.ck(clk),
	.d(n245091));
   ms00f80 regtop_v1_hpb_rd_reg_10_ (.o(wbb_dat_o[10]),
	.ck(clk),
	.d(n244972));
   ms00f80 busiftop_vmem_ch_r_reg (.o(busiftop_vmem_ch_r),
	.ck(clk),
	.d(vmem_ch));
   ms00f80 busiftop_vmem_add_reg_0_ (.o(vmem_add[0]),
	.ck(clk),
	.d(busiftop_N36));
   ms00f80 busiftop_vmem_add_reg_1_ (.o(vmem_add[1]),
	.ck(clk),
	.d(busiftop_N37));
   ms00f80 busiftop_vmem_add_reg_2_ (.o(vmem_add[2]),
	.ck(clk),
	.d(busiftop_N38));
   ms00f80 busiftop_vmem_add_reg_3_ (.o(vmem_add[3]),
	.ck(clk),
	.d(busiftop_N39));
   ms00f80 busiftop_vmem_add_reg_4_ (.o(vmem_add[4]),
	.ck(clk),
	.d(busiftop_N40));
   ms00f80 busiftop_vmem_add_reg_5_ (.o(vmem_add[5]),
	.ck(clk),
	.d(busiftop_N41));
   ms00f80 busiftop_vmem_add_reg_6_ (.o(vmem_add[6]),
	.ck(clk),
	.d(busiftop_N42));
   ms00f80 busiftop_vmem_add_reg_8_ (.o(vmem_add[8]),
	.ck(clk),
	.d(busiftop_N44));
   ms00f80 busiftop_vmem_add_reg_9_ (.o(vmem_add[9]),
	.ck(clk),
	.d(busiftop_N45));
   ms00f80 busiftop_vmem_add_reg_10_ (.o(vmem_add[10]),
	.ck(clk),
	.d(busiftop_N46));
   ms00f80 busiftop_vmem_add_reg_11_ (.o(vmem_add[11]),
	.ck(clk),
	.d(busiftop_N47));
   ms00f80 busiftop_vmem_add_reg_12_ (.o(vmem_add[12]),
	.ck(clk),
	.d(busiftop_N48));
   ms00f80 busiftop_vmem_add_reg_13_ (.o(vmem_add[13]),
	.ck(clk),
	.d(busiftop_N49));
   ms00f80 busiftop_vmem_add_reg_14_ (.o(vmem_add[14]),
	.ck(clk),
	.d(busiftop_N50));
   ms00f80 busiftop_vmem_add_reg_15_ (.o(vmem_add[15]),
	.ck(clk),
	.d(busiftop_N51));
   ms00f80 busiftop_vmem_add_reg_16_ (.o(vmem_add[16]),
	.ck(clk),
	.d(busiftop_N52));
   ms00f80 busiftop_vmem_add_reg_17_ (.o(vmem_add[17]),
	.ck(clk),
	.d(busiftop_N53));
   ms00f80 busiftop_vmem_add_reg_19_ (.o(vmem_add[19]),
	.ck(clk),
	.d(busiftop_N55));
   ms00f80 busiftop_vmem_add_reg_20_ (.o(vmem_add[20]),
	.ck(clk),
	.d(busiftop_N56));
   ms00f80 busiftop_vmem_add_reg_21_ (.o(vmem_add[21]),
	.ck(clk),
	.d(busiftop_N57));
   ms00f80 busiftop_vmem_add_reg_22_ (.o(vmem_add[22]),
	.ck(clk),
	.d(busiftop_N58));
   ms00f80 busiftop_vmem_add_reg_23_ (.o(vmem_add[23]),
	.ck(clk),
	.d(busiftop_N59));
   ms00f80 busiftop_vmem_add_reg_24_ (.o(vmem_add[24]),
	.ck(clk),
	.d(busiftop_N60));
   ms00f80 busiftop_vmem_add_reg_25_ (.o(vmem_add[25]),
	.ck(clk),
	.d(busiftop_N61));
   ms00f80 busiftop_vmem_ren_g_reg (.o(busiftop_vmem_ren_g),
	.ck(clk),
	.d(busiftop_N35));
   ms00f80 busiftop_vmem_add_reg_7_ (.o(vmem_add[7]),
	.ck(clk),
	.d(busiftop_N43));
   ms00f80 busiftop_vmem_add_reg_18_ (.o(vmem_add[18]),
	.ck(clk),
	.d(busiftop_N54));
   ms00f80 busiftop_vmem_data_out_reg_12_ (.o(vmem_data_out[12]),
	.ck(clk),
	.d(n244263));
   ms00f80 busiftop_vmem_data_out_reg_11_ (.o(vmem_data_out[11]),
	.ck(clk),
	.d(n244262));
   ms00f80 busiftop_vmem_data_out_reg_10_ (.o(vmem_data_out[10]),
	.ck(clk),
	.d(n253103));
   ms00f80 busiftop_vmem_data_out_reg_9_ (.o(vmem_data_out[9]),
	.ck(clk),
	.d(n253104));
   ms00f80 busiftop_vmem_data_out_reg_8_ (.o(vmem_data_out[8]),
	.ck(clk),
	.d(n253105));
   ms00f80 busiftop_vmem_data_out_reg_7_ (.o(vmem_data_out[7]),
	.ck(clk),
	.d(n253106));
   ms00f80 busiftop_vmem_data_out_reg_6_ (.o(vmem_data_out[6]),
	.ck(clk),
	.d(n253107));
   ms00f80 busiftop_vmem_data_out_reg_5_ (.o(vmem_data_out[5]),
	.ck(clk),
	.d(n253108));
   ms00f80 busiftop_vmem_data_out_reg_4_ (.o(vmem_data_out[4]),
	.ck(clk),
	.d(n253109));
   ms00f80 busiftop_vmem_data_out_reg_3_ (.o(vmem_data_out[3]),
	.ck(clk),
	.d(n253110));
   ms00f80 busiftop_vmem_data_out_reg_2_ (.o(vmem_data_out[2]),
	.ck(clk),
	.d(n253111));
   ms00f80 busiftop_vmem_data_out_reg_1_ (.o(vmem_data_out[1]),
	.ck(clk),
	.d(n253112));
   ms00f80 busiftop_vmem_data_out_reg_0_ (.o(vmem_data_out[0]),
	.ck(clk),
	.d(n253113));
   ms00f80 busiftop_vmem_data_out_reg_25_ (.o(vmem_data_out[25]),
	.ck(clk),
	.d(n244250));
   ms00f80 busiftop_vmem_data_out_reg_24_ (.o(vmem_data_out[24]),
	.ck(clk),
	.d(n253114));
   ms00f80 busiftop_vmem_data_out_reg_23_ (.o(vmem_data_out[23]),
	.ck(clk),
	.d(n253115));
   ms00f80 busiftop_vmem_data_out_reg_22_ (.o(vmem_data_out[22]),
	.ck(clk),
	.d(n253116));
   ms00f80 busiftop_vmem_data_out_reg_21_ (.o(vmem_data_out[21]),
	.ck(clk),
	.d(n253117));
   ms00f80 busiftop_vmem_data_out_reg_20_ (.o(vmem_data_out[20]),
	.ck(clk),
	.d(n244245));
   ms00f80 busiftop_vmem_data_out_reg_19_ (.o(vmem_data_out[19]),
	.ck(clk),
	.d(n253118));
   ms00f80 busiftop_vmem_data_out_reg_18_ (.o(vmem_data_out[18]),
	.ck(clk),
	.d(n253119));
   ms00f80 busiftop_vmem_data_out_reg_17_ (.o(vmem_data_out[17]),
	.ck(clk),
	.d(n253120));
   ms00f80 busiftop_vmem_data_out_reg_16_ (.o(vmem_data_out[16]),
	.ck(clk),
	.d(n253121));
   ms00f80 busiftop_vmem_data_out_reg_15_ (.o(vmem_data_out[15]),
	.ck(clk),
	.d(n253122));
   ms00f80 busiftop_vmem_data_out_reg_14_ (.o(vmem_data_out[14]),
	.ck(clk),
	.d(n253123));
   ms00f80 busiftop_vmem_data_out_reg_13_ (.o(vmem_data_out[13]),
	.ck(clk),
	.d(n253124));
   ms00f80 busiftop_vmem_wen_r_reg (.o(vmem_wen),
	.ck(clk),
	.d(busiftop_N28));
   ms00f80 busiftop_vmem_we_reg_3_ (.o(vmem_we[1]),
	.ck(clk),
	.d(busiftop_N32));
   na02f01 U261343 (.o(n211958),
	.a(n246862),
	.b(n246861));
   na02m01 U261344 (.o(n248957),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[27]));
   na02m01 U261345 (.o(n248966),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[28]));
   na02f01 U261346 (.o(n248969),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[29]));
   na02m01 U261347 (.o(n248972),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[30]));
   na02s01 U261348 (.o(n249181),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[2]));
   na02s01 U261349 (.o(n249174),
	.a(FE_OFN501_n246205),
	.b(regtop_g_wd_r[3]));
   na02s01 U261350 (.o(n249162),
	.a(FE_OFN501_n246205),
	.b(regtop_g_wd_r[5]));
   na02s01 U261351 (.o(n249157),
	.a(FE_OFN501_n246205),
	.b(regtop_g_wd_r[6]));
   na02s01 U261352 (.o(n249152),
	.a(FE_OFN501_n246205),
	.b(regtop_g_wd_r[7]));
   na02f01 U261353 (.o(n249168),
	.a(FE_OFN501_n246205),
	.b(regtop_g_wd_r[4]));
   na02f01 U261354 (.o(n249218),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[8]));
   na02f03 U261355 (.o(n249147),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[9]));
   na02s01 U261356 (.o(n249232),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[10]));
   na02f01 U261357 (.o(n249239),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[11]));
   na02f01 U261358 (.o(n249201),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[13]));
   na02s01 U261359 (.o(n249208),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[15]));
   na02f02 U261360 (.o(n249093),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[19]));
   na02f04 U261361 (.o(n249104),
	.a(FE_OFN501_n246205),
	.b(regtop_g_wd_r[20]));
   na02f02 U261362 (.o(n249124),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[21]));
   na02s01 U261363 (.o(n249194),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[0]));
   na02s01 U261364 (.o(n249187),
	.a(FE_OFN501_n246205),
	.b(regtop_g_wd_r[1]));
   na02f01 U261365 (.o(n249225),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[14]));
   na02f01 U261366 (.o(n249133),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[18]));
   na02f01 U261367 (.o(n249099),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[17]));
   na02m01 U261368 (.o(n246940),
	.a(regtop_g_udb2_r[6]),
	.b(n246939));
   in01m01 U261369 (.o(n246585),
	.a(FE_OFN366_n246266));
   in01f03 U261370 (.o(n252563),
	.a(n252561));
   no03f01 U261371 (.o(n247234),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[3]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   in01f03 U261372 (.o(n252671),
	.a(FE_OFN43_n252668));
   no02f03 U261373 (.o(n249077),
	.a(FE_OFN502_n246205),
	.b(regtop_N1990));
   na02f01 U261374 (.o(n248959),
	.a(regtop_g_paramdata_r[24]),
	.b(n248980));
   no04f04 U261376 (.o(n248676),
	.a(n248675),
	.b(n248674),
	.c(n248673),
	.d(n248672));
   no04f04 U261377 (.o(n248592),
	.a(n248591),
	.b(n248590),
	.c(n248589),
	.d(n248588));
   no04f03 U261378 (.o(n248032),
	.a(n248031),
	.b(n248030),
	.c(n248029),
	.d(n248028));
   no02s01 U261379 (.o(n249820),
	.a(n249819),
	.b(n249664));
   no04f04 U261380 (.o(n248269),
	.a(n248268),
	.b(n248267),
	.c(n248266),
	.d(n248265));
   no04f02 U261381 (.o(n247696),
	.a(n247695),
	.b(n247694),
	.c(n247693),
	.d(n247692));
   no04f03 U261382 (.o(n247780),
	.a(n247779),
	.b(FE_OFN554_n247778),
	.c(n247777),
	.d(n247776));
   no04f06 U261383 (.o(n247822),
	.a(n247821),
	.b(n247820),
	.c(n247819),
	.d(n247818));
   no04f04 U261384 (.o(n248550),
	.a(FE_OFN382_n248549),
	.b(n248548),
	.c(n248547),
	.d(n248546));
   no04f03 U261385 (.o(n248634),
	.a(n248633),
	.b(n248632),
	.c(n248631),
	.d(n248630));
   no04f04 U261386 (.o(n248227),
	.a(n248226),
	.b(n248225),
	.c(n248224),
	.d(n248223));
   na02s01 U261387 (.o(n246003),
	.a(n252485),
	.b(regtop_g_nfst_r[2]));
   no03f01 U261388 (.o(n247587),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[2]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no04f02 U261389 (.o(n247865),
	.a(n247843),
	.b(n247842),
	.c(n247841),
	.d(n247840));
   no04f02 U261390 (.o(n248951),
	.a(n248897),
	.b(n248896),
	.c(n248895),
	.d(n248894));
   na02m01 U261391 (.o(n245610),
	.a(n245609),
	.b(n245608));
   no03f01 U261392 (.o(n249766),
	.a(n249765),
	.b(n249664),
	.c(n249764));
   na02f01 U261393 (.o(n246873),
	.a(regtop_g_udb2_r[4]),
	.b(n246939));
   na02s01 U261394 (.o(n246911),
	.a(n247053),
	.b(n246910));
   no02s01 U261395 (.o(n249432),
	.a(n249430),
	.b(n249429));
   na02f01 U261396 (.o(n246862),
	.a(regtop_g_udb2_r[3]),
	.b(n246877));
   na02s01 U261397 (.o(n246906),
	.a(n247042),
	.b(n246905));
   no02f02 U261398 (.o(n249479),
	.a(n249477),
	.b(n249476));
   no02f02 U261399 (.o(n249491),
	.a(n249489),
	.b(n249488));
   no02f01 U261400 (.o(n249195),
	.a(n249193),
	.b(n249192));
   na04f01 U261401 (.o(n246872),
	.a(n246880),
	.b(n246871),
	.c(regtop_g_udb2_r[3]),
	.d(n246935));
   no02f01 U261402 (.o(n249447),
	.a(n249445),
	.b(n249444));
   no02f02 U261403 (.o(n249188),
	.a(n249186),
	.b(n249185));
   no04f02 U261404 (.o(n247584),
	.a(n247562),
	.b(n247561),
	.c(n247560),
	.d(n247559));
   no04f02 U261405 (.o(n247542),
	.a(n247518),
	.b(n247517),
	.c(n247516),
	.d(n247515));
   no04f04 U261406 (.o(n247123),
	.a(n247122),
	.b(n247121),
	.c(n247120),
	.d(n247119));
   no04f02 U261407 (.o(n247440),
	.a(n247416),
	.b(n247415),
	.c(n247414),
	.d(n247413));
   no04f02 U261408 (.o(n248424),
	.a(n248423),
	.b(n248422),
	.c(n248421),
	.d(n248420));
   no03f01 U261409 (.o(n249541),
	.a(n249539),
	.b(n249538),
	.c(n249537));
   no04f01 U261410 (.o(n247124),
	.a(n247090),
	.b(n247089),
	.c(n247088),
	.d(n247087));
   na03s01 U261411 (.o(n246691),
	.a(n246690),
	.b(n246689),
	.c(n246688));
   no03f01 U261412 (.o(n247376),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[0]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   ao12f01 U261413 (.o(n249202),
	.a(n249200),
	.b(n249252),
	.c(regtop_g_usrd_r[13]));
   ao22f02 U261414 (.o(n245596),
	.a(regtop_g_icnf_r),
	.b(n245592),
	.c(regtop_g_wd_r[16]),
	.d(n252269));
   ao12f02 U261415 (.o(n249380),
	.a(n249379),
	.b(regtop_g_mem_rd2_r[26]),
	.c(regtop_g_memr_ok_r));
   no03f01 U261416 (.o(n247380),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[1]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   ao22f01 U261417 (.o(n246934),
	.a(n246933),
	.b(n246932),
	.c(regtop_g_udb1_r[6]),
	.d(n246931));
   na02f01 U261421 (.o(n246939),
	.a(n246870),
	.b(n246869));
   na03f02 U261422 (.o(n249620),
	.a(n249619),
	.b(n249618),
	.c(n249617));
   na03f01 U261423 (.o(n247379),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247378));
   na04f02 U261424 (.o(n249750),
	.a(n249743),
	.b(n249742),
	.c(n249741),
	.d(n249740));
   na04f04 U261425 (.o(n248484),
	.a(n248483),
	.b(n248482),
	.c(n248481),
	.d(n248480));
   na04f04 U261426 (.o(n248652),
	.a(n248651),
	.b(n248650),
	.c(n248649),
	.d(n248648));
   na04f02 U261427 (.o(n248822),
	.a(n248811),
	.b(n248810),
	.c(n248809),
	.d(n248808));
   na04f02 U261428 (.o(n248445),
	.a(n248429),
	.b(n248428),
	.c(n248427),
	.d(n248426));
   na04f02 U261429 (.o(n248053),
	.a(n248037),
	.b(n248036),
	.c(n248035),
	.d(n248034));
   na04f02 U261430 (.o(n248095),
	.a(n248079),
	.b(n248078),
	.c(n248077),
	.d(n248076));
   na04f02 U261431 (.o(n248697),
	.a(n248681),
	.b(n248680),
	.c(n248679),
	.d(n248678));
   na04f01 U261432 (.o(n248739),
	.a(n248723),
	.b(n248722),
	.c(n248721),
	.d(n248720));
   na04f03 U261433 (.o(n248781),
	.a(n248765),
	.b(n248764),
	.c(n248763),
	.d(n248762));
   na04m01 U261434 (.o(n248571),
	.a(n248555),
	.b(n248554),
	.c(n248553),
	.d(n248552));
   na04f01 U261435 (.o(n248011),
	.a(n247995),
	.b(n247994),
	.c(n247993),
	.d(n247992));
   na04f03 U261436 (.o(n249707),
	.a(n249695),
	.b(n249694),
	.c(n249693),
	.d(n249692));
   na04f02 U261437 (.o(n249577),
	.a(n249571),
	.b(n249570),
	.c(n249569),
	.d(n249568));
   na04f03 U261438 (.o(n248823),
	.a(n248807),
	.b(n248806),
	.c(n248805),
	.d(n248804));
   no02f01 U261439 (.o(n249048),
	.a(n249047),
	.b(n249046));
   na04f02 U261440 (.o(n248245),
	.a(n248244),
	.b(n248243),
	.c(n248242),
	.d(n248241));
   na04f04 U261441 (.o(n247863),
	.a(n247847),
	.b(n247846),
	.c(n247845),
	.d(n247844));
   na04f04 U261442 (.o(n248308),
	.a(n248302),
	.b(n248301),
	.c(n248300),
	.d(n248299));
   na04f06 U261443 (.o(n248310),
	.a(n248294),
	.b(n248293),
	.c(n248292),
	.d(n248291));
   na04f06 U261444 (.o(n248287),
	.a(n248286),
	.b(n248285),
	.c(n248284),
	.d(n248283));
   na04f06 U261445 (.o(n248947),
	.a(n248933),
	.b(n248932),
	.c(n248931),
	.d(n248930));
   na04f03 U261446 (.o(n248949),
	.a(n248909),
	.b(n248908),
	.c(n248907),
	.d(n248906));
   na04f03 U261447 (.o(n247646),
	.a(n247645),
	.b(n247644),
	.c(n247643),
	.d(n247642));
   na04f03 U261448 (.o(n247798),
	.a(n247797),
	.b(n247796),
	.c(n247795),
	.d(n247794));
   na04f02 U261449 (.o(n247903),
	.a(n247897),
	.b(n247896),
	.c(n247895),
	.d(n247894));
   na04f02 U261451 (.o(n248115),
	.a(n248099),
	.b(n248098),
	.c(n248097),
	.d(n248096));
   na04f04 U261452 (.o(n248759),
	.a(n248743),
	.b(n248742),
	.c(n248741),
	.d(n248740));
   na04f04 U261453 (.o(n248350),
	.a(n248344),
	.b(n248343),
	.c(n248342),
	.d(n248341));
   na04f02 U261454 (.o(n248352),
	.a(n248336),
	.b(n248335),
	.c(n248334),
	.d(n248333));
   na04f02 U261455 (.o(n248329),
	.a(n248328),
	.b(n248327),
	.c(n248326),
	.d(n248325));
   na04f04 U261456 (.o(n248801),
	.a(n248785),
	.b(n248784),
	.c(n248783),
	.d(n248782));
   na04f03 U261457 (.o(n248799),
	.a(n248793),
	.b(n248792),
	.c(n248791),
	.d(n248790));
   na04f03 U261458 (.o(n248526),
	.a(n248525),
	.b(n248524),
	.c(n248523),
	.d(n248522));
   na04f06 U261459 (.o(n248203),
	.a(n248202),
	.b(n248201),
	.c(n248200),
	.d(n248199));
   na02s01 U261460 (.o(n249131),
	.a(n249130),
	.b(n249129));
   na02s01 U261461 (.o(n249092),
	.a(n249091),
	.b(n249090));
   na04f03 U261462 (.o(n249680),
	.a(n249672),
	.b(n249671),
	.c(n249670),
	.d(n249669));
   na04f06 U261463 (.o(n248246),
	.a(n248240),
	.b(n248239),
	.c(n248238),
	.d(n248237));
   na04f04 U261464 (.o(n248147),
	.a(n248137),
	.b(n248136),
	.c(n248135),
	.d(n248134));
   na04f02 U261465 (.o(n247862),
	.a(n247851),
	.b(n247850),
	.c(n247849),
	.d(n247848));
   na04f03 U261466 (.o(n248309),
	.a(n248298),
	.b(n248297),
	.c(n248296),
	.d(n248295));
   na04f02 U261467 (.o(n248307),
	.a(n248306),
	.b(n248305),
	.c(n248304),
	.d(n248303));
   na04f02 U261468 (.o(n248288),
	.a(n248282),
	.b(n248281),
	.c(n248280),
	.d(n248279));
   na04f01 U261469 (.o(n248289),
	.a(n248278),
	.b(n248277),
	.c(n248276),
	.d(n248275));
   na04f04 U261470 (.o(n248948),
	.a(n248921),
	.b(n248920),
	.c(n248919),
	.d(n248918));
   na04f06 U261471 (.o(n247758),
	.a(n247747),
	.b(n247746),
	.c(n247745),
	.d(n247744));
   na04f04 U261472 (.o(n247799),
	.a(n247793),
	.b(n247792),
	.c(n247791),
	.d(n247790));
   na04f01 U261473 (.o(n247884),
	.a(n247873),
	.b(n247872),
	.c(n247871),
	.d(n247870));
   na04f06 U261474 (.o(n247883),
	.a(n247877),
	.b(n247876),
	.c(n247875),
	.d(n247874));
   na04f02 U261475 (.o(n247904),
	.a(n247893),
	.b(n247892),
	.c(n247891),
	.d(n247890));
   na04f03 U261476 (.o(n247902),
	.a(n247901),
	.b(n247900),
	.c(n247899),
	.d(n247898));
   na04f04 U261477 (.o(n248462),
	.a(n248461),
	.b(n248460),
	.c(n248459),
	.d(n248458));
   na04f04 U261478 (.o(n248112),
	.a(n248111),
	.b(n248110),
	.c(n248109),
	.d(n248108));
   na04f04 U261479 (.o(n248758),
	.a(n248747),
	.b(n248746),
	.c(n248745),
	.d(n248744));
   na04f02 U261480 (.o(n248351),
	.a(n248340),
	.b(n248339),
	.c(n248338),
	.d(n248337));
   na04f04 U261481 (.o(n248349),
	.a(n248348),
	.b(n248347),
	.c(n248346),
	.d(n248345));
   na04f06 U261482 (.o(n248330),
	.a(n248324),
	.b(n248323),
	.c(n248322),
	.d(n248321));
   na04f03 U261483 (.o(n248331),
	.a(n248320),
	.b(n248319),
	.c(n248318),
	.d(n248317));
   na04f06 U261484 (.o(n248800),
	.a(n248789),
	.b(n248788),
	.c(n248787),
	.d(n248786));
   na04f02 U261485 (.o(n248612),
	.a(n248601),
	.b(n248600),
	.c(n248599),
	.d(n248598));
   na04f06 U261486 (.o(n248204),
	.a(n248198),
	.b(n248197),
	.c(n248196),
	.d(n248195));
   na04f01 U261487 (.o(n248247),
	.a(n248236),
	.b(n248235),
	.c(n248234),
	.d(n248233));
   na04f02 U261488 (.o(n247800),
	.a(n247789),
	.b(n247788),
	.c(n247787),
	.d(n247786));
   na04f02 U261489 (.o(n248205),
	.a(n248194),
	.b(n248193),
	.c(n248192),
	.d(n248191));
   na04f03 U261490 (.o(n248423),
	.a(n248397),
	.b(n248396),
	.c(n248395),
	.d(n248394));
   na04f04 U261491 (.o(n249681),
	.a(n249668),
	.b(n249667),
	.c(n249666),
	.d(n249665));
   na04f04 U261492 (.o(n249600),
	.a(n249599),
	.b(n249598),
	.c(n249597),
	.d(n249596));
   na04f01 U261493 (.o(n248248),
	.a(n248232),
	.b(n248231),
	.c(n248230),
	.d(n248229));
   na04f01 U261494 (.o(n247649),
	.a(n247614),
	.b(n247613),
	.c(n247612),
	.d(n247611));
   na04f04 U261495 (.o(n247759),
	.a(n247743),
	.b(n247742),
	.c(n247741),
	.d(n247740));
   na04f02 U261496 (.o(n247801),
	.a(n247785),
	.b(n247784),
	.c(n247783),
	.d(n247782));
   na04f02 U261497 (.o(n247885),
	.a(n247869),
	.b(n247868),
	.c(n247867),
	.d(n247866));
   na04f01 U261498 (.o(n248529),
	.a(n248513),
	.b(n248512),
	.c(n248511),
	.d(n248510));
   na04f06 U261499 (.o(n248613),
	.a(n248597),
	.b(n248596),
	.c(n248595),
	.d(n248594));
   na04f02 U261500 (.o(n248206),
	.a(n248190),
	.b(n248189),
	.c(n248188),
	.d(n248187));
   na04f03 U261501 (.o(n247715),
	.a(n247709),
	.b(n247708),
	.c(n247707),
	.d(n247706));
   na04f06 U261502 (.o(n247925),
	.a(n247919),
	.b(n247918),
	.c(n247917),
	.d(n247916));
   na04f03 U261503 (.o(n248443),
	.a(n248437),
	.b(n248436),
	.c(n248435),
	.d(n248434));
   na04f03 U261504 (.o(n248051),
	.a(n248045),
	.b(n248044),
	.c(n248043),
	.d(n248042));
   na04f02 U261505 (.o(n248093),
	.a(n248087),
	.b(n248086),
	.c(n248085),
	.d(n248084));
   na04f01 U261506 (.o(n248695),
	.a(n248689),
	.b(n248688),
	.c(n248687),
	.d(n248686));
   na04f02 U261507 (.o(n248737),
	.a(n248731),
	.b(n248730),
	.c(n248729),
	.d(n248728));
   na04f04 U261508 (.o(n248779),
	.a(n248773),
	.b(n248772),
	.c(n248771),
	.d(n248770));
   na04f02 U261509 (.o(n248569),
	.a(n248563),
	.b(n248562),
	.c(n248561),
	.d(n248560));
   na04f03 U261510 (.o(n248009),
	.a(n248003),
	.b(n248002),
	.c(n248001),
	.d(n248000));
   na04f06 U261511 (.o(n248387),
	.a(n248386),
	.b(n248385),
	.c(n248384),
	.d(n248383));
   na04f02 U261512 (.o(n249622),
	.a(n249613),
	.b(n249612),
	.c(n249611),
	.d(n249610));
   na04f03 U261513 (.o(n248485),
	.a(n248479),
	.b(n248478),
	.c(n248477),
	.d(n248476));
   na04f02 U261514 (.o(n248653),
	.a(n248647),
	.b(n248646),
	.c(n248645),
	.d(n248644));
   na03s01 U261515 (.o(n249464),
	.a(n249463),
	.b(n249462),
	.c(n249461));
   na04f02 U261516 (.o(n248390),
	.a(n248361),
	.b(n248360),
	.c(n248359),
	.d(n248358));
   na04f02 U261517 (.o(n248389),
	.a(n248368),
	.b(n248367),
	.c(n248366),
	.d(n248365));
   na04f03 U261518 (.o(n249751),
	.a(n249737),
	.b(n249736),
	.c(n249735),
	.d(n249734));
   na04f06 U261519 (.o(n248182),
	.a(n248172),
	.b(n248171),
	.c(n248170),
	.d(n248169));
   na04f03 U261520 (.o(n249708),
	.a(n249691),
	.b(n249690),
	.c(n249689),
	.d(n249688));
   na04f01 U261521 (.o(n249477),
	.a(n249471),
	.b(n249470),
	.c(n249469),
	.d(FE_OFN388_n249468));
   na04f01 U261522 (.o(n249489),
	.a(n249483),
	.b(n249482),
	.c(n249481),
	.d(FE_OFN390_n249480));
   oa12f04 U261523 (.o(n249255),
	.a(n247029),
	.b(n247031),
	.c(n247030));
   na04f02 U261524 (.o(n249678),
	.a(n249677),
	.b(n249676),
	.c(n249675),
	.d(n249674));
   na02s01 U261525 (.o(n245864),
	.a(n245863),
	.b(n245862));
   na04f04 U261526 (.o(n249601),
	.a(n249595),
	.b(n249594),
	.c(n249593),
	.d(n249592));
   no02f01 U261527 (.o(n248997),
	.a(n249031),
	.b(n248995));
   na04f06 U261528 (.o(n247560),
	.a(n247554),
	.b(n247553),
	.c(n247552),
	.d(n247551));
   na04f03 U261529 (.o(n247516),
	.a(n247508),
	.b(n247507),
	.c(n247506),
	.d(n247505));
   na04f02 U261530 (.o(n247581),
	.a(n247570),
	.b(n247569),
	.c(n247568),
	.d(n247567));
   na04f03 U261531 (.o(n247414),
	.a(n247407),
	.b(n247406),
	.c(n247405),
	.d(n247404));
   na04f04 U261532 (.o(n248388),
	.a(n248379),
	.b(n248378),
	.c(n248377),
	.d(n248376));
   na04f01 U261533 (.o(n249393),
	.a(n249387),
	.b(n249386),
	.c(n249385),
	.d(n249384));
   na04f04 U261534 (.o(n247088),
	.a(n247080),
	.b(n247079),
	.c(n247078),
	.d(n247077));
   na04f04 U261535 (.o(n247121),
	.a(n247105),
	.b(n247104),
	.c(n247103),
	.d(n247102));
   na04f02 U261536 (.o(n247438),
	.a(n247421),
	.b(n247420),
	.c(n247419),
	.d(n247418));
   na04m01 U261537 (.o(n247416),
	.a(n247398),
	.b(n247397),
	.c(n247396),
	.d(n247395));
   na04f02 U261538 (.o(n249705),
	.a(n249704),
	.b(n249703),
	.c(n249702),
	.d(n249701));
   na03f03 U261539 (.o(n249505),
	.a(n249494),
	.b(n249493),
	.c(n249492));
   na04f01 U261540 (.o(n249430),
	.a(n249424),
	.b(n249423),
	.c(n249422),
	.d(n249421));
   na04f04 U261541 (.o(n247580),
	.a(n247574),
	.b(n247573),
	.c(n247572),
	.d(n247571));
   na04f02 U261542 (.o(n248421),
	.a(n248412),
	.b(n248411),
	.c(n248410),
	.d(n248409));
   na04f01 U261543 (.o(n249465),
	.a(n249460),
	.b(n249459),
	.c(n249458),
	.d(n249457));
   na04f02 U261544 (.o(n248148),
	.a(n248133),
	.b(n248132),
	.c(n248131),
	.d(n248130));
   na04f02 U261545 (.o(n248149),
	.a(n248125),
	.b(n248124),
	.c(n248123),
	.d(n248122));
   na04f02 U261546 (.o(n248183),
	.a(n248166),
	.b(n248165),
	.c(n248164),
	.d(n248163));
   na04f02 U261547 (.o(n248181),
	.a(n248180),
	.b(n248179),
	.c(n248178),
	.d(n248177));
   na04f02 U261548 (.o(n247538),
	.a(n247530),
	.b(n247529),
	.c(n247528),
	.d(n247527));
   na04f02 U261549 (.o(n247120),
	.a(n247113),
	.b(n247112),
	.c(n247111),
	.d(n247110));
   na04f04 U261550 (.o(n247559),
	.a(n247558),
	.b(n247557),
	.c(n247556),
	.d(n247555));
   na04f03 U261551 (.o(n247515),
	.a(n247514),
	.b(n247513),
	.c(n247512),
	.d(n247511));
   na04f04 U261552 (.o(n247413),
	.a(n247412),
	.b(n247411),
	.c(n247410),
	.d(n247409));
   na04f02 U261553 (.o(n247561),
	.a(n247550),
	.b(n247549),
	.c(n247548),
	.d(n247547));
   na04f02 U261554 (.o(n247562),
	.a(n247546),
	.b(n247545),
	.c(n247544),
	.d(n247543));
   na04f03 U261555 (.o(n247579),
	.a(n247578),
	.b(n247577),
	.c(n247576),
	.d(n247575));
   na04f06 U261556 (.o(n247582),
	.a(n247566),
	.b(n247565),
	.c(n247564),
	.d(n247563));
   na04f04 U261557 (.o(n247517),
	.a(n247504),
	.b(n247503),
	.c(n247502),
	.d(n247501));
   na04f01 U261558 (.o(n247518),
	.a(n247500),
	.b(n247499),
	.c(n247498),
	.d(n247497));
   na04f01 U261559 (.o(n247090),
	.a(n247066),
	.b(n247065),
	.c(n247064),
	.d(n247063));
   na04f02 U261560 (.o(n247122),
	.a(n247098),
	.b(n247097),
	.c(n247096),
	.d(n247095));
   na04f01 U261561 (.o(n249562),
	.a(n249556),
	.b(n249555),
	.c(n249554),
	.d(n249553));
   na04f02 U261562 (.o(n247537),
	.a(n247536),
	.b(n247535),
	.c(n247534),
	.d(n247533));
   na04f02 U261563 (.o(n247089),
	.a(n247073),
	.b(n247072),
	.c(n247071),
	.d(n247070));
   na04f02 U261564 (.o(n247415),
	.a(n247403),
	.b(n247402),
	.c(n247401),
	.d(n247400));
   na04f02 U261565 (.o(n249522),
	.a(n249511),
	.b(n249510),
	.c(n249509),
	.d(n249508));
   na04f01 U261566 (.o(n249418),
	.a(n249412),
	.b(n249411),
	.c(n249410),
	.d(n249409));
   na04f03 U261567 (.o(n247435),
	.a(n247434),
	.b(n247433),
	.c(n247432),
	.d(n247431));
   na02s01 U261568 (.o(n249118),
	.a(n249117),
	.b(n249116));
   na04f01 U261569 (.o(n249539),
	.a(n249528),
	.b(n249527),
	.c(n249526),
	.d(n249525));
   na04s01 U261570 (.o(n249576),
	.a(n249575),
	.b(n249574),
	.c(n249573),
	.d(n249572));
   na04f02 U261571 (.o(n252242),
	.a(n252241),
	.b(n252312),
	.c(n252816),
	.d(n252750));
   na04f01 U261572 (.o(n249623),
	.a(n249609),
	.b(n249608),
	.c(n249685),
	.d(n249607));
   na04f03 U261573 (.o(n245509),
	.a(n245508),
	.b(n245507),
	.c(n245506),
	.d(n245505));
   no02f02 U261574 (.o(regtop_N1990),
	.a(n249113),
	.b(n252232));
   na02f01 U261575 (.o(n252728),
	.a(n252731),
	.b(n252711));
   na02f02 U261576 (.o(n252305),
	.a(n252377),
	.b(n252260));
   na02m01 U261577 (.o(n246874),
	.a(n246880),
	.b(n246859));
   na02f01 U261579 (.o(n246869),
	.a(n246880),
	.b(n246935));
   na02f01 U261580 (.o(n252748),
	.a(n252731),
	.b(n252730));
   no02s01 U261581 (.o(n252276),
	.a(n252275),
	.b(n252274));
   no02f02 U261582 (.o(n246838),
	.a(n249064),
	.b(n246352));
   na02f10 U261583 (.o(n252540),
	.a(n252523),
	.b(FE_OFN45_n252700));
   na02f01 U261584 (.o(n252257),
	.a(n252302),
	.b(regtop_g_ferror_r));
   no02f01 U261585 (.o(n249145),
	.a(n249144),
	.b(n249143));
   na02f02 U261586 (.o(n252602),
	.a(n252601),
	.b(n246909));
   no03s01 U261587 (.o(n252258),
	.a(n252250),
	.b(regtop_g_tmg_ferr_hit_r),
	.c(n252249));
   na02f01 U261588 (.o(n252996),
	.a(n253015),
	.b(n252972));
   ao12f01 U261589 (.o(n249927),
	.a(n252260),
	.b(regtop_g_prev_enfst_r),
	.c(n252948));
   oa12f02 U261591 (.o(n246896),
	.a(v_vldstatus_r[4]),
	.b(n246894),
	.c(n246893));
   na02f06 U261595 (.o(n252698),
	.a(n252687),
	.b(n252686));
   in01f08 U261596 (.o(n251619),
	.a(FE_OFN327_n251600));
   in01f08 U261597 (.o(n250484),
	.a(FE_OFN284_n250466));
   in01f06 U261598 (.o(n251229),
	.a(FE_OFN422_n251211));
   no02f02 U261599 (.o(n249317),
	.a(n246002),
	.b(FE_OFN492_n252377));
   in01f06 U261600 (.o(n250018),
	.a(FE_OFN402_n249999));
   in01f08 U261601 (.o(n252011),
	.a(FE_OFN434_n251996));
   na02s01 U261602 (.o(n246894),
	.a(n246888),
	.b(n247003));
   na02m02 U261603 (.o(n246893),
	.a(n246892),
	.b(n247015));
   na02f01 U261604 (.o(n249143),
	.a(n249142),
	.b(n249141));
   na02m02 U261605 (.o(n246978),
	.a(n246974),
	.b(n246973));
   no02f02 U261606 (.o(n249064),
	.a(y1_bs_wait_n),
	.b(FE_OFN68_n247591));
   na04f02 U261607 (.o(n249776),
	.a(n249775),
	.b(n249774),
	.c(n249773),
	.d(n249772));
   no02s01 U261608 (.o(n246230),
	.a(n253125),
	.b(n246233));
   na03s01 U261609 (.o(n245536),
	.a(n252826),
	.b(n252371),
	.c(n252604));
   na04f01 U261610 (.o(n245504),
	.a(n245496),
	.b(n245495),
	.c(n245494),
	.d(n245493));
   na02f02 U261611 (.o(n252510),
	.a(n252403),
	.b(n252384));
   na02f04 U261612 (.o(n249247),
	.a(n252596),
	.b(FE_OFN218_n246238));
   no02f03 U261613 (.o(n250144),
	.a(FE_OFN22_n250202),
	.b(n252122));
   no02m02 U261614 (.o(n247006),
	.a(n247005),
	.b(n247004));
   no02f01 U261615 (.o(n246002),
	.a(n252948),
	.b(FE_OFN439_n252264));
   in01f02 U261616 (.o(n252813),
	.a(FE_OFN6_n246618));
   na02f04 U261617 (.o(n252811),
	.a(n249135),
	.b(n249137));
   na02s01 U261618 (.o(n246976),
	.a(n246975),
	.b(n246723));
   na02s01 U261619 (.o(n249138),
	.a(n249137),
	.b(n249136));
   na02f01 U261620 (.o(n252252),
	.a(regtop_g_paramadr_r[6]),
	.b(n245581));
   no02f01 U261622 (.o(n246892),
	.a(n247028),
	.b(n247018));
   in01f01 U261623 (.o(n247125),
	.a(n247146));
   na03f01 U261624 (.o(n252832),
	.a(n252831),
	.b(n252866),
	.c(FE_OFN507_regtop_g_a_r_4_));
   na02f03 U261625 (.o(n245940),
	.a(n245939),
	.b(n252352));
   in01m01 U261626 (.o(n252448),
	.a(n252403));
   na02m01 U261627 (.o(n249863),
	.a(n249870),
	.b(vh_1_ph_add[7]));
   no02f02 U261628 (.o(n246956),
	.a(n246959),
	.b(n246912));
   na02s01 U261629 (.o(n252424),
	.a(n252462),
	.b(regtop_g_paramadr_r[6]));
   ao12f01 U261630 (.o(n249214),
	.a(n249213),
	.b(FE_OFN551_n249140),
	.c(regtop_g_atscd_r[8]));
   ao12m01 U261631 (.o(n249019),
	.a(n246895),
	.b(vldtop_vld_syndec_vld_vscdet_v_seqerr_r),
	.c(v_vldstatus_r[0]));
   na02f02 U261632 (.o(n252958),
	.a(n245447),
	.b(n245593));
   na02f03 U261633 (.o(n252050),
	.a(n250055),
	.b(n250201));
   na02f04 U261634 (.o(n252122),
	.a(n250128),
	.b(n250200));
   na02f04 U261635 (.o(n252196),
	.a(n250201),
	.b(n250200));
   no02f01 U261636 (.o(n248167),
	.a(n247109),
	.b(n250770));
   na03f01 U261637 (.o(n252159),
	.a(regtop_v1_hdi00_a[0]),
	.b(n250200),
	.c(n250164));
   no02f10 U261638 (.o(n248140),
	.a(n247082),
	.b(FE_OFN556_n250770));
   no02f01 U261639 (.o(n248356),
	.a(n247062),
	.b(n251053));
   no02f02 U261640 (.o(n249645),
	.a(regtop_g_a_r[7]),
	.b(n246204));
   no02m01 U261641 (.o(n252403),
	.a(n252382),
	.b(n252381));
   in01f03 U261642 (.o(n252523),
	.a(n252575));
   in01f02 U261643 (.o(n252567),
	.a(n252752));
   in01f04 U261644 (.o(n249823),
	.a(n245446));
   na02s01 U261645 (.o(n246883),
	.a(n246055),
	.b(n245986));
   no02s01 U261646 (.o(n246847),
	.a(n252254),
	.b(n252574));
   in01f02 U261647 (.o(n252352),
	.a(n245938));
   na02s01 U261648 (.o(n246233),
	.a(n246229),
	.b(busrtop_b_rreq_vrh_cnt_18byte_r[1]));
   no02f02 U261649 (.o(n252596),
	.a(regtop_g_adb_r[0]),
	.b(n252599));
   na02s01 U261650 (.o(n249316),
	.a(n249315),
	.b(n249314));
   na02f02 U261651 (.o(n252341),
	.a(regtop_g_paramadr_r[2]),
	.b(n245761));
   na02s01 U261652 (.o(n245820),
	.a(vh_1_ph_add[8]),
	.b(vh_1_ph_add[9]));
   na02f06 U261653 (.o(n245620),
	.a(n245417),
	.b(n245416));
   na02f06 U261654 (.o(n247082),
	.a(n249948),
	.b(n247081));
   na02f03 U261655 (.o(n247114),
	.a(n249948),
	.b(n250201));
   na03f10 U261656 (.o(n251621),
	.a(regtop_v1_hdi00_a[4]),
	.b(n247060),
	.c(n247056));
   no02s01 U261657 (.o(n247019),
	.a(n247018),
	.b(n247017));
   na02f03 U261658 (.o(n249827),
	.a(FE_OFN4_n245443),
	.b(n252874));
   na02s01 U261659 (.o(n245446),
	.a(FE_OFN4_n245443),
	.b(n249628));
   na02f01 U261660 (.o(n245477),
	.a(n245488),
	.b(FE_OFN520_regtop_g_a_r_6_));
   na02f02 U261661 (.o(n246889),
	.a(n246677),
	.b(n246676));
   na02f02 U261662 (.o(n245448),
	.a(n245447),
	.b(n252831));
   no02m03 U261663 (.o(n250200),
	.a(regtop_v1_hdi00_a[2]),
	.b(FE_OFN497_n249947));
   na02m01 U261664 (.o(n247001),
	.a(n246999),
	.b(n247024));
   no02m02 U261665 (.o(n246983),
	.a(n246982),
	.b(n246981));
   na03f01 U261666 (.o(n247076),
	.a(regtop_v1_hdi00_a[2]),
	.b(regtop_v1_hdi00_a[0]),
	.c(regtop_v1_hdi00_a[1]));
   na03f01 U261667 (.o(n251337),
	.a(regtop_v1_hdi00_a[3]),
	.b(regtop_v1_hdi00_a[4]),
	.c(n247056));
   na02s01 U261668 (.o(n245463),
	.a(FE_OFN4_n245443),
	.b(n249638));
   na02f03 U261669 (.o(n249828),
	.a(FE_OFN4_n245443),
	.b(n249639));
   in01m01 U261670 (.o(n245593),
	.a(n245481));
   na02f02 U261671 (.o(n245460),
	.a(FE_OFN4_n245443),
	.b(n249629));
   na03f01 U261672 (.o(n250486),
	.a(regtop_v1_hdi00_a[5]),
	.b(regtop_v1_hdi00_a[4]),
	.c(n247060));
   na02s01 U261673 (.o(n245938),
	.a(n252462),
	.b(n252379));
   na02f08 U261674 (.o(n251053),
	.a(regtop_v1_hdi00_a[5]),
	.b(n247055));
   na02f10 U261675 (.o(n250770),
	.a(regtop_v1_hdi00_a[5]),
	.b(n247061));
   na02f03 U261676 (.o(n247062),
	.a(regtop_v1_hdi00_a[0]),
	.b(n247091));
   na02m02 U261677 (.o(n249878),
	.a(n249885),
	.b(vh_1_ph_add[5]));
   na02f03 U261678 (.o(n247069),
	.a(regtop_v1_hdi00_a[2]),
	.b(n247081));
   na02f04 U261679 (.o(n247101),
	.a(regtop_v1_hdi00_a[2]),
	.b(n250201));
   na02f03 U261680 (.o(n249140),
	.a(n252591),
	.b(FE_OFN218_n246238));
   na02f01 U261681 (.o(n252820),
	.a(n245551),
	.b(n252238));
   no04s01 U261682 (.o(n246722),
	.a(n246705),
	.b(n246704),
	.c(n246703),
	.d(n246702));
   na02f01 U261683 (.o(n251904),
	.a(regtop_v1_hdi00_a[3]),
	.b(n247059));
   ao12f02 U261685 (.o(n246985),
	.a(n246387),
	.b(n246389),
	.c(n246388));
   na02s01 U261686 (.o(n246201),
	.a(n253015),
	.b(regtop_g_dmod_r));
   na02s01 U261687 (.o(n252383),
	.a(regtop_g_paramadr_r[2]),
	.b(regtop_g_paramadr_r[3]));
   na02m01 U261688 (.o(n252381),
	.a(n252380),
	.b(n252379));
   no02f02 U261689 (.o(n250128),
	.a(regtop_v1_hdi00_a[0]),
	.b(n250164));
   no02s01 U261690 (.o(n246853),
	.a(vldtop_vld_syndec_vld_vlfeed_dselect_r),
	.b(n247146));
   no02f01 U261691 (.o(n249636),
	.a(n249698),
	.b(n245461));
   no02f02 U261692 (.o(n247081),
	.a(FE_OFN516_regtop_v1_hdi00_a_0_),
	.b(regtop_v1_hdi00_a[1]));
   in01f01 U261693 (.o(n249725),
	.a(n245491));
   no02f01 U261695 (.o(n247091),
	.a(n250164),
	.b(regtop_v1_hdi00_a[2]));
   no02f01 U261696 (.o(n246984),
	.a(n246490),
	.b(n246489));
   no02f01 U261697 (.o(n246849),
	.a(n246865),
	.b(n246846));
   no02f08 U261698 (.o(n249211),
	.a(n252542),
	.b(n249106));
   no02f02 U261699 (.o(n245488),
	.a(n245458),
	.b(n245480));
   no02s01 U261700 (.o(n246677),
	.a(n246669),
	.b(n246668));
   na04f01 U261701 (.o(n247014),
	.a(n247013),
	.b(n247012),
	.c(n247011),
	.d(n247010));
   no03f01 U261702 (.o(n246388),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246552),
	.c(n246551));
   no02s01 U261703 (.o(n245887),
	.a(n245841),
	.b(n245856));
   no02s01 U261704 (.o(n245822),
	.a(n245828),
	.b(n245830));
   no02m01 U261705 (.o(n249885),
	.a(n249893),
	.b(n249886));
   in01f01 U261706 (.o(n249771),
	.a(n249542));
   no02f03 U261707 (.o(n247061),
	.a(n247060),
	.b(regtop_v1_hdi00_a[4]));
   no02f06 U261708 (.o(n249210),
	.a(n249111),
	.b(n249110));
   in01f02 U261710 (.o(n246909),
	.a(regtop_g_seqstrt_r));
   no02f01 U261711 (.o(n247059),
	.a(regtop_v1_hdi00_a[5]),
	.b(regtop_v1_hdi00_a[4]));
   no02f02 U261712 (.o(n250201),
	.a(regtop_v1_hdi00_a[0]),
	.b(regtop_v1_hdi00_a[1]));
   in01f01 U261713 (.o(n249948),
	.a(regtop_v1_hdi00_a[2]));
   no03f10 U261714 (.o(n252874),
	.a(regtop_g_a_r[6]),
	.b(FE_OFN491_regtop_g_a_r_3_),
	.c(n245457));
   in01f03 U261715 (.o(n245457),
	.a(n245459));
   na02f02 U261716 (.o(n246865),
	.a(n246902),
	.b(n245516));
   na02f06 U261717 (.o(n245470),
	.a(n245594),
	.b(n245449));
   na02s01 U261718 (.o(n246540),
	.a(n246532),
	.b(n246531));
   na02f01 U261719 (.o(n246968),
	.a(n246967),
	.b(n247007));
   na02f03 U261720 (.o(n245491),
	.a(FE_OFN490_regtop_g_a_r_3_),
	.b(FE_OFN534_regtop_g_a_r_5_));
   na02s01 U261721 (.o(n246504),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246503));
   na03f01 U261722 (.o(n246668),
	.a(n246667),
	.b(n246666),
	.c(n246665));
   na02f01 U261723 (.o(n249893),
	.a(n249902),
	.b(vh_1_ph_add[3]));
   ao12f02 U261724 (.o(n246988),
	.a(n246307),
	.b(n246309),
	.c(n246308));
   ao22s01 U261725 (.o(n246611),
	.a(n252462),
	.b(n252404),
	.c(n246608),
	.d(n246607));
   na02s01 U261726 (.o(n245827),
	.a(vh_1_ph_add[2]),
	.b(vh_1_ph_add[28]));
   no02f01 U261727 (.o(n252831),
	.a(regtop_g_a_r[6]),
	.b(n245445));
   no02f02 U261728 (.o(n249542),
	.a(n245497),
	.b(regtop_g_a_r[6]));
   na02s01 U261729 (.o(n247011),
	.a(n246461),
	.b(n246299));
   na02f01 U261730 (.o(n246307),
	.a(n246306),
	.b(n246305));
   no02f02 U261731 (.o(n247007),
	.a(n246427),
	.b(n246426));
   no02f02 U261732 (.o(n247013),
	.a(n246296),
	.b(n246295));
   in01f02 U261733 (.o(n252542),
	.a(n252684));
   no03f04 U261734 (.o(n245449),
	.a(regtop_g_a_r[8]),
	.b(FE_OFN510_regtop_g_a_r_7_),
	.c(FE_OFN520_regtop_g_a_r_6_));
   na02m01 U261735 (.o(n247012),
	.a(n246480),
	.b(n246324));
   na02s01 U261736 (.o(n245936),
	.a(n245935),
	.b(n245934));
   no02f01 U261737 (.o(n246350),
	.a(n246343),
	.b(n246342));
   na04f02 U261738 (.o(n247010),
	.a(n246670),
	.b(n246335),
	.c(n246334),
	.d(n246333));
   no03s01 U261739 (.o(n246308),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246303),
	.c(n246302));
   no02s01 U261740 (.o(n245410),
	.a(n245408),
	.b(n245407));
   na04f01 U261741 (.o(n246349),
	.a(n246348),
	.b(vldtop_vld_syndec_ADP[4]),
	.c(n246347),
	.d(n246346));
   in01f01 U261742 (.o(n252613),
	.a(n246943));
   no04f01 U261743 (.o(n245937),
	.a(n246402),
	.b(n246403),
	.c(n246670),
	.d(n246401));
   no02f01 U261744 (.o(n246967),
	.a(n246455),
	.b(n246454));
   na03s01 U261745 (.o(n246481),
	.a(n246480),
	.b(n246479),
	.c(n246478));
   no02m02 U261746 (.o(n246441),
	.a(n246440),
	.b(n246439));
   no02s01 U261747 (.o(n245427),
	.a(g_field_start_add_r[28]),
	.b(busrtop_b_rreq_vrh_rrq_fldstatadd_r[28]));
   no02f04 U261748 (.o(n252731),
	.a(regtop_g_paramadr_r[1]),
	.b(n246607));
   no02f03 U261749 (.o(n252568),
	.a(regtop_g_paramadr_r[6]),
	.b(n252575));
   no02f02 U261750 (.o(n245447),
	.a(regtop_g_a_r[2]),
	.b(FE_OFN504_regtop_g_a_r_4_));
   na02f03 U261751 (.o(n249698),
	.a(FE_OFN490_regtop_g_a_r_3_),
	.b(regtop_g_a_r[5]));
   na02f04 U261752 (.o(n245650),
	.a(n245393),
	.b(n245392));
   na02f01 U261753 (.o(n245775),
	.a(n246187),
	.b(n245765));
   na02f02 U261754 (.o(n246060),
	.a(n245774),
	.b(n249107));
   no02f01 U261755 (.o(n246022),
	.a(n246021),
	.b(n246020));
   na02f01 U261756 (.o(n246198),
	.a(n246197),
	.b(n246196));
   no02f03 U261757 (.o(n245459),
	.a(n245452),
	.b(n245458));
   in01m01 U261758 (.o(n245445),
	.a(n245451));
   na02s01 U261759 (.o(n246426),
	.a(n246425),
	.b(n246424));
   no02s01 U261760 (.o(n245397),
	.a(n245399),
	.b(n245398));
   na02f02 U261761 (.o(n245480),
	.a(regtop_g_a_r[2]),
	.b(FE_OFN505_regtop_g_a_r_4_));
   no02s01 U261762 (.o(n245402),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[25]),
	.b(n245406));
   ao12f01 U261763 (.o(n246366),
	.a(n246364),
	.b(n246803),
	.c(vldtop_vld_syndec_ADP[1]));
   na02f02 U261764 (.o(n246826),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246808));
   oa22f01 U261765 (.o(n246802),
	.a(v_vldstatus_r[4]),
	.b(n246801),
	.c(n246800),
	.d(n246799));
   no02m02 U261768 (.o(n246794),
	.a(vldtop_vld_syndec_ADP[2]),
	.b(n246806));
   na02f02 U261769 (.o(n246712),
	.a(n246009),
	.b(n246008));
   na02f01 U261770 (.o(n249107),
	.a(n249108),
	.b(n245773));
   na02m01 U261771 (.o(n245765),
	.a(n246194),
	.b(n245764));
   na02f01 U261772 (.o(n246188),
	.a(n246187),
	.b(n246186));
   no02f01 U261773 (.o(n246453),
	.a(n246452),
	.b(n246451));
   no02f06 U261774 (.o(n245393),
	.a(n245390),
	.b(n245389));
   no03s01 U261775 (.o(n246196),
	.a(n252576),
	.b(n246195),
	.c(n252575));
   no02s01 U261776 (.o(n245398),
	.a(n245396),
	.b(n245395));
   na02m02 U261777 (.o(n245458),
	.a(FE_OFN534_regtop_g_a_r_5_),
	.b(n245451));
   no02f02 U261778 (.o(n246197),
	.a(regtop_g_paramadr_r[5]),
	.b(n246614));
   ao12f02 U261779 (.o(n245774),
	.a(n248996),
	.b(n249108),
	.c(n249109));
   in01f01 U261780 (.o(n252379),
	.a(regtop_g_paramadr_r[6]));
   na02m01 U261781 (.o(n245764),
	.a(n252254),
	.b(n252575));
   no02s01 U261782 (.o(n245385),
	.a(n245387),
	.b(n245386));
   na02f01 U261783 (.o(n246614),
	.a(n246902),
	.b(n246845));
   no02f03 U261784 (.o(n248996),
	.a(n245771),
	.b(n245770));
   na02s01 U261785 (.o(n246797),
	.a(n246882),
	.b(n246796));
   no02f01 U261786 (.o(n245451),
	.a(regtop_g_a_r[7]),
	.b(regtop_g_a_r[8]));
   no02m02 U261787 (.o(n245376),
	.a(n245677),
	.b(n245678));
   no02s01 U261788 (.o(n245381),
	.a(n245378),
	.b(n245377));
   na02s01 U261789 (.o(n246192),
	.a(n248953),
	.b(n246191));
   no02f04 U261790 (.o(n252462),
	.a(regtop_g_paramadr_r[0]),
	.b(regtop_g_paramadr_r[1]));
   no02f03 U261791 (.o(n248953),
	.a(regtop_g_adb_r[0]),
	.b(regtop_g_adb_r[1]));
   in01f01 U261792 (.o(n246607),
	.a(regtop_g_paramadr_r[0]));
   in01f02 U261793 (.o(n249027),
	.a(v_seqstrt_r));
   no02f03 U261794 (.o(n249137),
	.a(n246165),
	.b(n246164));
   na02m02 U261795 (.o(n245544),
	.a(regtop_g_paramadr_r[3]),
	.b(n252380));
   na02m02 U261796 (.o(n245762),
	.a(regtop_g_paramadr_r[2]),
	.b(n252515));
   no02f04 U261797 (.o(n246565),
	.a(vldtop_vld_syndec_ADP[2]),
	.b(n246743));
   no02f01 U261798 (.o(n246171),
	.a(regtop_g_udb2_r[0]),
	.b(n246170));
   na02m02 U261799 (.o(n252449),
	.a(regtop_g_paramadr_r[4]),
	.b(n246608));
   in01f01 U261800 (.o(n246156),
	.a(n246109));
   no02f01 U261801 (.o(n245349),
	.a(n245344),
	.b(n245343));
   no02f01 U261802 (.o(n245352),
	.a(n245340),
	.b(n245339));
   in01f02 U261803 (.o(n252515),
	.a(regtop_g_paramadr_r[4]));
   no02f01 U261804 (.o(n245328),
	.a(n245326),
	.b(n245325));
   no02s01 U261805 (.o(n246732),
	.a(n246731),
	.b(n246882));
   no02f01 U261806 (.o(n245379),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[20]),
	.b(g_field_start_add_r[20]));
   na02f01 U261807 (.o(n246169),
	.a(n246168),
	.b(n246167));
   no02f01 U261808 (.o(n245343),
	.a(g_field_start_add_r[16]),
	.b(n245342));
   no02f01 U261809 (.o(n245339),
	.a(g_field_start_add_r[17]),
	.b(n245360));
   na02f01 U261810 (.o(n246780),
	.a(n249061),
	.b(vldtop_vld_syndec_vld_vscdet_v_search_1st_r));
   no02m02 U261811 (.o(n245361),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[18]),
	.b(g_field_start_add_r[18]));
   in01f02 U261812 (.o(n246087),
	.a(n246080));
   ao22f01 U261813 (.o(n246786),
	.a(vldtop_vld_syndec_vld_vscdet_v_prezerohld_r[0]),
	.b(v1_bs_req_n),
	.c(vldtop_vld_syndec_vld_vscdet_v_prezerotmp_r[0]),
	.d(n246237));
   in01m01 U261814 (.o(n246731),
	.a(v_vldstatus_r[4]));
   no02f02 U261815 (.o(n249007),
	.a(vldtop_vld_syndec_UREG[16]),
	.b(n246914));
   no02f02 U261816 (.o(n246166),
	.a(regtop_g_udb1_r[0]),
	.b(regtop_g_udb0_r[0]));
   no02f02 U261817 (.o(n246065),
	.a(n246066),
	.b(regtop_g_udb2_r[1]));
   in01f03 U261818 (.o(n246743),
	.a(vldtop_vld_syndec_ADP[3]));
   no02f02 U261819 (.o(n246659),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(vldtop_vld_syndec_ADP[3]));
   ao22f01 U261820 (.o(n246130),
	.a(regtop_g_udb0_r[6]),
	.b(regtop_g_udb2_r[6]),
	.c(n246128),
	.d(n246924));
   no02f01 U261821 (.o(n246361),
	.a(v_vldstatus_r[0]),
	.b(v_vldstatus_r[1]));
   na02f03 U261822 (.o(n246684),
	.a(n246419),
	.b(n246692));
   in01f01 U261823 (.o(n246359),
	.a(vldtop_vld_syndec_UREG[8]));
   na02f02 U261824 (.o(n246112),
	.a(regtop_g_udb2_r[4]),
	.b(n246095));
   in01f02 U261825 (.o(n246692),
	.a(vldtop_vld_syndec_ADP[2]));
   no03f02 U261826 (.o(n246354),
	.a(vldtop_vld_syndec_UREG[9]),
	.b(vldtop_vld_syndec_UREG[10]),
	.c(vldtop_vld_syndec_UREG[13]));
   in01f10 U261827 (.o(n246419),
	.a(vldtop_vld_syndec_ADP[1]));
   no04f02 U261828 (.o(n246355),
	.a(vldtop_vld_syndec_UREG[28]),
	.b(vldtop_vld_syndec_UREG[26]),
	.c(vldtop_vld_syndec_UREG[29]),
	.d(vldtop_vld_syndec_UREG[30]));
   no03f02 U261829 (.o(n246356),
	.a(vldtop_vld_syndec_UREG[27]),
	.b(vldtop_vld_syndec_UREG[25]),
	.c(vldtop_vld_syndec_UREG[31]));
   no04f02 U261830 (.o(n246353),
	.a(vldtop_vld_syndec_UREG[11]),
	.b(vldtop_vld_syndec_UREG[14]),
	.c(vldtop_vld_syndec_UREG[12]),
	.d(vldtop_vld_syndec_UREG[15]));
   na02f02 U261831 (.o(n246123),
	.a(regtop_g_udb0_r[5]),
	.b(regtop_g_udb1_r[5]));
   na02f04 U261832 (.o(n246069),
	.a(regtop_g_udb1_r[2]),
	.b(n246076));
   na02f01 U261833 (.o(n246144),
	.a(n246122),
	.b(n246121));
   na02f02 U261834 (.o(n246484),
	.a(n246570),
	.b(vldtop_vld_syndec_ADP[4]));
   no02f01 U261835 (.o(n249947),
	.a(regtop_v1_hdi00_bs),
	.b(regtop_v1_hdi00_we));
   na02f02 U261836 (.o(n248990),
	.a(n246158),
	.b(n246157));
   no02m02 U261837 (.o(n245517),
	.a(regtop_g_paramadr_r[4]),
	.b(regtop_g_paramadr_r[2]));
   na02s01 U261838 (.o(n246444),
	.a(n246565),
	.b(n246345));
   no02s01 U261839 (.o(n246460),
	.a(n246459),
	.b(n246458));
   no02s01 U261840 (.o(n246447),
	.a(n246446),
	.b(n246445));
   na02s01 U261841 (.o(n246363),
	.a(vldtop_vld_syndec_vld_seqhed_pre_SHIFT[1]),
	.b(n249027));
   na02f04 U261842 (.o(n249697),
	.a(n245447),
	.b(n245449));
   na02m02 U261843 (.o(n246200),
	.a(regtop_g_a_r[8]),
	.b(FE_OFN550_n249113));
   no02f03 U261844 (.o(n249108),
	.a(n252382),
	.b(n245763));
   na02f01 U261845 (.o(n246103),
	.a(n246100),
	.b(n246106));
   no02f01 U261846 (.o(n246164),
	.a(n246163),
	.b(n246162));
   na02s01 U261847 (.o(n245973),
	.a(n246706),
	.b(n245972));
   no02f01 U261848 (.o(n246438),
	.a(n246437),
	.b(n246436));
   in01f03 U261849 (.o(n246700),
	.a(n246527));
   na02f04 U261850 (.o(n246711),
	.a(n246565),
	.b(n246670));
   na02s01 U261851 (.o(n246462),
	.a(n246461),
	.b(n246460));
   na02s01 U261852 (.o(n246449),
	.a(n246448),
	.b(n246447));
   na02f03 U261853 (.o(n246795),
	.a(n246662),
	.b(n246659));
   no02s01 U261854 (.o(n245433),
	.a(g_field_start_add_r[29]),
	.b(busrtop_b_rreq_vrh_rrq_fldstatadd_r[29]));
   no02s01 U261855 (.o(n245401),
	.a(g_field_start_add_r[25]),
	.b(n245406));
   no02f01 U261856 (.o(n245340),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[17]),
	.b(n245360));
   na02s01 U261857 (.o(n245853),
	.a(vh_1_ph_add[4]),
	.b(vh_1_ph_add[30]));
   no02s01 U261858 (.o(n245841),
	.a(vh_1_ph_add[4]),
	.b(vh_1_ph_add[30]));
   no02f02 U261859 (.o(n249731),
	.a(n245444),
	.b(n249627));
   no02f03 U261860 (.o(n250055),
	.a(n249948),
	.b(FE_OFN497_n249947));
   na02s01 U261861 (.o(n246846),
	.a(n252379),
	.b(n246845));
   no03f01 U261862 (.o(n245766),
	.a(n245547),
	.b(n245579),
	.c(n245939));
   no03s01 U261863 (.o(n246324),
	.a(n246477),
	.b(n246476),
	.c(n246670));
   no02f02 U261864 (.o(n246528),
	.a(n246031),
	.b(n246030));
   na04f02 U261865 (.o(n246721),
	.a(n246720),
	.b(n246719),
	.c(n246718),
	.d(n246717));
   no04f02 U261866 (.o(n246520),
	.a(n246510),
	.b(n246671),
	.c(n246509),
	.d(n246508));
   na02s01 U261867 (.o(n246489),
	.a(n246488),
	.b(n246487));
   na02f02 U261868 (.o(n245481),
	.a(n252831),
	.b(n245479));
   no04f04 U261869 (.o(n246787),
	.a(n246786),
	.b(n249005),
	.c(n246785),
	.d(n246784));
   na02f01 U261870 (.o(n245497),
	.a(FE_OFN491_regtop_g_a_r_3_),
	.b(n245459));
   no02f01 U261871 (.o(n248408),
	.a(n247109),
	.b(FE_OFN28_n251337));
   no02f06 U261875 (.o(n245405),
	.a(n245402),
	.b(n245401));
   no02f01 U261876 (.o(n249855),
	.a(n249863),
	.b(n249856));
   na02s01 U261877 (.o(n246234),
	.a(busiftop_status_b_current_0_),
	.b(n246233));
   no04f02 U261878 (.o(n245590),
	.a(n245575),
	.b(n245574),
	.c(n245573),
	.d(n252368));
   no04f04 U261879 (.o(n245591),
	.a(n252376),
	.b(n252374),
	.c(n252372),
	.d(n245536));
   no02s02 U261880 (.o(n245505),
	.a(n245504),
	.b(n245503));
   na02f01 U261881 (.o(n249930),
	.a(n249929),
	.b(FE_OFN439_n252264));
   na03f03 U261882 (.o(n249388),
	.a(n245479),
	.b(n245492),
	.c(n245490));
   na02f03 U261883 (.o(n249829),
	.a(FE_OFN4_n245443),
	.b(FE_OFN398_n249646));
   na03f01 U261884 (.o(n250202),
	.a(regtop_v1_hdi00_a[5]),
	.b(regtop_v1_hdi00_a[3]),
	.c(regtop_v1_hdi00_a[4]));
   na02f04 U261885 (.o(n251977),
	.a(n250055),
	.b(n250128));
   na02s01 U261886 (.o(n252274),
	.a(n247595),
	.b(n247594));
   no02f02 U261887 (.o(n245761),
	.a(n252515),
	.b(n246845));
   no02f01 U261888 (.o(n252700),
	.a(n252449),
	.b(n252448));
   no02s01 U261889 (.o(n246612),
	.a(n246611),
	.b(n246610));
   no02f03 U261890 (.o(n248952),
	.a(n249137),
	.b(n249135));
   no02s01 U261891 (.o(n246581),
	.a(n246580),
	.b(n246579));
   na02f01 U261892 (.o(n245560),
	.a(n252379),
	.b(regtop_g_nferror_r));
   na02f03 U261893 (.o(n246799),
	.a(n249061),
	.b(n249011));
   no02f06 U261894 (.o(n246365),
	.a(n246366),
	.b(n246419));
   in01f01 U261895 (.o(n247149),
	.a(n247143));
   in01m01 U261896 (.o(n247144),
	.a(n246853));
   na02f02 U261897 (.o(n249789),
	.a(n245479),
	.b(n252867));
   na02f01 U261898 (.o(n245605),
	.a(n245429),
	.b(n245428));
   na02s01 U261899 (.o(n245642),
	.a(n245399),
	.b(n245398));
   no02f01 U261900 (.o(n245666),
	.a(n245712),
	.b(n245710));
   na04f02 U261901 (.o(n249520),
	.a(n249519),
	.b(n249518),
	.c(n249517),
	.d(n249516));
   na04f02 U261902 (.o(n249503),
	.a(n249502),
	.b(n249501),
	.c(n249500),
	.d(n249499));
   na04s01 U261903 (.o(n249504),
	.a(n249498),
	.b(n249497),
	.c(n249496),
	.d(n249495));
   na03f01 U261904 (.o(n249749),
	.a(n249748),
	.b(n249747),
	.c(n249685));
   na04f01 U261905 (.o(n249538),
	.a(n249532),
	.b(n249531),
	.c(n249530),
	.d(n249529));
   na04f04 U261906 (.o(n249406),
	.a(n249400),
	.b(n249399),
	.c(n249398),
	.d(n249397));
   na03f01 U261907 (.o(n249392),
	.a(FE_OFN445_n249391),
	.b(n249390),
	.c(n249389));
   in01f06 U261909 (.o(n250272),
	.a(FE_OFN278_n250254));
   no02f03 U261912 (.o(n250682),
	.a(n252086),
	.b(FE_OFN556_n250770));
   in01f08 U261913 (.o(n250804),
	.a(FE_OFN296_n250789));
   no02f01 U261916 (.o(n251211),
	.a(n252050),
	.b(FE_OFN28_n251337));
   in01f06 U261917 (.o(n251335),
	.a(FE_OFN316_n251317));
   no02f02 U261920 (.o(n251746),
	.a(n252013),
	.b(FE_OFN32_n251904));
   in01f08 U261921 (.o(n251867),
	.a(FE_OFN561_n251852));
   no02f08 U261924 (.o(n249252),
	.a(n249250),
	.b(n252811));
   na04f03 U261925 (.o(n246204),
	.a(regtop_g_a_r[8]),
	.b(n249725),
	.c(n245492),
	.d(FE_OFN520_regtop_g_a_r_6_));
   no02f02 U261926 (.o(n245492),
	.a(regtop_g_a_r[2]),
	.b(regtop_g_a_r[4]));
   na02f03 U261927 (.o(n246922),
	.a(n252462),
	.b(n246908));
   na02f01 U261928 (.o(n246877),
	.a(n246870),
	.b(n246874));
   na02f06 U261929 (.o(n252446),
	.a(n252775),
	.b(n252425));
   na02f03 U261930 (.o(n246930),
	.a(n252523),
	.b(n246908));
   no02f01 U261931 (.o(n252642),
	.a(regtop_g_paramadr_r[6]),
	.b(n246943));
   na02f02 U261932 (.o(n247018),
	.a(n246562),
	.b(n246561));
   na03m02 U261933 (.o(n247192),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247191));
   na04f03 U261934 (.o(n248821),
	.a(n248815),
	.b(n248814),
	.c(n248813),
	.d(n248812));
   na04f06 U261935 (.o(n248146),
	.a(n248145),
	.b(n248144),
	.c(n248143),
	.d(n248142));
   na04f01 U261936 (.o(n247540),
	.a(n247522),
	.b(n247521),
	.c(n247520),
	.d(n247519));
   na04f04 U261937 (.o(n247437),
	.a(n247425),
	.b(n247424),
	.c(n247423),
	.d(n247422));
   na04f06 U261938 (.o(n247861),
	.a(n247855),
	.b(n247854),
	.c(n247853),
	.d(n247852));
   na04f04 U261939 (.o(n248946),
	.a(n248945),
	.b(n248944),
	.c(n248943),
	.d(n248942));
   na04f01 U261940 (.o(n248487),
	.a(n248471),
	.b(n248470),
	.c(n248469),
	.d(n248468));
   na04f04 U261941 (.o(n247648),
	.a(n247624),
	.b(n247623),
	.c(n247622),
	.d(n247621));
   na04f04 U261942 (.o(n247757),
	.a(n247751),
	.b(n247750),
	.c(n247749),
	.d(n247748));
   na04f06 U261943 (.o(n247882),
	.a(n247881),
	.b(n247880),
	.c(n247879),
	.d(n247878));
   na04f02 U261944 (.o(n248465),
	.a(n248449),
	.b(n248448),
	.c(n248447),
	.d(n248446));
   na04f02 U261945 (.o(n248114),
	.a(n248103),
	.b(n248102),
	.c(n248101),
	.d(n248100));
   na04f03 U261946 (.o(n248757),
	.a(n248751),
	.b(n248750),
	.c(n248749),
	.d(n248748));
   na04f02 U261947 (.o(n248798),
	.a(n248797),
	.b(n248796),
	.c(n248795),
	.d(n248794));
   na04f01 U261948 (.o(n248655),
	.a(n248639),
	.b(n248638),
	.c(n248637),
	.d(n248636));
   na04f03 U261949 (.o(n248528),
	.a(n248517),
	.b(n248516),
	.c(n248515),
	.d(n248514));
   na04f04 U261950 (.o(n248611),
	.a(n248605),
	.b(n248604),
	.c(n248603),
	.d(n248602));
   no02s01 U261951 (.o(n245671),
	.a(n245670),
	.b(n245672));
   no03s01 U261952 (.o(n249524),
	.a(n249522),
	.b(n249521),
	.c(n249520));
   no03s01 U261953 (.o(n249507),
	.a(n249505),
	.b(n249504),
	.c(n249503));
   no04f03 U261954 (.o(n249604),
	.a(n249603),
	.b(n249602),
	.c(n249601),
	.d(n249600));
   in01f08 U261955 (.o(n245444),
	.a(FE_OFN4_n245443));
   no03f03 U261956 (.o(n249832),
	.a(n249664),
	.b(FE_OFN449_n249831),
	.c(n249830));
   no02f01 U261957 (.o(n249808),
	.a(n249806),
	.b(n249805));
   no02s01 U261958 (.o(n249408),
	.a(n249406),
	.b(n249405));
   no02f01 U261959 (.o(n248989),
	.a(regtop_N1990),
	.b(n245026));
   no02f01 U261961 (.o(n249169),
	.a(n249167),
	.b(n249166));
   na02f01 U261962 (.o(n249253),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[12]));
   na02f01 U261963 (.o(n249083),
	.a(regtop_g_paramdata_r[23]),
	.b(n249132));
   na02f01 U261964 (.o(n248956),
	.a(regtop_g_paramdata_r[20]),
	.b(n248980));
   na02s01 U261965 (.o(n249119),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[16]));
   na02f03 U261966 (.o(n252273),
	.a(n247595),
	.b(n249663));
   na02f01 U261967 (.o(n252829),
	.a(n253015),
	.b(n249725));
   na02f02 U261968 (.o(n247034),
	.a(n246909),
	.b(n246922));
   na02f08 U261969 (.o(n252401),
	.a(FE_OFN39_n252462),
	.b(n252730));
   na02f01 U261970 (.o(n252422),
	.a(FE_OFN39_n252462),
	.b(n252711));
   na02f02 U261971 (.o(n247045),
	.a(n246909),
	.b(n246930));
   na02f01 U261972 (.o(n252508),
	.a(n252523),
	.b(n252711));
   na02f02 U261973 (.o(n252676),
	.a(n245763),
	.b(n245525));
   na02f02 U261974 (.o(n252709),
	.a(n252731),
	.b(n252706));
   na02f03 U261975 (.o(n252780),
	.a(n252776),
	.b(n252775));
   no02f02 U261976 (.o(n246890),
	.a(n245937),
	.b(n245936));
   na03f02 U261977 (.o(n252816),
	.a(n252238),
	.b(regtop_g_ferror_r),
	.c(n252379));
   no02f02 U261978 (.o(n252818),
	.a(FE_OFN439_n252264),
	.b(n252894));
   no04s02 U261979 (.o(n249026),
	.a(n249020),
	.b(n249019),
	.c(n249018),
	.d(n249017));
   in01f06 U261981 (.o(n252834),
	.a(FE_OFN454_n252863));
   na02f01 U261982 (.o(n247146),
	.a(y1_bs_wait_n),
	.b(vldtop_vld_syndec_vld_vlfeed_feed_on));
   na02f01 U261983 (.o(n252905),
	.a(FE_OFN499_n253015),
	.b(n252874));
   na02f04 U261985 (.o(n253012),
	.a(n253015),
	.b(n252998));
   na02f04 U261986 (.o(n253029),
	.a(n253015),
	.b(n253014));
   no04f04 U261987 (.o(n248186),
	.a(n248149),
	.b(n248148),
	.c(n248147),
	.d(n248146));
   no04f06 U261988 (.o(n248950),
	.a(n248949),
	.b(n248948),
	.c(n248947),
	.d(n248946));
   no04f01 U261989 (.o(n247907),
	.a(n247885),
	.b(n247884),
	.c(n247883),
	.d(n247882));
   no04f06 U261990 (.o(n248802),
	.a(n248801),
	.b(n248800),
	.c(FE_OFN252_n248799),
	.d(n248798));
   na03s01 U261991 (.o(n157834),
	.a(n249877),
	.b(n249876),
	.c(n249875));
   na04f04 U261992 (.o(n244218),
	.a(n245486),
	.b(n245485),
	.c(n245484),
	.d(n245483));
   na04f02 U261993 (.o(n244977),
	.a(n249456),
	.b(n249455),
	.c(n249454),
	.d(n249453));
   na04f02 U261994 (.o(n244985),
	.a(n249366),
	.b(n249365),
	.c(n249364),
	.d(n249363));
   na02m02 U261995 (.o(n245026),
	.a(n246206),
	.b(FE_OFN503_n246205));
   na02f02 U261996 (.o(n244994),
	.a(n249195),
	.b(n249194));
   na02f04 U261997 (.o(n245008),
	.a(n249226),
	.b(n249225));
   na03f02 U261998 (.o(n245025),
	.a(n248961),
	.b(n248960),
	.c(n248959));
   no02f01 U261999 (.o(n211948),
	.a(regtop_g_seqstrt_r),
	.b(n246926));
   no02s01 U262000 (.o(n212049),
	.a(regtop_g_seqstrt_r),
	.b(n246934));
   na02s01 U262001 (.o(n212286),
	.a(n246748),
	.b(n246747));
   na02f01 U262002 (.o(n212425),
	.a(n247254),
	.b(n247138));
   na02f01 U262003 (.o(n212594),
	.a(n247154),
	.b(n247153));
   na02f01 U262004 (.o(n212608),
	.a(n247209),
	.b(n247208));
   na02f01 U262005 (.o(n212624),
	.a(n247307),
	.b(n247306));
   no02f01 U262006 (.o(n253047),
	.a(n247359),
	.b(n247358));
   no02f01 U262007 (.o(n253062),
	.a(n247458),
	.b(n247457));
   na02f10 U262008 (.o(n247126),
	.a(n247125),
	.b(n247143));
   oa22f04 U262011 (.o(n248980),
	.a(n248955),
	.b(n249250),
	.c(n248954),
	.d(n249081));
   no02f08 U262012 (.o(n247494),
	.a(n247143),
	.b(n247144));
   na02f08 U262013 (.o(n247143),
	.a(n246822),
	.b(n246821));
   no02f02 U262015 (.o(n246908),
	.a(n246904),
	.b(n246903));
   na02f02 U262016 (.o(n246819),
	.a(n246818),
	.b(n246365));
   no03m02 U262017 (.o(n246820),
	.a(n246817),
	.b(n246816),
	.c(n246815));
   no02f04 U262018 (.o(n249113),
	.a(n245776),
	.b(n252542));
   no02f04 U262019 (.o(n248978),
	.a(n248952),
	.b(n252813));
   na02f03 U262020 (.o(n246830),
	.a(n246737),
	.b(n246743));
   in01m01 U262021 (.o(n252601),
	.a(n252595));
   ao12f02 U262022 (.o(n246815),
	.a(n246802),
	.b(n246804),
	.c(n246803));
   in01f02 U262023 (.o(n246791),
	.a(n246790));
   in01f04 U262024 (.o(n252995),
	.a(FE_OFN458_n252996));
   na02f06 U262025 (.o(n252460),
	.a(FE_OFN39_n252462),
	.b(FE_OFN45_n252700));
   no02f03 U262026 (.o(n252711),
	.a(n252448),
	.b(n252405));
   in01f06 U262027 (.o(n252339),
	.a(FE_OFN354_n252338));
   in01f02 U262028 (.o(n249041),
	.a(n246198));
   in01f02 U262029 (.o(n252270),
	.a(n252264));
   no02f01 U262030 (.o(n246162),
	.a(n246161),
	.b(n246163));
   no02f08 U262031 (.o(n252871),
	.a(FE_OFN498_n253015),
	.b(n249771));
   in01f04 U262032 (.o(n252941),
	.a(FE_OFN456_n252942));
   no02f04 U262033 (.o(n252969),
	.a(FE_OFN498_n253015),
	.b(n252958));
   in01m01 U262034 (.o(n246685),
	.a(n246803));
   in01f04 U262035 (.o(n252972),
	.a(n249789));
   in01f06 U262036 (.o(n252875),
	.a(FE_OFN441_n252905));
   in01f04 U262037 (.o(n252445),
	.a(FE_OFN37_n252446));
   na03f04 U262038 (.o(n252264),
	.a(n253015),
	.b(n245594),
	.c(n245593));
   na02f02 U262039 (.o(n246121),
	.a(n246120),
	.b(n246119));
   no02f02 U262040 (.o(n246803),
	.a(n246778),
	.b(n246780));
   na02f01 U262041 (.o(n252668),
	.a(n252764),
	.b(n252642));
   in01f02 U262042 (.o(n252697),
	.a(n252698));
   na02f08 U262043 (.o(n252561),
	.a(n252568),
	.b(n252764));
   na02f03 U262044 (.o(n245924),
	.a(n252597),
	.b(FE_OFN218_n246238));
   in01m01 U262045 (.o(n246804),
	.a(n246795));
   in01m01 U262046 (.o(n252867),
	.a(n245487));
   no02f06 U262047 (.o(n249663),
	.a(n246372),
	.b(n245448));
   no02f04 U262048 (.o(n252998),
	.a(n249698),
	.b(n249720));
   no02f08 U262049 (.o(n249825),
	.a(n245444),
	.b(n249388));
   na02f03 U262050 (.o(n252382),
	.a(n246863),
	.b(n245762));
   in01m01 U262051 (.o(n245899),
	.a(n245840));
   na02m01 U262052 (.o(n245627),
	.a(n245411),
	.b(n245410));
   na02f01 U262053 (.o(n245826),
	.a(n245824),
	.b(n245887));
   no02s01 U262054 (.o(n245423),
	.a(n245419),
	.b(n245418));
   in01f02 U262055 (.o(n246662),
	.a(n246684));
   na02f10 U262056 (.o(n252195),
	.a(n247056),
	.b(n247055));
   in01m01 U262058 (.o(n246362),
	.a(n246361));
   in01f01 U262059 (.o(n245514),
	.a(n245517));
   no02f01 U262061 (.o(n246206),
	.a(n249072),
	.b(n249073));
   no02f02 U262062 (.o(n247350),
	.a(n247149),
	.b(n247144));
   in01f01 U262063 (.o(n246941),
	.a(n246880));
   no02f02 U262064 (.o(n246880),
	.a(n246904),
	.b(n246848));
   na02f02 U262065 (.o(n246821),
	.a(n246820),
	.b(n246819));
   no02f02 U262068 (.o(n246818),
	.a(n246794),
	.b(n246793));
   in01f01 U262069 (.o(n246203),
	.a(n246202));
   in01f02 U262070 (.o(n246810),
	.a(n246816));
   no02f02 U262071 (.o(n246202),
	.a(n246201),
	.b(n246200));
   na02f02 U262072 (.o(n246793),
	.a(n246830),
	.b(n246827));
   na03f02 U262073 (.o(n247026),
	.a(n247025),
	.b(n247024),
	.c(n247023));
   in01f02 U262074 (.o(n246827),
	.a(n246809));
   in01f01 U262075 (.o(n246817),
	.a(n246826));
   no03f08 U262076 (.o(n249945),
	.a(n249928),
	.b(n249927),
	.c(n249926));
   no02f03 U262077 (.o(n246647),
	.a(n249082),
	.b(n252813));
   in01f02 U262078 (.o(n246808),
	.a(n246792));
   na02f03 U262079 (.o(n246773),
	.a(n248952),
	.b(FE_OFN6_n246618));
   in01f03 U262080 (.o(n252459),
	.a(n252460));
   in01f03 U262081 (.o(n252421),
	.a(FE_OFN212_n252422));
   in01f04 U262082 (.o(n252400),
	.a(n252401));
   in01f04 U262084 (.o(n252629),
	.a(FE_OFN558_n252630));
   in01f04 U262085 (.o(n252727),
	.a(FE_OFN360_n252728));
   in01f04 U262086 (.o(n252747),
	.a(FE_OFN362_n252748));
   in01f04 U262087 (.o(n252507),
	.a(FE_OFN356_n252508));
   na02f03 U262088 (.o(n246738),
	.a(n246736),
	.b(n249027));
   na02f08 U262089 (.o(n246189),
	.a(n246197),
	.b(n246188));
   no03f03 U262090 (.o(n252595),
	.a(n252576),
	.b(n252575),
	.c(n252574));
   na02s02 U262096 (.o(n252574),
	.a(n246849),
	.b(n246909));
   in01f02 U262102 (.o(n252970),
	.a(n252969));
   no02f02 U262103 (.o(n246806),
	.a(n246685),
	.b(n246662));
   in01f06 U262115 (.o(n252730),
	.a(n252510));
   na02f08 U262122 (.o(n249081),
	.a(n252684),
	.b(n249041));
   in01m01 U262123 (.o(n248985),
	.a(n249107));
   no02f08 U262162 (.o(n249664),
	.a(n245444),
	.b(FE_OFN526_n249548));
   no02f03 U262165 (.o(n247603),
	.a(n249588),
	.b(n252274));
   na02f01 U262167 (.o(n246187),
	.a(n249108),
	.b(n246607));
   no02f01 U262168 (.o(n252863),
	.a(FE_OFN548_regtop_g_a_r_2_),
	.b(n252832));
   in01f02 U262172 (.o(n253028),
	.a(n253029));
   na02f01 U262176 (.o(n246903),
	.a(n246902),
	.b(n246901));
   in01f02 U262177 (.o(n253011),
	.a(n253012));
   in01s01 U262182 (.o(n246800),
	.a(n246798));
   no02f02 U262185 (.o(n249135),
	.a(n246172),
	.b(n246171));
   na02f04 U262187 (.o(n246247),
	.a(n248953),
	.b(FE_OFN218_n246238));
   na02f02 U262195 (.o(n246161),
	.a(n246160),
	.b(n246159));
   in01f04 U262197 (.o(n252482),
	.a(FE_OFN214_n252483));
   na02f06 U262198 (.o(n252773),
	.a(n252776),
	.b(n252764));
   na02f06 U262220 (.o(n252350),
	.a(n252352),
	.b(n252764));
   na02f04 U262222 (.o(n252361),
	.a(n252567),
	.b(n252352));
   na02f02 U262224 (.o(n252954),
	.a(FE_OFN499_n253015),
	.b(n252944));
   no02f04 U262231 (.o(n253014),
	.a(n246372),
	.b(n245487));
   in01f01 U262232 (.o(n252866),
	.a(n252829));
   no02f04 U262233 (.o(n246778),
	.a(n246795),
	.b(n246782));
   no02f03 U262234 (.o(n252944),
	.a(n245448),
	.b(n245491));
   no02f06 U262235 (.o(n252912),
	.a(FE_OFN491_regtop_g_a_r_3_),
	.b(n245477));
   no02f01 U262236 (.o(n246261),
	.a(n252234),
	.b(n246225));
   ao12s01 U262237 (.o(n245879),
	.a(n245877),
	.b(n245878),
	.c(n245899));
   no02f01 U262238 (.o(n246172),
	.a(n246169),
	.b(n246170));
   no02f01 U262239 (.o(n249648),
	.a(FE_OFN509_regtop_g_a_r_7_),
	.b(n246204));
   no02s01 U262241 (.o(n245409),
	.a(n245411),
	.b(n245410));
   no02f02 U262242 (.o(n246863),
	.a(n245848),
	.b(n245761));
   in01m01 U262243 (.o(n252687),
	.a(n252517));
   in01s01 U262244 (.o(n246613),
	.a(n246612));
   in01m01 U262245 (.o(n252314),
	.a(n245848));
   na02f02 U262246 (.o(n249720),
	.a(n245594),
	.b(n245490));
   oa12f06 U262247 (.o(n245942),
	.a(n245825),
	.b(n245826),
	.c(n245840));
   na02f02 U262248 (.o(n246729),
	.a(n246662),
	.b(n246743));
   in01f01 U262249 (.o(n246706),
	.a(n246578));
   na02s01 U262251 (.o(n245612),
	.a(n245423),
	.b(n245422));
   na02f01 U262252 (.o(n245849),
	.a(n245848),
	.b(n252568));
   no02f02 U262253 (.o(n245490),
	.a(n245445),
	.b(FE_OFN520_regtop_g_a_r_6_));
   ao12f02 U262254 (.o(n245840),
	.a(n245821),
	.b(n245823),
	.c(n245822));
   no02s01 U262255 (.o(n245429),
	.a(n245426),
	.b(n245425));
   no02f02 U262256 (.o(n245848),
	.a(n245514),
	.b(n245518));
   na02f02 U262257 (.o(n245825),
	.a(n245824),
	.b(n245886));
   no02f02 U262258 (.o(n249061),
	.a(n246731),
	.b(n246362));
   na02s01 U262259 (.o(n252685),
	.a(n252684),
	.b(n252731));
   in01f03 U262260 (.o(n246570),
	.a(n246693));
   na02f04 U262261 (.o(n249005),
	.a(n246358),
	.b(n246357));
   no02s01 U262262 (.o(n247147),
	.a(n247146),
	.b(n247145));
   no02f02 U262263 (.o(n245594),
	.a(FE_OFN549_regtop_g_a_r_2_),
	.b(FE_OFN506_regtop_g_a_r_4_));
   na02s01 U262264 (.o(n252463),
	.a(n252684),
	.b(n252462));
   no02f01 U262265 (.o(n245824),
	.a(n245895),
	.b(n245820));
   na02f02 U262266 (.o(n245528),
	.a(n245527),
	.b(n252515));
   in01s01 U262267 (.o(n252384),
	.a(n252383));
   in01s01 U262268 (.o(n247478),
	.a(n247476));
   in01s01 U262269 (.o(n247194),
	.a(n247192));
   in01s01 U262270 (.o(n247327),
	.a(n247325));
   in01f01 U262271 (.o(n247496),
	.a(n247493));
   in01f01 U262272 (.o(n247474),
	.a(n247472));
   in01f01 U262273 (.o(n247359),
	.a(n247357));
   no02f01 U262274 (.o(n247334),
	.a(FE_OCPN583_n247126),
	.b(n247333));
   no02f01 U262275 (.o(n247216),
	.a(n247126),
	.b(n247215));
   no02f01 U262276 (.o(n247224),
	.a(FE_OCPN583_n247126),
	.b(n247223));
   no02f02 U262277 (.o(n247260),
	.a(FE_OFN577_n247126),
	.b(n247259));
   no02s01 U262278 (.o(n247165),
	.a(FE_OCPN583_n247126),
	.b(n247164));
   no02f01 U262279 (.o(n247201),
	.a(FE_OFN577_n247126),
	.b(n247200));
   no02f01 U262280 (.o(n247129),
	.a(FE_OFN577_n247126),
	.b(n247128));
   no02f01 U262281 (.o(n247175),
	.a(FE_OCPN583_n247126),
	.b(n247174));
   no02f01 U262282 (.o(n247185),
	.a(FE_OCPN583_n247126),
	.b(n247184));
   no02f01 U262283 (.o(n247197),
	.a(FE_OCPN583_n247126),
	.b(n247196));
   no02s01 U262284 (.o(n247230),
	.a(FE_OFN577_n247126),
	.b(n247229));
   no02f01 U262285 (.o(n247266),
	.a(FE_OCPN583_n247126),
	.b(n247265));
   no02f01 U262286 (.o(n247181),
	.a(n247126),
	.b(n247180));
   no02f02 U262287 (.o(n247141),
	.a(n247126),
	.b(n247140));
   no02f01 U262288 (.o(n247161),
	.a(n247126),
	.b(n247160));
   no02f01 U262289 (.o(n247212),
	.a(n247126),
	.b(n247211));
   no02f02 U262290 (.o(n247310),
	.a(FE_OFN577_n247126),
	.b(n247309));
   no02f01 U262291 (.o(n247314),
	.a(FE_OFN577_n247126),
	.b(n247313));
   no02s01 U262292 (.o(n247291),
	.a(n247126),
	.b(n247290));
   no02f01 U262293 (.o(n247318),
	.a(FE_OCPN583_n247126),
	.b(n247317));
   no02f01 U262294 (.o(n247278),
	.a(FE_OCPN583_n247126),
	.b(n247277));
   no02f01 U262295 (.o(n247295),
	.a(FE_OFN577_n247126),
	.b(n247294));
   no02f02 U262296 (.o(n247366),
	.a(FE_OFN577_n247126),
	.b(n247365));
   no02f01 U262297 (.o(n247370),
	.a(FE_OCPN583_n247126),
	.b(n247369));
   no02f01 U262298 (.o(n247274),
	.a(FE_OCPN583_n247126),
	.b(n247273));
   no02f02 U262299 (.o(n247171),
	.a(FE_OFN577_n247126),
	.b(n247170));
   no02f01 U262300 (.o(n247133),
	.a(FE_OFN577_n247126),
	.b(n247132));
   no02f01 U262301 (.o(n247157),
	.a(FE_OCPN583_n247126),
	.b(n247156));
   no02f01 U262302 (.o(n247242),
	.a(n247126),
	.b(n247241));
   no02f10 U262307 (.o(n249189),
	.a(n249252),
	.b(FE_OFN551_n249140));
   in01f01 U262308 (.o(n247441),
	.a(FE_OFN18_n247494));
   no02f02 U262309 (.o(n247150),
	.a(n247149),
	.b(n247148));
   oa22f04 U262310 (.o(n249132),
	.a(n249250),
	.b(n249082),
	.c(n249081),
	.d(n249080));
   in01f02 U262311 (.o(n248992),
	.a(n248993));
   na02f04 U262312 (.o(n249073),
	.a(n249250),
	.b(n249081));
   no03f02 U262313 (.o(n246925),
	.a(n246922),
	.b(n247039),
	.c(n246921));
   oa12f02 U262314 (.o(n246870),
	.a(n246909),
	.b(n246904),
	.c(n246850));
   in01f02 U262315 (.o(n246822),
	.a(n246814));
   na02f02 U262316 (.o(n247254),
	.a(n247137),
	.b(n249255));
   na02f02 U262317 (.o(n246814),
	.a(n246813),
	.b(n246812));
   no02f08 U262318 (.o(n246904),
	.a(n249029),
	.b(n246185));
   na02f06 U262319 (.o(n246185),
	.a(n249042),
	.b(n246184));
   na03f02 U262320 (.o(n246813),
	.a(n246818),
	.b(n246815),
	.c(n246365));
   oa12f02 U262321 (.o(n246812),
	.a(n246815),
	.b(n246806),
	.c(n246811));
   na02s01 U262322 (.o(n245626),
	.a(n245622),
	.b(n245623));
   no02s01 U262323 (.o(n245633),
	.a(n245629),
	.b(n245630));
   na02m02 U262324 (.o(n246811),
	.a(n246826),
	.b(n246810));
   na03f02 U262326 (.o(n247030),
	.a(n247028),
	.b(n247027),
	.c(n247026));
   no02s01 U262327 (.o(n245630),
	.a(n245629),
	.b(n245631));
   no02f02 U262328 (.o(n246816),
	.a(n246809),
	.b(n246828));
   no02f04 U262329 (.o(n249029),
	.a(n246105),
	.b(n246104));
   no02f02 U262330 (.o(n247008),
	.a(n246996),
	.b(n246995));
   na03s02 U262331 (.o(n246995),
	.a(n246994),
	.b(n246993),
	.c(n246992));
   no02m02 U262332 (.o(n246104),
	.a(n246103),
	.b(n246102));
   no02f02 U262333 (.o(n246102),
	.a(n246101),
	.b(n246103));
   na02f06 U262334 (.o(n252824),
	.a(n249317),
	.b(n246909));
   na02m02 U262335 (.o(n246148),
	.a(n246145),
	.b(n246144));
   na02f01 U262336 (.o(n246140),
	.a(n246137),
	.b(n246136));
   no02f01 U262338 (.o(n246831),
	.a(n246805),
	.b(n246794));
   in01f02 U262339 (.o(n246737),
	.a(n246738));
   no02f03 U262340 (.o(n248977),
	.a(n248953),
	.b(n249081));
   na02f02 U262341 (.o(n245986),
	.a(n245985),
	.b(n245984));
   no02f01 U262342 (.o(n246165),
	.a(n246161),
	.b(n246162));
   no02m02 U262343 (.o(n246736),
	.a(n246735),
	.b(n246734));
   ao12f02 U262345 (.o(n246735),
	.a(n249012),
	.b(n249014),
	.c(n246730));
   no02m02 U262346 (.o(n246789),
	.a(n246781),
	.b(n246780));
   no02f04 U262347 (.o(n249020),
	.a(n246798),
	.b(n246799));
   in01f08 U262348 (.o(n252157),
	.a(FE_OFN346_n252141));
   in01f08 U262350 (.o(n251548),
	.a(FE_OFN204_n251530));
   in01f06 U262351 (.o(n251796),
	.a(FE_OFN432_n251781));
   in01f08 U262352 (.o(n250378),
	.a(FE_OFN410_n250360));
   in01f08 U262353 (.o(n250237),
	.a(FE_OFN276_n250218));
   in01f08 U262355 (.o(n251477),
	.a(FE_OFN322_n251459));
   in01f08 U262356 (.o(n250945),
	.a(FE_OFN418_n250930));
   in01f08 U262358 (.o(n250981),
	.a(FE_OFN200_n250965));
   in01f08 U262361 (.o(n252120),
	.a(FE_OFN208_n252105));
   in01f06 U262362 (.o(n250662),
	.a(FE_OFN414_n250646));
   in01f08 U262364 (.o(n251016),
	.a(FE_OFN302_n251001));
   in01f08 U262366 (.o(n252193),
	.a(FE_OFN348_n252178));
   in01f08 U262368 (.o(n250591),
	.a(FE_OFN412_n250576));
   in01f08 U262370 (.o(n251513),
	.a(FE_OFN428_n251494));
   in01f06 U262371 (.o(n250162),
	.a(FE_OFN272_n250144));
   in01f08 U262372 (.o(n250413),
	.a(FE_OFN195_n250395));
   in01f08 U262373 (.o(n251442),
	.a(FE_OFN426_n251424));
   in01f08 U262374 (.o(n252230),
	.a(FE_OFN350_n252215));
   in01f08 U262375 (.o(n251832),
	.a(FE_OFN206_n251816));
   in01f06 U262376 (.o(n251051),
	.a(FE_OFN304_n251036));
   in01f06 U262377 (.o(n250626),
	.a(FE_OFN290_n250611));
   in01f06 U262379 (.o(n251902),
	.a(FE_OFN337_n251887));
   in01f06 U262380 (.o(n250198),
	.a(FE_OFN274_n250180));
   in01f06 U262381 (.o(n250053),
	.a(FE_OFN270_n250035));
   in01f08 U262382 (.o(n251655),
	.a(FE_OFN329_n251637));
   in01f10 U262383 (.o(n251158),
	.a(FE_OFN420_n251140));
   in01f08 U262385 (.o(n250307),
	.a(FE_OFN408_n250289));
   in01f04 U262386 (.o(n249824),
	.a(n245472));
   in01f08 U262387 (.o(n250732),
	.a(FE_OFN292_n250717));
   in01f06 U262388 (.o(n250556),
	.a(FE_OFN288_n250540));
   no02f02 U262389 (.o(n249014),
	.a(n246778),
	.b(n246728));
   in01f08 U262390 (.o(n250875),
	.a(FE_OFN416_n250859));
   in01f06 U262391 (.o(n250343),
	.a(FE_OFN280_n250324));
   in01f06 U262392 (.o(n251194),
	.a(FE_OFN311_n251175));
   in01f06 U262393 (.o(n250839),
	.a(n250824));
   in01f06 U262394 (.o(n252048),
	.a(FE_OFN343_n252032));
   in01f08 U262395 (.o(n251726),
	.a(FE_OFN430_n251710));
   in01f06 U262396 (.o(n250768),
	.a(FE_OFN294_n250752));
   in01f03 U262397 (.o(n251300),
	.a(FE_OFN314_n251281));
   in01f06 U262398 (.o(n251975),
	.a(FE_OFN341_n251960));
   na02f02 U262399 (.o(n246098),
	.a(n246097),
	.b(n246096));
   na02f01 U262400 (.o(n252640),
	.a(n252758),
	.b(n252642));
   in01f06 U262401 (.o(n251690),
	.a(FE_OFN331_n251675));
   in01f06 U262402 (.o(n251264),
	.a(FE_OFN202_n251246));
   no02f03 U262403 (.o(n246798),
	.a(n246788),
	.b(n246787));
   in01f06 U262404 (.o(n249982),
	.a(n249964));
   no02s01 U262405 (.o(n246901),
	.a(n252382),
	.b(n246900));
   in01f08 U262406 (.o(n250520),
	.a(n250502));
   in01f06 U262407 (.o(n251407),
	.a(FE_OFN320_n251388));
   in01f06 U262408 (.o(n250126),
	.a(FE_OFN193_n250107));
   in01f08 U262409 (.o(n250697),
	.a(FE_OFN197_n250682));
   in01f08 U262410 (.o(n251088),
	.a(FE_OFN307_n251072));
   in01f08 U262411 (.o(n250449),
	.a(FE_OFN282_n250430));
   in01f08 U262412 (.o(n251583),
	.a(FE_OFN324_n251565));
   in01f06 U262413 (.o(n250910),
	.a(FE_OFN300_n250895));
   in01f08 U262415 (.o(n251371),
	.a(FE_OFN318_n251353));
   na02f04 U262416 (.o(n252232),
	.a(n246204),
	.b(n245778));
   in01f06 U262417 (.o(n251761),
	.a(FE_OFN333_n251746));
   in01f06 U262418 (.o(n250089),
	.a(FE_OFN404_n250071));
   in01f06 U262419 (.o(n251123),
	.a(FE_OFN309_n251105));
   in01f06 U262420 (.o(n252084),
	.a(FE_OFN437_n252069));
   na02f01 U262421 (.o(n252338),
	.a(n252352),
	.b(n252775));
   in01f08 U262422 (.o(n251939),
	.a(FE_OFN339_n251923));
   no02f01 U262424 (.o(n251353),
	.a(n252196),
	.b(FE_OFN28_n251337));
   no02f03 U262425 (.o(n250466),
	.a(FE_OFN210_n252159),
	.b(FE_OFN24_n250486));
   no02f01 U262427 (.o(n251494),
	.a(n252050),
	.b(n251621));
   no02f01 U262429 (.o(n250611),
	.a(n252013),
	.b(FE_OFN556_n250770));
   no02f01 U262430 (.o(n250324),
	.a(n252013),
	.b(FE_OFN24_n250486));
   no02f01 U262431 (.o(n251246),
	.a(n252086),
	.b(FE_OFN28_n251337));
   no02f01 U262432 (.o(n251530),
	.a(n252086),
	.b(n251621));
   no02f01 U262434 (.o(n251960),
	.a(n251941),
	.b(n252195));
   no02f01 U262435 (.o(n251637),
	.a(n252196),
	.b(n251621));
   no02f01 U262439 (.o(n251852),
	.a(n252122),
	.b(FE_OFN33_n251904));
   no02f01 U262440 (.o(n250646),
	.a(n252050),
	.b(n250770));
   no02f03 U262441 (.o(n251887),
	.a(FE_OFN210_n252159),
	.b(FE_OFN32_n251904));
   no02f01 U262442 (.o(n251281),
	.a(n252122),
	.b(FE_OFN28_n251337));
   no02f01 U262443 (.o(n251600),
	.a(FE_OFN210_n252159),
	.b(n251621));
   no02f01 U262444 (.o(n250752),
	.a(FE_OFN210_n252159),
	.b(FE_OFN556_n250770));
   no02f01 U262445 (.o(n251317),
	.a(FE_OFN210_n252159),
	.b(FE_OFN28_n251337));
   no02f01 U262446 (.o(n250540),
	.a(n251941),
	.b(FE_OFN556_n250770));
   no02f01 U262447 (.o(n251424),
	.a(n251977),
	.b(n251621));
   no02f01 U262449 (.o(n251816),
	.a(n252086),
	.b(FE_OFN32_n251904));
   no02f01 U262450 (.o(n250360),
	.a(n252050),
	.b(FE_OFN24_n250486));
   no02f01 U262451 (.o(n251675),
	.a(n251941),
	.b(FE_OFN32_n251904));
   no02f01 U262453 (.o(n251459),
	.a(n252013),
	.b(n251621));
   no02f01 U262454 (.o(n251565),
	.a(n252122),
	.b(n251621));
   no02f01 U262455 (.o(n251388),
	.a(n251941),
	.b(n251621));
   no02f01 U262456 (.o(n250717),
	.a(n252122),
	.b(n250770));
   no02f01 U262457 (.o(n251781),
	.a(n252050),
	.b(FE_OFN32_n251904));
   no02f01 U262458 (.o(n250576),
	.a(n251977),
	.b(n250770));
   no02f01 U262460 (.o(n250395),
	.a(n252086),
	.b(FE_OFN24_n250486));
   no02f01 U262461 (.o(n251923),
	.a(n252196),
	.b(FE_OFN32_n251904));
   no02f02 U262462 (.o(n251710),
	.a(n251977),
	.b(FE_OFN33_n251904));
   no02f08 U262463 (.o(n250502),
	.a(n252196),
	.b(FE_OFN24_n250486));
   no02f01 U262464 (.o(n250430),
	.a(n252122),
	.b(FE_OFN24_n250486));
   no02f02 U262466 (.o(n250071),
	.a(FE_OFN22_n250202),
	.b(n252050));
   no02f01 U262467 (.o(n251001),
	.a(n252122),
	.b(n251053));
   no02f01 U262468 (.o(n252141),
	.a(n252122),
	.b(n252195));
   no02f01 U262470 (.o(n250180),
	.a(FE_OFN22_n250202),
	.b(FE_OFN210_n252159));
   no02f01 U262471 (.o(n252178),
	.a(FE_OFN210_n252159),
	.b(n252195));
   no02f01 U262473 (.o(n251175),
	.a(n252013),
	.b(FE_OFN28_n251337));
   no02f01 U262474 (.o(n250859),
	.a(n251977),
	.b(n251053));
   no02f01 U262476 (.o(n252215),
	.a(n252196),
	.b(n252195));
   no02f04 U262477 (.o(n250824),
	.a(n251941),
	.b(n251053));
   no02f02 U262478 (.o(n249964),
	.a(n251941),
	.b(FE_OFN22_n250202));
   no02f01 U262479 (.o(n250107),
	.a(FE_OFN22_n250202),
	.b(n252086));
   no02f06 U262481 (.o(n249999),
	.a(FE_OFN22_n250202),
	.b(n251977));
   no02f01 U262482 (.o(n251036),
	.a(FE_OFN210_n252159),
	.b(n251053));
   no02f01 U262483 (.o(n250930),
	.a(n252050),
	.b(n251053));
   no02f01 U262484 (.o(n250035),
	.a(FE_OFN22_n250202),
	.b(n252013));
   no02f01 U262485 (.o(n251140),
	.a(n251977),
	.b(FE_OFN28_n251337));
   no02f01 U262486 (.o(n250789),
	.a(n252196),
	.b(n250770));
   no02f01 U262487 (.o(n250965),
	.a(n252086),
	.b(n251053));
   no02f01 U262488 (.o(n251072),
	.a(n252196),
	.b(n251053));
   no02f01 U262489 (.o(n250289),
	.a(n251977),
	.b(FE_OFN24_n250486));
   no02f01 U262490 (.o(n251996),
	.a(n251977),
	.b(n252195));
   no02f01 U262492 (.o(n252032),
	.a(n252013),
	.b(n252195));
   no02f01 U262493 (.o(n250895),
	.a(n252013),
	.b(n251053));
   no02f02 U262494 (.o(n251105),
	.a(n251941),
	.b(FE_OFN28_n251337));
   no02f01 U262495 (.o(n252105),
	.a(n252086),
	.b(n252195));
   no02f01 U262496 (.o(n250218),
	.a(FE_OFN22_n250202),
	.b(n252196));
   in01s02 U262498 (.o(n252764),
	.a(n252341));
   no02f01 U262499 (.o(n252069),
	.a(n252050),
	.b(n252195));
   no02f01 U262500 (.o(n250254),
	.a(n251941),
	.b(FE_OFN24_n250486));
   no02f01 U262501 (.o(n248129),
	.a(n247069),
	.b(FE_OFN32_n251904));
   na02s01 U262502 (.o(n245515),
	.a(n245529),
	.b(n246899));
   no02f06 U262503 (.o(n249640),
	.a(n249698),
	.b(n245470));
   na02f04 U262504 (.o(n246782),
	.a(n249007),
	.b(n246360));
   na02s01 U262505 (.o(n246900),
	.a(n246899),
	.b(n252379));
   na02f01 U262506 (.o(n245487),
	.a(n245447),
	.b(n245490));
   no02f01 U262507 (.o(n248126),
	.a(n247069),
	.b(n251621));
   no02f01 U262508 (.o(n248362),
	.a(n247069),
	.b(FE_OFN24_n250486));
   no02f01 U262509 (.o(n248364),
	.a(n247069),
	.b(n252195));
   no02f01 U262510 (.o(n248363),
	.a(n247069),
	.b(n251053));
   no02f01 U262511 (.o(n248127),
	.a(n247069),
	.b(FE_OFN28_n251337));
   no02f01 U262512 (.o(n248128),
	.a(n247069),
	.b(FE_OFN556_n250770));
   no02s01 U262513 (.o(n245421),
	.a(n245423),
	.b(n245422));
   na02f04 U262514 (.o(n247094),
	.a(FE_OFN516_regtop_v1_hdi00_a_0_),
	.b(n247091));
   in01f01 U262515 (.o(n245479),
	.a(n249698));
   no02f02 U262516 (.o(n245939),
	.a(n245529),
	.b(n245528));
   na02f02 U262517 (.o(n246902),
	.a(n245537),
	.b(n246845));
   no03f02 U262518 (.o(n246727),
	.a(n246726),
	.b(n246785),
	.c(n246725));
   na02f03 U262519 (.o(n246785),
	.a(n246356),
	.b(n246355));
   na02f02 U262520 (.o(n246914),
	.a(n246354),
	.b(n246353));
   na02s01 U262521 (.o(n246610),
	.a(n252684),
	.b(n246609));
   ao22s01 U262523 (.o(n249475),
	.a(g_hs60p_r[5]),
	.b(FE_OFN398_n249646),
	.c(n249548),
	.d(1'b1));
   ao22s01 U262524 (.o(n249526),
	.a(n249548),
	.b(1'b1),
	.c(n253014),
	.d(g_cbcr_offset_r[9]));
   ao22s01 U262525 (.o(n249487),
	.a(n249548),
	.b(1'b1),
	.c(n249638),
	.d(regtop_g_tc_r[4]));
   ao22s01 U262526 (.o(n249550),
	.a(n249548),
	.b(1'b1),
	.c(n253014),
	.d(g_cbcr_offset_r[8]));
   ao22s01 U262527 (.o(n249448),
	.a(n249548),
	.b(1'b1),
	.c(n249584),
	.d(regtop_g_nfst_r[15]));
   ao22s01 U262529 (.o(n249493),
	.a(n249547),
	.b(regtop_g_icdc_r),
	.c(n249548),
	.d(1'b1));
   no02m02 U262530 (.o(n245568),
	.a(n245550),
	.b(n246902));
   ao12f01 U262531 (.o(n245559),
	.a(n245552),
	.b(n245763),
	.c(n245553));
   oa12f04 U262532 (.o(n244966),
	.a(n249661),
	.b(n245444),
	.c(n249662));
   oa12f04 U262533 (.o(n245599),
	.a(n245605),
	.b(n245607),
	.c(n245604));
   ao12f02 U262535 (.o(n249035),
	.a(n249072),
	.b(n249034),
	.c(n249073));
   in01f01 U262536 (.o(n246237),
	.a(v1_bs_req_n));
   in01m01 U262537 (.o(n246145),
	.a(n246143));
   no02m02 U262538 (.o(n246143),
	.a(n246122),
	.b(n246121));
   oa12f02 U262539 (.o(n244989),
	.a(n249058),
	.b(n249077),
	.c(FE_OFN532_regtop_g_a_r_5_));
   na02f02 U262540 (.o(n249055),
	.a(n249037),
	.b(n249053));
   ao12f02 U262541 (.o(n249049),
	.a(n249072),
	.b(n249048),
	.c(n249073));
   oa12f02 U262542 (.o(n244988),
	.a(n249049),
	.b(n249077),
	.c(FE_OFN517_regtop_g_a_r_6_));
   na02f02 U262543 (.o(n246119),
	.a(regtop_g_udb2_r[5]),
	.b(n246124));
   ao12f02 U262545 (.o(n249075),
	.a(n249072),
	.b(n249074),
	.c(n249073));
   na03m02 U262546 (.o(n247489),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247487));
   na03m02 U262547 (.o(n247343),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247342));
   na03m02 U262548 (.o(n247484),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247483));
   na03m02 U262549 (.o(n247586),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247585));
   na03m02 U262550 (.o(n247321),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247320));
   na03f01 U262551 (.o(n247325),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247494),
	.c(n247324));
   na02f04 U262552 (.o(n246845),
	.a(regtop_g_paramadr_r[3]),
	.b(n245527));
   in01s01 U262553 (.o(n247015),
	.a(n246891));
   na02s02 U262554 (.o(n246891),
	.a(n246890),
	.b(n246025));
   no02f02 U262555 (.o(n247024),
	.a(n246998),
	.b(n246997));
   no02f01 U262556 (.o(n249646),
	.a(regtop_g_a_r[3]),
	.b(n245477));
   no02f01 U262557 (.o(n245773),
	.a(n246943),
	.b(n245772));
   no02f06 U262559 (.o(n252684),
	.a(regtop_g_paramadr_r[6]),
	.b(regtop_g_paramadr_r[4]));
   oa22s01 U262560 (.o(n246417),
	.a(n246430),
	.b(n246527),
	.c(n246528),
	.d(n246693));
   ao12f02 U262561 (.o(n247027),
	.a(n247006),
	.b(n247008),
	.c(n247007));
   no03f01 U262562 (.o(n245443),
	.a(regtop_g_ms_r_n),
	.b(regtop_g_memr_ok_r),
	.c(regtop_g_read_r_n));
   no02f03 U262563 (.o(n245420),
	.a(g_field_start_add_r[27]),
	.b(busrtop_b_rreq_vrh_rrq_fldstatadd_r[27]));
   na02f01 U262564 (.o(n246457),
	.a(n246570),
	.b(n246345));
   na02f02 U262565 (.o(n246464),
	.a(n246700),
	.b(vldtop_vld_syndec_ADP[4]));
   na02s02 U262566 (.o(n246466),
	.a(n246568),
	.b(vldtop_vld_syndec_ADP[4]));
   in01f02 U262567 (.o(n246697),
	.a(n246565));
   no02f02 U262568 (.o(n246707),
	.a(n246011),
	.b(n246010));
   no02s02 U262569 (.o(n249870),
	.a(n249878),
	.b(n249871));
   ao12f06 U262570 (.o(n249668),
	.a(n249664),
	.b(n249738),
	.c(regtop_g_ispi_r));
   in01s01 U262571 (.o(n249685),
	.a(n249664));
   ao12f02 U262572 (.o(n249752),
	.a(n245444),
	.b(n249727),
	.c(n249726));
   ao12s01 U262573 (.o(n249726),
	.a(n249723),
	.b(n249725),
	.c(n249724));
   no02f08 U262574 (.o(n249548),
	.a(n245481),
	.b(n245480));
   no02f03 U262575 (.o(n249635),
	.a(n245471),
	.b(n245470));
   no02f08 U262576 (.o(n249638),
	.a(n245471),
	.b(n249697));
   no02f06 U262577 (.o(n249628),
	.a(n252286),
	.b(n245471));
   no02f06 U262578 (.o(n249629),
	.a(n245471),
	.b(n245461));
   ao22f01 U262579 (.o(n249212),
	.a(n249211),
	.b(regtop_g_paramdata_r[11]),
	.c(n249210),
	.d(regtop_g_paramdata_r[15]));
   na02s01 U262580 (.o(n246186),
	.a(n252462),
	.b(n246194));
   in01s01 U262581 (.o(n247595),
	.a(n246201));
   in01f01 U262582 (.o(n249588),
	.a(n249645));
   no03f01 U262583 (.o(n245580),
	.a(n245579),
	.b(n252239),
	.c(n245578));
   in01f01 U262584 (.o(n252254),
	.a(n252462));
   no02f02 U262585 (.o(n245579),
	.a(regtop_g_paramadr_r[4]),
	.b(n245531));
   na02f02 U262586 (.o(n245531),
	.a(n246608),
	.b(n252380));
   na02f02 U262587 (.o(n249082),
	.a(n249135),
	.b(n246617));
   no02f01 U262588 (.o(n246170),
	.a(regtop_g_udb2_r[0]),
	.b(n246169));
   ao22s01 U262589 (.o(n246309),
	.a(n246570),
	.b(n246699),
	.c(n246568),
	.d(n246712));
   no02f02 U262590 (.o(n247023),
	.a(n247022),
	.b(n247021));
   na02f01 U262591 (.o(n247021),
	.a(n247020),
	.b(n247019));
   na02f01 U262592 (.o(n246973),
	.a(n246989),
	.b(n246972));
   no02s02 U262593 (.o(n246972),
	.a(n246971),
	.b(n246970));
   na02s02 U262594 (.o(n246970),
	.a(n246988),
	.b(n246969));
   no03f01 U262595 (.o(n246979),
	.a(n246980),
	.b(n246982),
	.c(n246966));
   ao12f02 U262619 (.o(n245355),
	.a(n245353),
	.b(n245665),
	.c(n245354));
   na02f02 U262620 (.o(n245356),
	.a(n245666),
	.b(n245354));
   no02f02 U262621 (.o(n245354),
	.a(n245667),
	.b(n245702));
   in01s01 U262622 (.o(n249871),
	.a(vh_1_ph_add[6]));
   na04f02 U262623 (.o(n245478),
	.a(n245476),
	.b(n245475),
	.c(n245474),
	.d(n245473));
   ao22s01 U262624 (.o(n249599),
	.a(FE_OFN552_n245462),
	.b(regtop_g_vd_r[6]),
	.c(n249812),
	.d(regtop_g_tmc_r[6]));
   oa12s01 U262625 (.o(n249603),
	.a(n249583),
	.b(n249827),
	.c(n252884));
   ao12s01 U262626 (.o(n249583),
	.a(n249664),
	.b(regtop_g_mem_rd2_r[6]),
	.c(regtop_g_memr_ok_r));
   ao22f01 U262627 (.o(n249618),
	.a(FE_OFN545_n245460),
	.b(regtop_g_brv_r[5]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcvo0_r[5]));
   ao22f02 U262628 (.o(n249672),
	.a(n249731),
	.b(g_field_offset_r[2]),
	.c(n249732),
	.d(g_cbcr_offset_r[2]));
   ao22s01 U262629 (.o(n249671),
	.a(n249812),
	.b(regtop_g_tmc_r[2]),
	.c(n249757),
	.d(regtop_g_scp_r[2]));
   ao22s01 U262630 (.o(n249695),
	.a(n249812),
	.b(regtop_g_tmc_r[1]),
	.c(n249757),
	.d(regtop_g_scp_r[1]));
   na04f02 U262631 (.o(n249805),
	.a(n249804),
	.b(n249803),
	.c(n249802),
	.d(n249801));
   na04f01 U262632 (.o(n249796),
	.a(n249795),
	.b(n249794),
	.c(n249793),
	.d(n249792));
   na04f01 U262634 (.o(n249765),
	.a(n249761),
	.b(n249760),
	.c(n249759),
	.d(n249758));
   na02f06 U262635 (.o(n249242),
	.a(n252684),
	.b(n248985));
   na02f10 U262636 (.o(n249250),
	.a(n252684),
	.b(n249066));
   ao12f02 U262637 (.o(n245776),
	.a(n246060),
	.b(n246197),
	.c(n245775));
   no03f02 U262638 (.o(n246933),
	.a(n246930),
	.b(n247050),
	.c(n246929));
   no03m02 U262639 (.o(n246427),
	.a(n246418),
	.b(n246417),
	.c(n246416));
   na02f08 U262640 (.o(n246088),
	.a(regtop_g_udb1_r[3]),
	.b(regtop_g_udb2_r[3]));
   na02f01 U262641 (.o(n246071),
	.a(regtop_g_udb0_r[2]),
	.b(n246077));
   na02f01 U262642 (.o(n246072),
	.a(n246070),
	.b(n246077));
   in01f01 U262643 (.o(n246074),
	.a(n246073));
   na02f04 U262644 (.o(n246152),
	.a(n246087),
	.b(n246086));
   no02s01 U262645 (.o(n245413),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[26]),
	.b(g_field_start_add_r[26]));
   no02s01 U262646 (.o(n245403),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[24]),
	.b(g_field_start_add_r[24]));
   no02s01 U262647 (.o(n245394),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[23]),
	.b(g_field_start_add_r[23]));
   no02s01 U262648 (.o(n245391),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[22]),
	.b(g_field_start_add_r[22]));
   no02f01 U262649 (.o(n245382),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[21]),
	.b(g_field_start_add_r[21]));
   no02f01 U262650 (.o(n245364),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[19]),
	.b(g_field_start_add_r[19]));
   no02f02 U262651 (.o(n245360),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[17]),
	.b(g_field_start_add_r[17]));
   na02f01 U262652 (.o(n245770),
	.a(n245769),
	.b(n245768));
   no02s01 U262653 (.o(n246553),
	.a(n246498),
	.b(n246693));
   ao22s01 U262654 (.o(n246488),
	.a(n246512),
	.b(n246528),
	.c(n246511),
	.d(n246526));
   oa22s01 U262655 (.o(n246486),
	.a(n246485),
	.b(n246525),
	.c(n246484),
	.d(n246483));
   no02s02 U262656 (.o(n246992),
	.a(n246991),
	.b(n246990));
   na02s02 U262657 (.o(n246990),
	.a(n246989),
	.b(n246988));
   no02s02 U262658 (.o(n246999),
	.a(n247017),
	.b(n247009));
   na04f02 U262659 (.o(n246996),
	.a(n246986),
	.b(n246985),
	.c(n246984),
	.d(n246983));
   no02f02 U262660 (.o(n246969),
	.a(n246987),
	.b(n246968));
   no02f02 U262661 (.o(n245348),
	.a(n245334),
	.b(n245333));
   no02f02 U262662 (.o(n245334),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[15]),
	.b(n245341));
   no02f02 U262663 (.o(n245333),
	.a(g_field_start_add_r[15]),
	.b(n245341));
   na02s01 U262664 (.o(n245895),
	.a(vh_1_ph_add[6]),
	.b(vh_1_ph_add[7]));
   oa12f01 U262665 (.o(n245886),
	.a(n245857),
	.b(n245856),
	.c(n245853));
   ao12s01 U262666 (.o(n245859),
	.a(n245854),
	.b(n245899),
	.c(n245855));
   na03f06 U262667 (.o(n251941),
	.a(regtop_v1_hdi00_a[1]),
	.b(regtop_v1_hdi00_a[0]),
	.c(n250055));
   na03f04 U262668 (.o(n252013),
	.a(regtop_v1_hdi00_a[0]),
	.b(n250055),
	.c(n250164));
   na03f06 U262669 (.o(n252086),
	.a(regtop_v1_hdi00_a[1]),
	.b(regtop_v1_hdi00_a[0]),
	.c(n250200));
   na02f01 U262670 (.o(n245530),
	.a(n252462),
	.b(n245551));
   no02f01 U262671 (.o(n252576),
	.a(n246193),
	.b(n246192));
   na03s01 U262672 (.o(n246193),
	.a(regtop_g_adb_r[2]),
	.b(regtop_g_adb_r[6]),
	.c(regtop_g_adb_r[4]));
   na02f01 U262673 (.o(n252564),
	.a(n245761),
	.b(n252404));
   no02f03 U262674 (.o(n245527),
	.a(regtop_g_paramadr_r[5]),
	.b(regtop_g_paramadr_r[7]));
   in01f02 U262675 (.o(n249241),
	.a(n249138));
   oa22f01 U262676 (.o(n246401),
	.a(n246379),
	.b(n246695),
	.c(n246380),
	.d(n246527));
   no02s01 U262677 (.o(n246446),
	.a(n246338),
	.b(n246695));
   na02s02 U262678 (.o(n245975),
	.a(n245974),
	.b(n245973));
   ao22s01 U262679 (.o(n246448),
	.a(n246700),
	.b(n246344),
	.c(n246570),
	.d(n246465));
   oa22s01 U262680 (.o(n246051),
	.a(n246535),
	.b(n246578),
	.c(n246435),
	.d(n246714));
   oa22s01 U262681 (.o(n246580),
	.a(n246575),
	.b(n246708),
	.c(n246714),
	.d(n246574));
   ao22s01 U262682 (.o(n246573),
	.a(n246570),
	.b(n246569),
	.c(n246568),
	.d(n246567));
   in01s01 U262683 (.o(n246343),
	.a(n246339));
   ao22s01 U262684 (.o(n246339),
	.a(n246706),
	.b(n246338),
	.c(n246658),
	.d(n246337));
   oa22s01 U262685 (.o(n246342),
	.a(n246714),
	.b(n246341),
	.c(n246711),
	.d(n246340));
   na02s01 U262686 (.o(n246347),
	.a(n246570),
	.b(n246463));
   in01s01 U262687 (.o(n246439),
	.a(n246438));
   oa22s01 U262688 (.o(n246437),
	.a(n246536),
	.b(n246578),
	.c(n246535),
	.d(n246711));
   oa22s01 U262689 (.o(n246436),
	.a(n246533),
	.b(n246714),
	.c(n246435),
	.d(n246708));
   no02s01 U262690 (.o(n246440),
	.a(n246434),
	.b(n246433));
   oa22s01 U262691 (.o(n246313),
	.a(n246714),
	.b(n246340),
	.c(n246708),
	.d(n246341));
   oa22s01 U262692 (.o(n246314),
	.a(n246578),
	.b(n246344),
	.c(n246711),
	.d(n246312));
   ao22s01 U262693 (.o(n246517),
	.a(n246694),
	.b(n246516),
	.c(n246515),
	.d(n246514));
   ao22s01 U262694 (.o(n246518),
	.a(n246513),
	.b(n246512),
	.c(n246698),
	.d(n246511));
   oa22s01 U262695 (.o(n246396),
	.a(n246709),
	.b(n246714),
	.c(n246394),
	.d(n246708));
   oa22s01 U262696 (.o(n246469),
	.a(n246468),
	.b(n246484),
	.c(n246485),
	.d(n246467));
   oa22s01 U262697 (.o(n246470),
	.a(n246466),
	.b(n246465),
	.c(n246464),
	.d(n246463));
   no03f01 U262698 (.o(n246404),
	.a(n246403),
	.b(n246402),
	.c(n246401));
   in01s01 U262699 (.o(n246515),
	.a(n246484));
   no02f01 U262700 (.o(n247020),
	.a(n246055),
	.b(n245986));
   na02s01 U262701 (.o(n246796),
	.a(v_vldstatus_r[1]),
	.b(n249021));
   na02f01 U262702 (.o(n246882),
	.a(v_vldstatus_r[0]),
	.b(n246898));
   no02f01 U262703 (.o(n247003),
	.a(n246887),
	.b(n246886));
   no02f06 U262704 (.o(n245619),
	.a(n245417),
	.b(n245416));
   no02f04 U262705 (.o(n245634),
	.a(n245405),
	.b(n245404));
   na02f04 U262706 (.o(n245635),
	.a(n245405),
	.b(n245404));
   in01s01 U262707 (.o(n245643),
	.a(n245397));
   no02f04 U262708 (.o(n245649),
	.a(n245393),
	.b(n245392));
   ao12f02 U262709 (.o(n245676),
	.a(n245371),
	.b(n245688),
	.c(n245372));
   in01f01 U262710 (.o(n245372),
	.a(n245720));
   na02f02 U262711 (.o(n245677),
	.a(n245688),
	.b(n245721));
   in01f01 U262712 (.o(n245688),
	.a(n245359));
   no02f01 U262713 (.o(n245359),
	.a(n245370),
	.b(n245369));
   na02f01 U262714 (.o(n245668),
	.a(n245352),
	.b(n245351));
   na02m02 U262715 (.o(n245703),
	.a(n245350),
	.b(n245349));
   no02f02 U262716 (.o(n245702),
	.a(n245350),
	.b(n245349));
   no02f02 U262717 (.o(n245712),
	.a(n245348),
	.b(n245347));
   na02f01 U262718 (.o(n245713),
	.a(n245348),
	.b(n245347));
   no02f02 U262720 (.o(n245332),
	.a(n245735),
	.b(n245743));
   na04s01 U262721 (.o(n245992),
	.a(n245991),
	.b(n245990),
	.c(n245989),
	.d(n245988));
   na04s01 U262722 (.o(n245997),
	.a(n245996),
	.b(n245995),
	.c(n245994),
	.d(n245993));
   ao12s01 U262723 (.o(n249849),
	.a(n249848),
	.b(vh_1_ph_add[9]),
	.c(n249855));
   oa12s01 U262724 (.o(n249848),
	.a(n249916),
	.b(vh_1_ph_add[9]),
	.c(n249855));
   ao12s01 U262725 (.o(n249857),
	.a(n249855),
	.b(n249863),
	.c(n249856));
   oa12s01 U262726 (.o(n249864),
	.a(n249863),
	.b(n249870),
	.c(vh_1_ph_add[7]));
   ao12s01 U262727 (.o(n249872),
	.a(n249870),
	.b(n249878),
	.c(n249871));
   in01f02 U262728 (.o(n249913),
	.a(n246230));
   in01f02 U262729 (.o(n249916),
	.a(n246234));
   no02f01 U262730 (.o(n249273),
	.a(n249272),
	.b(busrtop_b_rreq_vrh_add1_r[8]));
   in01f01 U262731 (.o(n249924),
	.a(n246002));
   na04f02 U262732 (.o(n245574),
	.a(n245559),
	.b(n252489),
	.c(n252547),
	.d(n252491));
   ao22f02 U262733 (.o(n249784),
	.a(FE_OFN4_n245443),
	.b(n249781),
	.c(g_hsdc_r[0]),
	.d(n249786));
   na03f02 U262734 (.o(n249781),
	.a(n249780),
	.b(n249779),
	.c(n249778));
   ao22f02 U262735 (.o(n249611),
	.a(n249812),
	.b(regtop_g_tmc_r[5]),
	.c(regtop_g_scp_r[5]),
	.d(n249757));
   na04f02 U262736 (.o(n249657),
	.a(n249656),
	.b(n249655),
	.c(n249654),
	.d(n249653));
   na04f02 U262737 (.o(n249658),
	.a(n249644),
	.b(n249643),
	.c(n249642),
	.d(n249641));
   no02f04 U262738 (.o(n249841),
	.a(n245444),
	.b(FE_OFN544_n252912));
   no04f02 U262739 (.o(n249753),
	.a(n249752),
	.b(n249751),
	.c(n249750),
	.d(n249749));
   no03f08 U262740 (.o(n249944),
	.a(n249930),
	.b(regtop_g_prev_efbst_r),
	.c(regtop_g_prev_enfst_r));
   na04f03 U262741 (.o(n249563),
	.a(n249552),
	.b(n249551),
	.c(n249550),
	.d(n249549));
   no02m02 U262742 (.o(n249928),
	.a(regtop_g_prev_efbst_r),
	.b(n249924));
   in01s01 U262743 (.o(n249926),
	.a(n249929));
   no02f08 U262744 (.o(n249812),
	.a(n245444),
	.b(n249396));
   in01f08 U262745 (.o(n249811),
	.a(n249827));
   na02f03 U262746 (.o(n249763),
	.a(FE_OFN4_n245443),
	.b(FE_OFN396_n249640));
   in01f04 U262747 (.o(n249786),
	.a(n249829));
   no02f04 U262749 (.o(n249836),
	.a(n245444),
	.b(n249789));
   na04f02 U262750 (.o(n249445),
	.a(n249439),
	.b(n249438),
	.c(n249437),
	.d(n249436));
   no02f02 U262751 (.o(n249072),
	.a(n246061),
	.b(n252542));
   in01f02 U262752 (.o(n249031),
	.a(n249039));
   no02f01 U262753 (.o(n249193),
	.a(n249189),
	.b(n252656));
   no02f01 U262754 (.o(n249179),
	.a(n249189),
	.b(n252660));
   no02f01 U262755 (.o(n249173),
	.a(n249189),
	.b(n252662));
   no02f01 U262756 (.o(n249167),
	.a(n249189),
	.b(n252664));
   no02f01 U262757 (.o(n249161),
	.a(n249189),
	.b(n252666));
   no02f01 U262758 (.o(n249156),
	.a(n249189),
	.b(n252778));
   no02f01 U262759 (.o(n249151),
	.a(n249189),
	.b(n252755));
   in01s01 U262760 (.o(n249199),
	.a(n249198));
   oa22f01 U262761 (.o(n249126),
	.a(FE_OFN483_n249211),
	.b(n252664),
	.c(n249242),
	.d(n252778));
   ao22s01 U262762 (.o(n249102),
	.a(n249211),
	.b(regtop_g_paramdata_r[23]),
	.c(n249127),
	.d(regtop_g_atscd_r[20]));
   ao22s01 U262763 (.o(n249122),
	.a(n249211),
	.b(regtop_g_paramdata_r[24]),
	.c(n249127),
	.d(regtop_g_atscd_r[21]));
   in01f02 U262764 (.o(n249127),
	.a(n249078));
   in01f04 U262765 (.o(n249128),
	.a(n249079));
   ao12s01 U262766 (.o(n249097),
	.a(n249095),
	.b(n249127),
	.c(regtop_g_atscd_r[17]));
   oa22s01 U262767 (.o(n249095),
	.a(FE_OFN483_n249211),
	.b(n252662),
	.c(n249242),
	.d(n252666));
   na02f02 U262768 (.o(n252260),
	.a(n252270),
	.b(regtop_g_wd_r[17]));
   in01f02 U262769 (.o(n252269),
	.a(n252273));
   no03f01 U262770 (.o(n252289),
	.a(n245794),
	.b(n245793),
	.c(n245792));
   na02s01 U262771 (.o(n245792),
	.a(n252908),
	.b(n245791));
   oa22f01 U262772 (.o(n252302),
	.a(n252253),
	.b(n252252),
	.c(n252251),
	.d(n252254));
   in01s01 U262773 (.o(n252300),
	.a(n252305));
   oa22f01 U262774 (.o(n252307),
	.a(n245588),
	.b(n252252),
	.c(regtop_g_paramadr_r[1]),
	.d(n252251));
   na02f02 U262775 (.o(n247039),
	.a(n246949),
	.b(n246920));
   na02f02 U262776 (.o(n247040),
	.a(n247034),
	.b(n247033));
   na02s02 U262777 (.o(n247033),
	.a(n247042),
	.b(n247039));
   no02f02 U262778 (.o(n247042),
	.a(regtop_g_seqstrt_r),
	.b(n246922));
   na02s01 U262779 (.o(n246952),
	.a(regtop_g_udb0_r[0]),
	.b(regtop_g_udb0_r[1]));
   in01f01 U262780 (.o(n246954),
	.a(n247042));
   na02f01 U262781 (.o(n246935),
	.a(n246871),
	.b(n246868));
   in01s01 U262782 (.o(n246848),
	.a(n246847));
   in01f01 U262783 (.o(n246062),
	.a(regtop_g_udb2_r[0]));
   na02f01 U262784 (.o(n246850),
	.a(n252462),
	.b(n246849));
   na02s02 U262785 (.o(n247050),
	.a(n246956),
	.b(n246928));
   na02f02 U262786 (.o(n247051),
	.a(n247045),
	.b(n247044));
   na02s02 U262787 (.o(n247044),
	.a(n247053),
	.b(n247050));
   no02f04 U262788 (.o(n247053),
	.a(regtop_g_seqstrt_r),
	.b(n246930));
   in01f01 U262789 (.o(n246963),
	.a(n247053));
   na02f04 U262790 (.o(n252521),
	.a(n252523),
	.b(n252706));
   na02f04 U262791 (.o(n252575),
	.a(regtop_g_paramadr_r[1]),
	.b(n246607));
   na02f01 U262792 (.o(n252630),
	.a(n252711),
	.b(n252613));
   no02f02 U262793 (.o(n252680),
	.a(n245546),
	.b(n245545));
   in01f01 U262794 (.o(n252485),
	.a(n252824));
   na02f02 U262795 (.o(n252704),
	.a(n252731),
	.b(FE_OFN45_n252700));
   na02f02 U262796 (.o(n252752),
	.a(n245547),
	.b(n246609));
   na02f03 U262797 (.o(n249079),
	.a(n249137),
	.b(FE_OFN6_n246618));
   in01f04 U262798 (.o(n252660),
	.a(regtop_g_paramdata_r[19]));
   in01f04 U262799 (.o(n252662),
	.a(regtop_g_paramdata_r[20]));
   in01f04 U262800 (.o(n252666),
	.a(regtop_g_paramdata_r[22]));
   in01f04 U262801 (.o(n252778),
	.a(regtop_g_paramdata_r[23]));
   no02f01 U262802 (.o(n246618),
	.a(n246614),
	.b(n246613));
   ao22s01 U262804 (.o(n245935),
	.a(n246658),
	.b(n246543),
	.c(n246664),
	.d(n246492));
   na02f02 U262805 (.o(n247000),
	.a(n246890),
	.b(n247020));
   ao12s02 U262806 (.o(n246025),
	.a(n246023),
	.b(n246309),
	.c(n246024));
   no03f01 U262807 (.o(n246024),
	.a(n246303),
	.b(n246302),
	.c(n246670));
   ao12f01 U262808 (.o(n249018),
	.a(n249012),
	.b(n249014),
	.c(n249013));
   oa12s01 U262809 (.o(n249013),
	.a(n249009),
	.b(n249011),
	.c(n249010));
   na02s01 U262810 (.o(n246370),
	.a(FE_OFN2_g_swrst_r_n),
	.b(y1_bs_wait_n));
   ao12f02 U262811 (.o(n247031),
	.a(n246977),
	.b(n246979),
	.c(n246978));
   ao12f01 U262812 (.o(n246834),
	.a(n246829),
	.b(n246831),
	.c(n246830));
   in01s01 U262813 (.o(n247148),
	.a(n247147));
   na02s02 U262814 (.o(n246836),
	.a(n246964),
	.b(vldtop_vld_syndec_vld_vlfeed_feed_on));
   na02f06 U262815 (.o(n252377),
	.a(regtop_g_wd_r[0]),
	.b(n252871));
   in01f01 U262816 (.o(n252957),
	.a(n252954));
   na04f01 U262817 (.o(n248267),
	.a(n248256),
	.b(n248255),
	.c(n248254),
	.d(n248253));
   na04f03 U262818 (.o(n248265),
	.a(n248264),
	.b(n248263),
	.c(n248262),
	.d(n248261));
   na04f06 U262819 (.o(n248266),
	.a(n248260),
	.b(n248259),
	.c(n248258),
	.d(n248257));
   na04f04 U262820 (.o(n248268),
	.a(n248252),
	.b(n248251),
	.c(n248250),
	.d(n248249));
   na04f03 U262821 (.o(n247436),
	.a(n247429),
	.b(n247428),
	.c(n247427),
	.d(n247426));
   na04f04 U262822 (.o(n248420),
	.a(n248419),
	.b(n248418),
	.c(n248417),
	.d(n248416));
   na04f01 U262823 (.o(n248422),
	.a(n248403),
	.b(n248402),
	.c(n248401),
	.d(n248400));
   na04f06 U262824 (.o(n247840),
	.a(n247839),
	.b(n247838),
	.c(n247837),
	.d(n247836));
   na04f04 U262825 (.o(n247841),
	.a(n247835),
	.b(n247834),
	.c(n247833),
	.d(n247832));
   na04s02 U262826 (.o(n247843),
	.a(n247827),
	.b(n247826),
	.c(n247825),
	.d(n247824));
   na04f01 U262827 (.o(n247842),
	.a(n247831),
	.b(n247830),
	.c(n247829),
	.d(n247828));
   na04f06 U262828 (.o(n248894),
	.a(n248893),
	.b(n248892),
	.c(n248891),
	.d(n248890));
   na04f06 U262829 (.o(n248895),
	.a(n248881),
	.b(n248880),
	.c(n248879),
	.d(n248878));
   na04f01 U262830 (.o(n248897),
	.a(n248857),
	.b(n248856),
	.c(n248855),
	.d(n248854));
   na04f02 U262831 (.o(n247988),
	.a(n247977),
	.b(n247976),
	.c(n247975),
	.d(n247974));
   na04f01 U262832 (.o(n247986),
	.a(n247985),
	.b(n247984),
	.c(n247983),
	.d(n247982));
   na04f03 U262833 (.o(n247987),
	.a(n247981),
	.b(n247980),
	.c(n247979),
	.d(n247978));
   na04f04 U262834 (.o(n247989),
	.a(n247973),
	.b(n247972),
	.c(n247971),
	.d(n247970));
   na04f04 U262835 (.o(n247966),
	.a(n247965),
	.b(n247964),
	.c(n247963),
	.d(n247962));
   na04f04 U262836 (.o(n247967),
	.a(n247961),
	.b(n247960),
	.c(n247959),
	.d(n247958));
   na04f01 U262837 (.o(n247969),
	.a(n247953),
	.b(n247952),
	.c(n247951),
	.d(n247950));
   na04f03 U262838 (.o(n247694),
	.a(n247670),
	.b(n247669),
	.c(n247668),
	.d(n247667));
   na04f02 U262839 (.o(n247692),
	.a(n247691),
	.b(n247690),
	.c(n247689),
	.d(n247688));
   na04f03 U262840 (.o(n247693),
	.a(n247681),
	.b(n247680),
	.c(n247679),
	.d(n247678));
   na04f01 U262841 (.o(n247695),
	.a(n247659),
	.b(n247658),
	.c(n247657),
	.d(n247656));
   na04f04 U262842 (.o(n247736),
	.a(n247725),
	.b(n247724),
	.c(n247723),
	.d(n247722));
   na04f02 U262843 (.o(n247734),
	.a(n247733),
	.b(n247732),
	.c(n247731),
	.d(n247730));
   na04f02 U262844 (.o(n247735),
	.a(n247729),
	.b(n247728),
	.c(n247727),
	.d(n247726));
   na04f02 U262845 (.o(n247737),
	.a(n247721),
	.b(n247720),
	.c(n247719),
	.d(n247718));
   na04f03 U262846 (.o(n247714),
	.a(n247713),
	.b(n247712),
	.c(n247711),
	.d(n247710));
   na04f01 U262847 (.o(n247717),
	.a(n247701),
	.b(n247700),
	.c(n247699),
	.d(n247698));
   na04f01 U262848 (.o(n247778),
	.a(n247767),
	.b(n247766),
	.c(n247765),
	.d(n247764));
   na04f01 U262849 (.o(n247776),
	.a(n247775),
	.b(n247774),
	.c(n247773),
	.d(n247772));
   na04s02 U262850 (.o(n247777),
	.a(n247771),
	.b(n247770),
	.c(n247769),
	.d(n247768));
   na04f03 U262851 (.o(n247779),
	.a(n247763),
	.b(n247762),
	.c(n247761),
	.d(n247760));
   na04f03 U262852 (.o(n247820),
	.a(n247809),
	.b(n247808),
	.c(n247807),
	.d(n247806));
   na04f02 U262853 (.o(n247818),
	.a(n247817),
	.b(n247816),
	.c(n247815),
	.d(n247814));
   na04f06 U262854 (.o(n247819),
	.a(n247813),
	.b(n247812),
	.c(n247811),
	.d(n247810));
   na04f04 U262855 (.o(n247821),
	.a(n247805),
	.b(n247804),
	.c(n247803),
	.d(n247802));
   ao22s01 U262856 (.o(n247874),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2030]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1006]));
   na04f02 U262857 (.o(n247946),
	.a(n247935),
	.b(n247934),
	.c(n247933),
	.d(n247932));
   na04f03 U262858 (.o(n247944),
	.a(n247943),
	.b(n247942),
	.c(n247941),
	.d(n247940));
   ao22s01 U262859 (.o(n247943),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1037]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[13]));
   na04f04 U262860 (.o(n247945),
	.a(n247939),
	.b(n247938),
	.c(n247937),
	.d(n247936));
   na04f04 U262861 (.o(n247947),
	.a(n247931),
	.b(n247930),
	.c(n247929),
	.d(n247928));
   na04f04 U262862 (.o(n247924),
	.a(n247923),
	.b(n247922),
	.c(n247921),
	.d(n247920));
   ao22s01 U262863 (.o(n247922),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1581]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[557]));
   na04f01 U262864 (.o(n247927),
	.a(n247911),
	.b(n247910),
	.c(n247909),
	.d(n247908));
   ao22s01 U262865 (.o(n248429),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1132]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[108]));
   na04f03 U262866 (.o(n248444),
	.a(n248433),
	.b(n248432),
	.c(n248431),
	.d(n248430));
   na04f01 U262867 (.o(n248442),
	.a(n248441),
	.b(n248440),
	.c(n248439),
	.d(n248438));
   ao22s01 U262868 (.o(n248438),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1836]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[812]));
   na04f01 U262869 (.o(n248072),
	.a(n248061),
	.b(n248060),
	.c(n248059),
	.d(n248058));
   na04f02 U262870 (.o(n248070),
	.a(n248069),
	.b(n248068),
	.c(n248067),
	.d(n248066));
   na04f04 U262871 (.o(n248071),
	.a(n248065),
	.b(n248064),
	.c(n248063),
	.d(n248062));
   na04f03 U262872 (.o(n248073),
	.a(n248057),
	.b(n248056),
	.c(n248055),
	.d(n248054));
   ao22s01 U262873 (.o(n248056),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1611]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[587]));
   na04f02 U262874 (.o(n248050),
	.a(n248049),
	.b(n248048),
	.c(n248047),
	.d(n248046));
   na04f04 U262875 (.o(n248092),
	.a(n248091),
	.b(n248090),
	.c(n248089),
	.d(n248088));
   na04f02 U262876 (.o(n248094),
	.a(n248083),
	.b(n248082),
	.c(n248081),
	.d(n248080));
   ao22s01 U262877 (.o(n248083),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1194]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[170]));
   na04f06 U262878 (.o(n248714),
	.a(n248713),
	.b(n248712),
	.c(n248711),
	.d(n248710));
   na04f06 U262879 (.o(n248715),
	.a(n248709),
	.b(n248708),
	.c(n248707),
	.d(n248706));
   na04f03 U262880 (.o(n248716),
	.a(n248705),
	.b(n248704),
	.c(n248703),
	.d(n248702));
   ao22s01 U262881 (.o(n248704),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1673]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[649]));
   na04f06 U262882 (.o(n248717),
	.a(n248701),
	.b(n248700),
	.c(n248699),
	.d(n248698));
   na04f02 U262883 (.o(n248694),
	.a(n248693),
	.b(n248692),
	.c(n248691),
	.d(n248690));
   na04f04 U262884 (.o(n248736),
	.a(n248735),
	.b(n248734),
	.c(n248733),
	.d(n248732));
   ao22s01 U262885 (.o(n248731),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1256]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[232]));
   na04f03 U262886 (.o(n248738),
	.a(n248727),
	.b(n248726),
	.c(n248725),
	.d(n248724));
   ao22s01 U262887 (.o(n248790),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1990]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[966]));
   na04f06 U262888 (.o(n248778),
	.a(n248777),
	.b(n248776),
	.c(n248775),
	.d(n248774));
   ao22s01 U262889 (.o(n248777),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1062]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[38]));
   na04f02 U262890 (.o(n248590),
	.a(n248579),
	.b(n248578),
	.c(n248577),
	.d(n248576));
   na04f02 U262891 (.o(n248589),
	.a(n248583),
	.b(n248582),
	.c(n248581),
	.d(n248580));
   na04f03 U262892 (.o(n248591),
	.a(n248575),
	.b(n248574),
	.c(n248573),
	.d(n248572));
   ao22s01 U262893 (.o(n248575),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1092]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[68]));
   na04f02 U262894 (.o(n248588),
	.a(n248587),
	.b(n248586),
	.c(n248585),
	.d(n248584));
   ao22s01 U262895 (.o(n248584),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1796]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[772]));
   na04f03 U262896 (.o(n248568),
	.a(n248567),
	.b(n248566),
	.c(n248565),
	.d(n248564));
   ao22s01 U262897 (.o(n248554),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1636]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[612]));
   na04f03 U262898 (.o(n248548),
	.a(n248537),
	.b(n248536),
	.c(n248535),
	.d(n248534));
   na04f02 U262899 (.o(n248546),
	.a(n248545),
	.b(n248544),
	.c(n248543),
	.d(n248542));
   na04f04 U262900 (.o(n248547),
	.a(n248541),
	.b(n248540),
	.c(n248539),
	.d(n248538));
   na04f02 U262901 (.o(n248549),
	.a(n248533),
	.b(n248532),
	.c(n248531),
	.d(n248530));
   ao22s01 U262902 (.o(n247998),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1698]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[674]));
   na04f01 U262903 (.o(n248030),
	.a(n248019),
	.b(n248018),
	.c(n248017),
	.d(n248016));
   ao22s01 U262904 (.o(n248019),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1154]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[130]));
   na04f02 U262905 (.o(n248028),
	.a(n248027),
	.b(n248026),
	.c(n248025),
	.d(n248024));
   na04f06 U262906 (.o(n248029),
	.a(n248023),
	.b(n248022),
	.c(n248021),
	.d(n248020));
   na04f03 U262907 (.o(n248031),
	.a(n248015),
	.b(n248014),
	.c(n248013),
	.d(n248012));
   na04f04 U262908 (.o(n248008),
	.a(n248007),
	.b(n248006),
	.c(n248005),
	.d(n248004));
   na04f03 U262909 (.o(n248632),
	.a(n248621),
	.b(n248620),
	.c(n248619),
	.d(n248618));
   na04f02 U262910 (.o(n248630),
	.a(n248629),
	.b(n248628),
	.c(n248627),
	.d(n248626));
   na04f04 U262911 (.o(n248631),
	.a(n248625),
	.b(n248624),
	.c(n248623),
	.d(n248622));
   na04f06 U262912 (.o(n248633),
	.a(n248617),
	.b(n248616),
	.c(n248615),
	.d(n248614));
   na04f04 U262913 (.o(n248225),
	.a(n248214),
	.b(n248213),
	.c(n248212),
	.d(n248211));
   na04f03 U262914 (.o(n248223),
	.a(n248222),
	.b(n248221),
	.c(n248220),
	.d(n248219));
   na04f04 U262915 (.o(n248224),
	.a(n248218),
	.b(n248217),
	.c(n248216),
	.d(n248215));
   ao22s01 U262916 (.o(n248218),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1216]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[192]));
   na04f06 U262917 (.o(n248226),
	.a(n248210),
	.b(n248209),
	.c(n248208),
	.d(n248207));
   oa12s01 U262918 (.o(n245670),
	.a(n245703),
	.b(n245705),
	.c(n245702));
   ao12f02 U262919 (.o(n245705),
	.a(n245665),
	.b(n245729),
	.c(n245666));
   na02f02 U262920 (.o(n246097),
	.a(n246095),
	.b(n246112));
   na02f02 U262921 (.o(n246096),
	.a(regtop_g_udb2_r[4]),
	.b(n246112));
   in01f01 U262922 (.o(n246099),
	.a(n246092));
   in01s01 U262923 (.o(n246091),
	.a(n246088));
   in01f01 U262924 (.o(n246090),
	.a(n246089));
   na02f03 U262925 (.o(n246073),
	.a(regtop_g_udb1_r[1]),
	.b(regtop_g_udb0_r[1]));
   na02f02 U262926 (.o(n246120),
	.a(n246118),
	.b(n246124));
   in01f01 U262927 (.o(n246122),
	.a(n246115));
   no02f02 U262928 (.o(n246115),
	.a(n246114),
	.b(n246113));
   in01f01 U262929 (.o(n246113),
	.a(n246112));
   no02f01 U262930 (.o(n246080),
	.a(n246079),
	.b(n246078));
   in01f01 U262931 (.o(n246078),
	.a(n246077));
   na02f02 U262932 (.o(n246106),
	.a(n246099),
	.b(n246098));
   in01f01 U262933 (.o(n245452),
	.a(n245492));
   na02f01 U262934 (.o(n246134),
	.a(n246132),
	.b(n246131));
   na02f01 U262935 (.o(n246132),
	.a(regtop_g_udb1_r[6]),
	.b(n246129));
   na02f01 U262936 (.o(n246131),
	.a(n246130),
	.b(n246129));
   na02f01 U262937 (.o(n246129),
	.a(regtop_g_udb1_r[6]),
	.b(n246130));
   in01f01 U262938 (.o(n246135),
	.a(n246127));
   no02f01 U262939 (.o(n246127),
	.a(n246126),
	.b(n246125));
   in01s01 U262940 (.o(n246100),
	.a(n246107));
   na03f01 U262941 (.o(n246730),
	.a(vldtop_vld_syndec_vld_vscdet_v_search_1st_r),
	.b(n246729),
	.c(n248999));
   no02f01 U262942 (.o(n246733),
	.a(n246732),
	.b(vldtop_vld_syndec_vld_seqhed_pre_SHIFT[3]));
   no02f80 U262944 (.o(n245406),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[25]),
	.b(g_field_start_add_r[25]));
   no02f02 U262945 (.o(n245342),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[16]),
	.b(g_field_start_add_r[16]));
   no02f02 U262946 (.o(n245341),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[15]),
	.b(g_field_start_add_r[15]));
   no02f02 U262947 (.o(n245336),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[14]),
	.b(g_field_start_add_r[14]));
   no02f02 U262948 (.o(n245335),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[13]),
	.b(g_field_start_add_r[13]));
   no02f03 U262949 (.o(n245324),
	.a(g_field_start_add_r[11]),
	.b(g_field_start_add_r[12]));
   no02f01 U262950 (.o(n245828),
	.a(vh_1_ph_add[2]),
	.b(vh_1_ph_add[28]));
   ao22f02 U262951 (.o(n245465),
	.a(regtop_g_brv_r[16]),
	.b(FE_OFN546_n245460),
	.c(regtop_g_tr_r[0]),
	.d(FE_OFN552_n245462));
   ao22f02 U262952 (.o(n245464),
	.a(regtop_g_fcho2_r[0]),
	.b(FE_OFN527_n249828),
	.c(regtop_g_cp_r[0]),
	.d(n249813));
   ao22f01 U262953 (.o(n249773),
	.a(n249824),
	.b(regtop_g_dhs_r[8]),
	.c(n249823),
	.d(regtop_g_hsv_r[8]));
   ao22f01 U262954 (.o(n249772),
	.a(FE_OFN546_n245460),
	.b(regtop_g_frc_r[0]),
	.c(FE_OFN552_n245462),
	.d(regtop_g_tr_r[8]));
   ao22s01 U262955 (.o(n249775),
	.a(FE_OFN527_n249828),
	.b(regtop_g_fcho2_r[8]),
	.c(n249813),
	.d(regtop_g_cd_r));
   na02f06 U262956 (.o(n245471),
	.a(regtop_g_a_r[3]),
	.b(FE_OFN534_regtop_g_a_r_5_));
   na02f04 U262957 (.o(n245461),
	.a(n245450),
	.b(n245449));
   in01f02 U262958 (.o(n247060),
	.a(regtop_v1_hdi00_a[3]));
   in01f01 U262959 (.o(n250164),
	.a(regtop_v1_hdi00_a[1]));
   no02f03 U262960 (.o(n247055),
	.a(regtop_v1_hdi00_a[3]),
	.b(regtop_v1_hdi00_a[4]));
   in01f03 U262961 (.o(n247056),
	.a(regtop_v1_hdi00_a[5]));
   na02f01 U262962 (.o(n246136),
	.a(n246135),
	.b(n246134));
   in01f01 U262963 (.o(n246137),
	.a(n246133));
   no02f01 U262964 (.o(n246133),
	.a(n246135),
	.b(n246134));
   na02f02 U262965 (.o(n246176),
	.a(n246175),
	.b(n246174));
   ao12f02 U262966 (.o(n246178),
	.a(n246067),
	.b(n246163),
	.c(n246160));
   no02f01 U262967 (.o(n249109),
	.a(n245772),
	.b(n252254));
   in01s01 U262968 (.o(n252275),
	.a(n249648));
   oa12s01 U262969 (.o(n246899),
	.a(regtop_g_paramadr_r[7]),
	.b(regtop_g_paramadr_r[5]),
	.c(n245514));
   oa12f01 U262970 (.o(n246163),
	.a(n246167),
	.b(n246166),
	.c(n246062));
   in01f01 U262971 (.o(n246653),
	.a(n246714));
   na02s01 U262972 (.o(n246445),
	.a(n246670),
	.b(n246444));
   oa22s01 U262973 (.o(n246452),
	.a(n246466),
	.b(n246463),
	.c(n246464),
	.d(n246467));
   oa22s01 U262974 (.o(n246451),
	.a(n246468),
	.b(n246485),
	.c(n246450),
	.d(n246484));
   in01f01 U262975 (.o(n245529),
	.a(n246608));
   na03s02 U262976 (.o(n247004),
	.a(n247003),
	.b(n247018),
	.c(n247002));
   ao12f02 U262977 (.o(n246781),
	.a(n246778),
	.b(n246795),
	.c(n246779));
   oa12s02 U262978 (.o(n246734),
	.a(n246733),
	.b(n246782),
	.c(n246799));
   in01s01 U262979 (.o(n246801),
	.a(n246797));
   na02f06 U262980 (.o(n246372),
	.a(regtop_g_a_r[3]),
	.b(regtop_g_a_r[5]));
   na03f08 U262981 (.o(n247109),
	.a(regtop_v1_hdi00_a[2]),
	.b(regtop_v1_hdi00_a[1]),
	.c(FE_OFN516_regtop_v1_hdi00_a_0_));
   no02f04 U262982 (.o(n245416),
	.a(n245415),
	.b(n245414));
   no02s01 U262983 (.o(n245408),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[26]),
	.b(n245413));
   no02f01 U262984 (.o(n245386),
	.a(n245384),
	.b(n245383));
   no02s01 U262985 (.o(n245377),
	.a(g_field_start_add_r[21]),
	.b(n245382));
   no02f01 U262986 (.o(n245370),
	.a(n245358),
	.b(n245357));
   no02f01 U262987 (.o(n245367),
	.a(n245363),
	.b(n245362));
   no02f01 U262988 (.o(n245363),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[18]),
	.b(n245361));
   no02f01 U262989 (.o(n245362),
	.a(g_field_start_add_r[18]),
	.b(n245361));
   oa12f02 U262990 (.o(n245353),
	.a(n245668),
	.b(n245667),
	.c(n245703));
   no02f01 U262991 (.o(n245344),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[16]),
	.b(n245342));
   no02f02 U262992 (.o(n245345),
	.a(n245338),
	.b(n245337));
   no02f02 U262993 (.o(n245338),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[14]),
	.b(n245336));
   no02f02 U262994 (.o(n245337),
	.a(g_field_start_add_r[14]),
	.b(n245336));
   no02f01 U262995 (.o(n245710),
	.a(n245346),
	.b(n245345));
   no02f01 U262996 (.o(n245330),
	.a(n245323),
	.b(n245322));
   no02f01 U262997 (.o(n245323),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[13]),
	.b(n245335));
   no02f01 U262998 (.o(n245322),
	.a(g_field_start_add_r[13]),
	.b(n245335));
   no02f01 U262999 (.o(n245326),
	.a(g_field_start_add_r[11]),
	.b(n245324));
   no02f01 U263000 (.o(n245325),
	.a(g_field_start_add_r[12]),
	.b(n245324));
   ao12s01 U263001 (.o(n245868),
	.a(n245866),
	.b(n245899),
	.c(n245867));
   ao12s01 U263002 (.o(n245900),
	.a(n245897),
	.b(n245899),
	.c(n245898));
   ao12s01 U263003 (.o(n245888),
	.a(n245886),
	.b(n245899),
	.c(n245887));
   no02s01 U263004 (.o(n245856),
	.a(vh_1_ph_add[5]),
	.b(vh_1_ph_add[31]));
   oa12s01 U263005 (.o(n245821),
	.a(n245831),
	.b(n245830),
	.c(n245827));
   no02s01 U263006 (.o(n245830),
	.a(vh_1_ph_add[3]),
	.b(vh_1_ph_add[29]));
   oa12s01 U263007 (.o(n245823),
	.a(n245810),
	.b(n245812),
	.c(n245811));
   no02s01 U263008 (.o(n249902),
	.a(n249910),
	.b(n249903));
   na02s01 U263009 (.o(n249910),
	.a(vh_1_ph_add[0]),
	.b(vh_1_ph_add[1]));
   na03f01 U263010 (.o(n245552),
	.a(n252673),
	.b(n252487),
	.c(n252820));
   no02f01 U263011 (.o(n249778),
	.a(n249777),
	.b(n249776));
   oa12s01 U263012 (.o(n249777),
	.a(n249770),
	.b(n249771),
	.c(n252828));
   ao22s01 U263013 (.o(n249770),
	.a(n249769),
	.b(regtop_g_ps_r),
	.c(n249811),
	.d(g_pcut_r[8]));
   na04f06 U263014 (.o(n245503),
	.a(n245502),
	.b(n245501),
	.c(n245500),
	.d(n245499));
   no02f02 U263015 (.o(n249728),
	.a(n245444),
	.b(n249588));
   no02f02 U263016 (.o(n249729),
	.a(n245444),
	.b(n252275));
   ao22s01 U263017 (.o(n249748),
	.a(n249811),
	.b(g_mbc_r[0]),
	.c(n249744),
	.d(regtop_g_fbst_r[0]));
   ao22f01 U263018 (.o(n249740),
	.a(n249813),
	.b(regtop_g_mc_r[0]),
	.c(n249824),
	.d(regtop_g_dvs_r[0]));
   ao22f04 U263019 (.o(n249743),
	.a(n249823),
	.b(regtop_g_vsv_r[0]),
	.c(n249812),
	.d(regtop_g_tmc_r[0]));
   ao12f01 U263020 (.o(n249929),
	.a(FE_OFN493_n252377),
	.b(n252309),
	.c(n249925));
   no02f06 U263021 (.o(n249769),
	.a(n245491),
	.b(n245470));
   na02f02 U263022 (.o(n246158),
	.a(n246154),
	.b(n246155));
   na02f02 U263023 (.o(n246157),
	.a(n246156),
	.b(n246155));
   na02f06 U263024 (.o(n249039),
	.a(n248992),
	.b(n248994));
   no02f01 U263025 (.o(n246194),
	.a(regtop_g_paramadr_r[2]),
	.b(n246608));
   na02f01 U263026 (.o(n246943),
	.a(regtop_g_paramadr_r[0]),
	.b(regtop_g_paramadr_r[1]));
   na02f01 U263027 (.o(n245545),
	.a(regtop_g_paramadr_r[4]),
	.b(n245763));
   na02f03 U263028 (.o(n245763),
	.a(n245544),
	.b(n252517));
   no02f01 U263029 (.o(n245547),
	.a(regtop_g_paramadr_r[7]),
	.b(n252449));
   no02f02 U263030 (.o(n252775),
	.a(regtop_g_paramadr_r[7]),
	.b(n252314));
   in01f01 U263031 (.o(n252776),
	.a(n252757));
   in01f03 U263032 (.o(n246609),
	.a(regtop_g_paramadr_r[5]));
   ao22f01 U263033 (.o(n245934),
	.a(n246706),
	.b(n246377),
	.c(n246653),
	.d(n246546));
   oa22s01 U263034 (.o(n246537),
	.a(n246536),
	.b(n246711),
	.c(n246535),
	.d(n246714));
   oa22s01 U263035 (.o(n246538),
	.a(n246534),
	.b(n246578),
	.c(n246533),
	.d(n246708));
   ao22s01 U263036 (.o(n246306),
	.a(n246512),
	.b(n246698),
	.c(n246511),
	.d(n246694));
   in01s01 U263037 (.o(n246455),
	.a(n246449));
   in01s01 U263038 (.o(n246454),
	.a(n246453));
   ao22s01 U263039 (.o(n246425),
	.a(n246512),
	.b(n246526),
	.c(n246511),
	.d(n246482));
   oa22s01 U263040 (.o(n246423),
	.a(n246485),
	.b(n246483),
	.c(n246484),
	.d(n246422));
   in01s01 U263041 (.o(n252234),
	.a(n245939));
   oa22s01 U263042 (.o(n246020),
	.a(n246709),
	.b(n246711),
	.c(n246394),
	.d(n246714));
   oa22s01 U263043 (.o(n246021),
	.a(n246651),
	.b(n246708),
	.c(n246715),
	.d(n246578));
   no02s02 U263044 (.o(n246728),
	.a(vldtop_vld_syndec_vld_vscdet_v_search_1st_r),
	.b(n249011));
   in01s01 U263045 (.o(n249012),
	.a(n249061));
   na02s01 U263046 (.o(n249008),
	.a(n249007),
	.b(n249006));
   no04s02 U263047 (.o(n249006),
	.a(vldtop_vld_syndec_UREG[8]),
	.b(vldtop_vld_syndec_UREG[3]),
	.c(n249005),
	.d(n249004));
   na04f01 U263048 (.o(n249004),
	.a(vldtop_vld_syndec_UREG[0]),
	.b(n249003),
	.c(n249002),
	.d(n249001));
   no02f03 U263049 (.o(n249011),
	.a(vldtop_vld_syndec_vld_vscdet_v_search_1st_r),
	.b(n246727));
   na02f01 U263050 (.o(n246725),
	.a(vldtop_vld_syndec_UREG[24]),
	.b(vldtop_vld_syndec_vld_vscdet_v_detvald_r[1]));
   na02s01 U263051 (.o(n249015),
	.a(n246361),
	.b(n246731));
   no04f02 U263052 (.o(n249003),
	.a(vldtop_vld_syndec_UREG[1]),
	.b(vldtop_vld_syndec_UREG[2]),
	.c(vldtop_vld_syndec_UREG[4]),
	.d(vldtop_vld_syndec_UREG[5]));
   na02f04 U263053 (.o(n246828),
	.a(vldtop_vld_syndec_ADP[3]),
	.b(n246738));
   in01s01 U263054 (.o(n246364),
	.a(n246363));
   no02f01 U263056 (.o(n245604),
	.a(n245429),
	.b(n245428));
   na02f01 U263057 (.o(n245657),
	.a(n245387),
	.b(n245386));
   in01s01 U263058 (.o(n245658),
	.a(n245385));
   no02f03 U263059 (.o(n245694),
	.a(n245381),
	.b(n245380));
   na02s02 U263060 (.o(n245695),
	.a(n245381),
	.b(n245380));
   no02f01 U263061 (.o(n245686),
	.a(n245368),
	.b(n245367));
   na02f01 U263062 (.o(n245720),
	.a(n245368),
	.b(n245367));
   no02f02 U263063 (.o(n245667),
	.a(n245352),
	.b(n245351));
   na02f02 U263064 (.o(n245727),
	.a(n245346),
	.b(n245345));
   na02f01 U263065 (.o(n245736),
	.a(n245330),
	.b(n245329));
   no02f02 U263066 (.o(n245735),
	.a(n245330),
	.b(n245329));
   na02f02 U263067 (.o(n245744),
	.a(n245328),
	.b(busrtop_b_rreq_N229));
   no02m02 U263068 (.o(n245743),
	.a(n245328),
	.b(busrtop_b_rreq_N229));
   no04f03 U263069 (.o(n249319),
	.a(y1_bs_data_r[3]),
	.b(y1_bs_data_r[5]),
	.c(y1_bs_data_r[28]),
	.d(y1_bs_data_r[30]));
   ao12s01 U263071 (.o(n246229),
	.a(n246213),
	.b(n246214),
	.c(n246215));
   na02f01 U263072 (.o(n249282),
	.a(n249257),
	.b(n249287));
   no02f80 U263073 (.o(n249287),
	.a(busrtop_b_rreq_vrh_add1_r[0]),
	.b(busrtop_b_rreq_vrh_add1_r[1]));
   ao22f01 U263075 (.o(n249044),
	.a(n249042),
	.b(n249066),
	.c(regtop_g_adb_r[6]),
	.d(n249041));
   na02f02 U263077 (.o(n249056),
	.a(n249052),
	.b(n249053));
   in01f03 U263079 (.o(n248994),
	.a(n248991));
   in01s01 U263080 (.o(n249216),
	.a(n249215));
   oa12f01 U263081 (.o(n249215),
	.a(n249214),
	.b(n252656),
	.c(n249247));
   ao22f01 U263083 (.o(n249142),
	.a(n249211),
	.b(regtop_g_paramdata_r[12]),
	.c(FE_OFN496_n249242),
	.d(regtop_g_paramdata_r[14]));
   in01s01 U263084 (.o(n249230),
	.a(n249229));
   oa12f01 U263085 (.o(n249229),
	.a(n249228),
	.b(n252660),
	.c(n249247));
   ao12f01 U263086 (.o(n249228),
	.a(n249227),
	.b(FE_OFN551_n249140),
	.c(regtop_g_atscd_r[10]));
   oa22f01 U263087 (.o(n249227),
	.a(FE_OFN483_n249211),
	.b(n252648),
	.c(n249242),
	.d(n252652));
   in01s01 U263088 (.o(n249237),
	.a(n249236));
   oa12s01 U263089 (.o(n249236),
	.a(n249235),
	.b(n252662),
	.c(n249247));
   ao12f01 U263090 (.o(n249235),
	.a(n249234),
	.b(FE_OFN551_n249140),
	.c(regtop_g_atscd_r[11]));
   oa22f01 U263091 (.o(n249234),
	.a(FE_OFN483_n249211),
	.b(n252650),
	.c(n249242),
	.d(n252654));
   in01s01 U263092 (.o(n249249),
	.a(n249248));
   oa12f01 U263093 (.o(n249248),
	.a(n249246),
	.b(n252664),
	.c(n249247));
   ao12f01 U263094 (.o(n249246),
	.a(n249244),
	.b(FE_OFN551_n249140),
	.c(regtop_g_atscd_r[12]));
   oa22f01 U263095 (.o(n249244),
	.a(FE_OFN483_n249211),
	.b(n252652),
	.c(n249242),
	.d(n252656));
   in01s01 U263096 (.o(n249223),
	.a(n249222));
   oa12f01 U263097 (.o(n249222),
	.a(n249221),
	.b(n252778),
	.c(n249247));
   ao12f01 U263098 (.o(n249221),
	.a(n249220),
	.b(FE_OFN551_n249140),
	.c(regtop_g_atscd_r[14]));
   oa22f01 U263099 (.o(n249220),
	.a(FE_OFN483_n249211),
	.b(n252656),
	.c(n249242),
	.d(n252660));
   in01s01 U263100 (.o(n249206),
	.a(n249205));
   oa12f01 U263101 (.o(n249205),
	.a(n249204),
	.b(n252755),
	.c(n249247));
   ao12f01 U263102 (.o(n249204),
	.a(n249203),
	.b(FE_OFN551_n249140),
	.c(regtop_g_atscd_r[15]));
   oa22f01 U263103 (.o(n249203),
	.a(FE_OFN483_n249211),
	.b(n252658),
	.c(n249242),
	.d(n252662));
   ao12s01 U263104 (.o(n249091),
	.a(n249089),
	.b(n249127),
	.c(regtop_g_atscd_r[19]));
   oa22s01 U263105 (.o(n249089),
	.a(FE_OFN483_n249211),
	.b(n252666),
	.c(n249242),
	.d(n252755));
   ao12f01 U263106 (.o(n249117),
	.a(n249115),
	.b(n249127),
	.c(regtop_g_atscd_r[16]));
   ao22f01 U263107 (.o(n249114),
	.a(n249113),
	.b(n249112),
	.c(regtop_g_paramdata_r[24]),
	.d(n249210));
   na02f01 U263108 (.o(n245777),
	.a(FE_OFN4_n245443),
	.b(regtop_g_a_r[8]));
   no02f02 U263109 (.o(n252283),
	.a(n252276),
	.b(regtop_g_hclr_r_s));
   in01f01 U263110 (.o(n252285),
	.a(n252276));
   na02f02 U263111 (.o(n252286),
	.a(n245492),
	.b(n245449));
   no04f01 U263112 (.o(n246679),
	.a(n252949),
	.b(n249720),
	.c(n252829),
	.d(n246680));
   no02s01 U263113 (.o(n249925),
	.a(regtop_g_fbst_r[9]),
	.b(n249316));
   no03s01 U263114 (.o(n249314),
	.a(regtop_g_fbst_r[0]),
	.b(regtop_g_fbst_r[3]),
	.c(regtop_g_fbst_r[1]));
   no04s01 U263115 (.o(n249315),
	.a(regtop_g_fbst_r[6]),
	.b(regtop_g_fbst_r[4]),
	.c(regtop_g_fbst_r[7]),
	.d(regtop_g_fbst_r[5]));
   na03f01 U263116 (.o(n252288),
	.a(n252289),
	.b(1'b1),
	.c(n252947));
   no02f01 U263117 (.o(n252245),
	.a(n246865),
	.b(n246864));
   in01s01 U263118 (.o(n252309),
	.a(regtop_g_nfst_r[22]));
   in01f08 U263119 (.o(n252349),
	.a(n252350));
   in01f02 U263120 (.o(n252360),
	.a(n252361));
   no02f01 U263121 (.o(n246266),
	.a(regtop_g_ferror_r),
	.b(FE_OFN486_n245940));
   in01s01 U263122 (.o(n252425),
	.a(n252424));
   na02f01 U263123 (.o(n252483),
	.a(n252687),
	.b(n252464));
   in01s01 U263124 (.o(n252464),
	.a(n252463));
   no02f01 U263125 (.o(n246238),
	.a(n246614),
	.b(n245849));
   in01s01 U263126 (.o(n252758),
	.a(n252564));
   na02f02 U263127 (.o(n252571),
	.a(n252568),
	.b(n252567));
   in01f02 U263128 (.o(n246260),
	.a(FE_OFN220_n246261));
   in01s01 U263129 (.o(n246225),
	.a(n252568));
   in01f01 U263130 (.o(n252591),
	.a(n245944));
   na02s01 U263131 (.o(n245944),
	.a(regtop_g_adb_r[0]),
	.b(regtop_g_adb_r[1]));
   no02f08 U263132 (.o(n252597),
	.a(regtop_g_adb_r[1]),
	.b(n252600));
   no02f02 U263133 (.o(n252706),
	.a(n252517),
	.b(n252516));
   in01f02 U263134 (.o(n252639),
	.a(FE_OFN41_n252640));
   na02f01 U263135 (.o(n252757),
	.a(n252731),
	.b(n252379));
   na02f03 U263136 (.o(n252762),
	.a(n252776),
	.b(n252758));
   in01f02 U263137 (.o(n252772),
	.a(n252773));
   na04f01 U263138 (.o(n246676),
	.a(n246675),
	.b(n246674),
	.c(n246673),
	.d(n246672));
   na02f01 U263139 (.o(n246885),
	.a(n247013),
	.b(n247011));
   na02f01 U263140 (.o(n246884),
	.a(n247012),
	.b(n247010));
   no02s02 U263141 (.o(n245985),
	.a(n245976),
	.b(n245975));
   oa12s02 U263142 (.o(n246055),
	.a(n246053),
	.b(n246417),
	.c(n246054));
   no02f01 U263143 (.o(n246053),
	.a(n246052),
	.b(n246051));
   oa22s01 U263144 (.o(n246052),
	.a(n246042),
	.b(n246708),
	.c(n246533),
	.d(n246711));
   na02s01 U263145 (.o(n246582),
	.a(n246573),
	.b(n246572));
   na02f02 U263146 (.o(n246997),
	.a(n246350),
	.b(n246349));
   na02f02 U263147 (.o(n246998),
	.a(n246442),
	.b(n246441));
   na02f02 U263148 (.o(n246991),
	.a(n246505),
	.b(n246504));
   oa22s01 U263149 (.o(n246493),
	.a(n246714),
	.b(n246576),
	.c(n246711),
	.d(n246577));
   na02s02 U263150 (.o(n246982),
	.a(n246321),
	.b(n246320));
   na04f01 U263151 (.o(n246320),
	.a(n246319),
	.b(vldtop_vld_syndec_ADP[4]),
	.c(n246318),
	.d(n246317));
   no02f01 U263152 (.o(n246321),
	.a(n246314),
	.b(n246313));
   oa12f02 U263153 (.o(n246980),
	.a(n246539),
	.b(n246670),
	.c(n246540));
   no02f01 U263154 (.o(n246539),
	.a(n246538),
	.b(n246537));
   no02s01 U263155 (.o(n246531),
	.a(n246530),
	.b(n246529));
   ao12f02 U263156 (.o(n246994),
	.a(n246519),
	.b(n246520),
	.c(n246670));
   no02f01 U263157 (.o(n246397),
	.a(n246396),
	.b(n246395));
   no02s02 U263158 (.o(n246989),
	.a(n246473),
	.b(n246472));
   ao22s01 U263159 (.o(n246305),
	.a(n246516),
	.b(n246514),
	.c(n246515),
	.d(n246304));
   oa12f02 U263160 (.o(n246987),
	.a(n246410),
	.b(n246412),
	.c(n246411));
   in01s01 U263161 (.o(n246981),
	.a(n246967));
   ao22s01 U263162 (.o(n246276),
	.a(n246516),
	.b(n246304),
	.c(n246515),
	.d(n246275));
   na02f01 U263163 (.o(n248999),
	.a(vldtop_vld_syndec_ADP[3]),
	.b(n246684));
   na02f02 U263164 (.o(n246779),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246729));
   na02f01 U263165 (.o(n249060),
	.a(n249026),
	.b(n249025));
   ao12f02 U263166 (.o(n249063),
	.a(n249019),
	.b(n246897),
	.c(n246896));
   ao22f01 U263167 (.o(n246726),
	.a(vldtop_vld_syndec_vld_vscdet_v_prezerohld_r[1]),
	.b(v1_bs_req_n),
	.c(vldtop_vld_syndec_vld_vscdet_v_prezerotmp_r[1]),
	.d(n246237));
   in01f02 U263168 (.o(n249028),
	.a(n249064));
   na02f02 U263169 (.o(n252942),
	.a(n253015),
	.b(n252912));
   in01f01 U263170 (.o(n252948),
	.a(regtop_g_wd_r[16]));
   na04s02 U263171 (.o(n248842),
	.a(n248831),
	.b(n248830),
	.c(n248829),
	.d(n248828));
   na04f06 U263172 (.o(n248840),
	.a(n248839),
	.b(n248838),
	.c(n248837),
	.d(n248836));
   na04f03 U263173 (.o(n248841),
	.a(n248835),
	.b(n248834),
	.c(n248833),
	.d(n248832));
   na04f02 U263174 (.o(n248843),
	.a(n248827),
	.b(n248826),
	.c(n248825),
	.d(n248824));
   na04f04 U263175 (.o(n248506),
	.a(n248495),
	.b(n248494),
	.c(n248493),
	.d(n248492));
   na04f02 U263176 (.o(n248504),
	.a(n248503),
	.b(n248502),
	.c(n248501),
	.d(n248500));
   na04f02 U263177 (.o(n248505),
	.a(n248499),
	.b(n248498),
	.c(n248497),
	.d(n248496));
   na04f01 U263178 (.o(n248507),
	.a(n248491),
	.b(n248490),
	.c(n248489),
	.d(n248488));
   ao22f01 U263179 (.o(n248481),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1332]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[308]));
   na04f02 U263180 (.o(n248674),
	.a(n248663),
	.b(n248662),
	.c(n248661),
	.d(n248660));
   na04f04 U263181 (.o(n248672),
	.a(n248671),
	.b(n248670),
	.c(n248669),
	.d(n248668));
   na04f04 U263182 (.o(n248673),
	.a(n248667),
	.b(n248666),
	.c(n248665),
	.d(n248664));
   na04f04 U263183 (.o(n248675),
	.a(n248659),
	.b(n248658),
	.c(n248657),
	.d(n248656));
   ao22s01 U263184 (.o(n248649),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1317]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[293]));
   na02s01 U263185 (.o(n245601),
	.a(n245598),
	.b(n245597));
   na02s01 U263186 (.o(n245639),
	.a(n245636),
	.b(n245635));
   oa12m02 U263187 (.o(n245375),
	.a(n245679),
	.b(n245676),
	.c(n245678));
   na02s01 U263188 (.o(n245683),
	.a(n245680),
	.b(n245679));
   oa12s01 U263189 (.o(n245689),
	.a(n245720),
	.b(n245722),
	.c(n245686));
   na02s01 U263190 (.o(n245717),
	.a(n245714),
	.b(n245713));
   na02f02 U263191 (.o(n246000),
	.a(n245999),
	.b(n245998));
   na02s01 U263192 (.o(n245862),
	.a(n245861),
	.b(n245860));
   oa12f02 U263193 (.o(n244972),
	.a(n249523),
	.b(n245444),
	.c(n249524));
   na04s01 U263194 (.o(n249521),
	.a(n249515),
	.b(n249514),
	.c(n249513),
	.d(n249512));
   na03f01 U263195 (.o(n157831),
	.a(n249854),
	.b(n249853),
	.c(n249852));
   in01s01 U263196 (.o(n249853),
	.a(n249849));
   na03f01 U263197 (.o(n157832),
	.a(n249862),
	.b(n249861),
	.c(n249860));
   na02s01 U263198 (.o(n249861),
	.a(n249916),
	.b(n249857));
   na02s01 U263199 (.o(n157833),
	.a(n249869),
	.b(n249868));
   ao12s01 U263200 (.o(n249868),
	.a(n249866),
	.b(n249916),
	.c(n249867));
   na02s01 U263201 (.o(n249876),
	.a(n249916),
	.b(n249872));
   ao12s01 U263202 (.o(n249883),
	.a(n249881),
	.b(n249916),
	.c(n249882));
   na03f01 U263203 (.o(n157836),
	.a(n249892),
	.b(n249891),
	.c(n249890));
   na02s01 U263204 (.o(n249271),
	.a(n249273),
	.b(n249269));
   na02f01 U263205 (.o(n170951),
	.a(n245596),
	.b(n245595));
   na04f02 U263207 (.o(n244220),
	.a(n249785),
	.b(n249784),
	.c(n249783),
	.d(n249782));
   na03f03 U263208 (.o(n244968),
	.a(n249606),
	.b(n249605),
	.c(n249604));
   in01s01 U263209 (.o(n170952),
	.a(n249931));
   na03f06 U263210 (.o(n244967),
	.a(n249626),
	.b(n249625),
	.c(n249624));
   no04f03 U263211 (.o(n249624),
	.a(n249623),
	.b(n249622),
	.c(n249621),
	.d(n249620));
   in01s01 U263212 (.o(n170953),
	.a(n249932));
   na04f02 U263213 (.o(n244213),
	.a(n245513),
	.b(n245512),
	.c(n245511),
	.d(n245510));
   in01s01 U263214 (.o(n170954),
	.a(n249933));
   no04f04 U263215 (.o(n249662),
	.a(n249660),
	.b(n249659),
	.c(n249658),
	.d(n249657));
   in01s01 U263216 (.o(n170955),
	.a(n249934));
   na03f04 U263217 (.o(n244965),
	.a(n249684),
	.b(n249683),
	.c(n249682));
   no04f02 U263218 (.o(n249682),
	.a(n249681),
	.b(n249680),
	.c(n249679),
	.d(n249678));
   in01s01 U263219 (.o(n170956),
	.a(n249935));
   na03f01 U263220 (.o(n244964),
	.a(n249711),
	.b(n249710),
	.c(n249709));
   ao12s01 U263221 (.o(n249711),
	.a(n249687),
	.b(n249746),
	.c(regtop_g_embv_adr_r[1]));
   no04f02 U263222 (.o(n249709),
	.a(n249708),
	.b(n249707),
	.c(n249706),
	.d(n249705));
   in01s01 U263223 (.o(n170957),
	.a(n249936));
   na04s02 U263224 (.o(n244222),
	.a(n249756),
	.b(n249755),
	.c(n249754),
	.d(n249753));
   in01s01 U263225 (.o(n170958),
	.a(n249937));
   in01s01 U263226 (.o(n170959),
	.a(n249938));
   na04s01 U263227 (.o(n249476),
	.a(n249475),
	.b(n249474),
	.c(n249473),
	.d(n249472));
   in01s01 U263228 (.o(n170960),
	.a(n249939));
   na04f04 U263229 (.o(n249488),
	.a(n249487),
	.b(n249486),
	.c(n249485),
	.d(n249484));
   in01s01 U263230 (.o(n170961),
	.a(n249940));
   in01s01 U263231 (.o(n170962),
	.a(n249941));
   in01s01 U263232 (.o(n170963),
	.a(n249942));
   oa12s01 U263233 (.o(n244971),
	.a(n249540),
	.b(n245444),
	.c(n249541));
   in01s01 U263234 (.o(n170964),
	.a(n249943));
   oa12f02 U263235 (.o(n244970),
	.a(n249565),
	.b(n245444),
	.c(n249566));
   no04f02 U263236 (.o(n249566),
	.a(n249564),
	.b(n249563),
	.c(n249562),
	.d(n249561));
   na04f06 U263237 (.o(n249561),
	.a(n249560),
	.b(n249559),
	.c(n249558),
	.d(n249557));
   in01s01 U263238 (.o(n170965),
	.a(n249946));
   ao12f01 U263239 (.o(n249946),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embh_adr_r[0]));
   na04s02 U263240 (.o(n244214),
	.a(FE_OFN466_n249845),
	.b(n249844),
	.c(n249843),
	.d(n249842));
   na04f04 U263241 (.o(n244215),
	.a(n249835),
	.b(n249834),
	.c(n249833),
	.d(n249832));
   na04f03 U263242 (.o(n244217),
	.a(n249810),
	.b(n249809),
	.c(n249808),
	.d(n249807));
   na04f01 U263243 (.o(n244219),
	.a(FE_OFN478_n249800),
	.b(n249799),
	.c(n249798),
	.d(n249797));
   na03f01 U263244 (.o(n244216),
	.a(n249822),
	.b(FE_OFN464_n249821),
	.c(n249820));
   na04f01 U263245 (.o(n249405),
	.a(n249404),
	.b(n249403),
	.c(n249402),
	.d(n249401));
   na04s02 U263246 (.o(n244983),
	.a(n249383),
	.b(n249382),
	.c(n249381),
	.d(n249380));
   na04f01 U263247 (.o(n249429),
	.a(n249428),
	.b(n249427),
	.c(n249426),
	.d(n249425));
   na04s02 U263248 (.o(n244984),
	.a(n249374),
	.b(n249373),
	.c(n249372),
	.d(n249371));
   na04s01 U263249 (.o(n249417),
	.a(n249416),
	.b(n249415),
	.c(n249414),
	.d(n249413));
   oa12f02 U263250 (.o(n244978),
	.a(n249446),
	.b(FE_OFN575_n245444),
	.c(n249447));
   na04f03 U263251 (.o(n249444),
	.a(n249443),
	.b(n249442),
	.c(n249441),
	.d(n249440));
   no04f02 U263252 (.o(n249581),
	.a(n249579),
	.b(n249578),
	.c(n249577),
	.d(n249576));
   ao22s01 U263253 (.o(n246842),
	.a(n252269),
	.b(regtop_g_wd_r[0]),
	.c(regtop_g_issh_r),
	.d(n246841));
   oa22s01 U263254 (.o(n249949),
	.a(n249982),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[511]),
	.d(n249964));
   oa22s01 U263255 (.o(n249950),
	.a(n249982),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[510]),
	.d(FE_OFN268_n249964));
   oa22s01 U263256 (.o(n249951),
	.a(n249982),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[509]),
	.d(FE_OFN268_n249964));
   oa22s01 U263257 (.o(n249952),
	.a(n249982),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[508]),
	.d(FE_OFN268_n249964));
   oa22s01 U263258 (.o(n249953),
	.a(n249982),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[507]),
	.d(FE_OFN268_n249964));
   oa22s01 U263259 (.o(n249955),
	.a(n249982),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[505]),
	.d(FE_OFN268_n249964));
   oa22s01 U263260 (.o(n249956),
	.a(n249982),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[504]),
	.d(FE_OFN268_n249964));
   oa22s01 U263261 (.o(n249957),
	.a(n249982),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[503]),
	.d(FE_OFN268_n249964));
   oa22s01 U263262 (.o(n249958),
	.a(n249982),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[502]),
	.d(FE_OFN268_n249964));
   oa22s01 U263263 (.o(n249959),
	.a(n249982),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[501]),
	.d(FE_OFN268_n249964));
   oa22s01 U263264 (.o(n249960),
	.a(n249982),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[500]),
	.d(FE_OFN268_n249964));
   oa22s01 U263265 (.o(n249961),
	.a(n249982),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[499]),
	.d(FE_OFN268_n249964));
   oa22s01 U263266 (.o(n249962),
	.a(n249982),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[498]),
	.d(FE_OFN268_n249964));
   oa22s01 U263267 (.o(n249963),
	.a(n249982),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[497]),
	.d(FE_OFN268_n249964));
   oa22s01 U263268 (.o(n249965),
	.a(n249982),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[496]),
	.d(FE_OFN268_n249964));
   oa22s01 U263269 (.o(n249966),
	.a(n249982),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[495]),
	.d(FE_OFN268_n249964));
   oa22s01 U263270 (.o(n249967),
	.a(n249982),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[494]),
	.d(FE_OFN268_n249964));
   oa22s01 U263271 (.o(n249968),
	.a(n249982),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[493]),
	.d(FE_OFN268_n249964));
   oa22s01 U263272 (.o(n249969),
	.a(n249982),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[492]),
	.d(FE_OFN268_n249964));
   oa22s01 U263273 (.o(n249971),
	.a(n249982),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[490]),
	.d(FE_OFN268_n249964));
   oa22s01 U263274 (.o(n249972),
	.a(n249982),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[489]),
	.d(n249964));
   oa22s01 U263275 (.o(n249973),
	.a(n249982),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[488]),
	.d(FE_OFN268_n249964));
   oa22s01 U263276 (.o(n249974),
	.a(n249982),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[487]),
	.d(FE_OFN268_n249964));
   oa22s01 U263277 (.o(n249976),
	.a(n249982),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[486]),
	.d(FE_OFN268_n249964));
   oa22s01 U263278 (.o(n249984),
	.a(n250018),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[479]),
	.d(n249999));
   oa22s01 U263279 (.o(n249985),
	.a(n250018),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[478]),
	.d(FE_OFN402_n249999));
   oa22s01 U263280 (.o(n249986),
	.a(n250018),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[477]),
	.d(FE_OFN402_n249999));
   oa22s01 U263281 (.o(n249988),
	.a(n250018),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[475]),
	.d(FE_OFN402_n249999));
   oa22s01 U263282 (.o(n249989),
	.a(n250018),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[474]),
	.d(FE_OFN402_n249999));
   oa22s01 U263283 (.o(n249990),
	.a(n250018),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[473]),
	.d(n249999));
   oa22s01 U263284 (.o(n249991),
	.a(n250018),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[472]),
	.d(n249999));
   oa22s01 U263285 (.o(n249992),
	.a(n250018),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[471]),
	.d(FE_OFN402_n249999));
   oa22s01 U263286 (.o(n249993),
	.a(n250018),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[470]),
	.d(FE_OFN402_n249999));
   oa22s01 U263287 (.o(n249994),
	.a(n250018),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[469]),
	.d(FE_OFN402_n249999));
   oa22s01 U263288 (.o(n249995),
	.a(n250018),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[468]),
	.d(FE_OFN402_n249999));
   oa22s01 U263289 (.o(n249996),
	.a(n250018),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[467]),
	.d(FE_OFN402_n249999));
   oa22s01 U263290 (.o(n249997),
	.a(n250018),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[466]),
	.d(FE_OFN402_n249999));
   oa22s01 U263291 (.o(n249998),
	.a(n250018),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[465]),
	.d(FE_OFN402_n249999));
   oa22s01 U263292 (.o(n250000),
	.a(n250018),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[464]),
	.d(FE_OFN402_n249999));
   oa22s01 U263293 (.o(n250001),
	.a(n250018),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[463]),
	.d(FE_OFN402_n249999));
   oa22s01 U263294 (.o(n250002),
	.a(n250018),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[462]),
	.d(FE_OFN402_n249999));
   oa22s01 U263295 (.o(n250004),
	.a(n250018),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[460]),
	.d(FE_OFN402_n249999));
   oa22s01 U263296 (.o(n250005),
	.a(n250018),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[459]),
	.d(FE_OFN402_n249999));
   oa22s01 U263297 (.o(n250006),
	.a(n250018),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[458]),
	.d(FE_OFN402_n249999));
   oa22s01 U263298 (.o(n250008),
	.a(n250018),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[456]),
	.d(FE_OFN402_n249999));
   oa22s01 U263299 (.o(n250009),
	.a(n250018),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[455]),
	.d(n249999));
   oa22s01 U263300 (.o(n250011),
	.a(n250018),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[454]),
	.d(FE_OFN402_n249999));
   oa22s01 U263301 (.o(n250020),
	.a(n250053),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[447]),
	.d(FE_OFN270_n250035));
   oa22s01 U263302 (.o(n250022),
	.a(n250053),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[445]),
	.d(FE_OFN270_n250035));
   oa22s01 U263303 (.o(n250023),
	.a(n250053),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[444]),
	.d(FE_OFN270_n250035));
   oa22s01 U263304 (.o(n250024),
	.a(n250053),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[443]),
	.d(FE_OFN270_n250035));
   oa22s01 U263305 (.o(n250025),
	.a(n250053),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[442]),
	.d(FE_OFN270_n250035));
   oa22s01 U263306 (.o(n250026),
	.a(n250053),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[441]),
	.d(FE_OFN270_n250035));
   oa22s01 U263307 (.o(n250027),
	.a(n250053),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[440]),
	.d(FE_OFN270_n250035));
   oa22s01 U263308 (.o(n250028),
	.a(n250053),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[439]),
	.d(FE_OFN270_n250035));
   oa22s01 U263309 (.o(n250029),
	.a(n250053),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[438]),
	.d(FE_OFN270_n250035));
   oa22s01 U263310 (.o(n250030),
	.a(n250053),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[437]),
	.d(FE_OFN270_n250035));
   oa22s01 U263311 (.o(n250031),
	.a(n250053),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[436]),
	.d(FE_OFN270_n250035));
   oa22s01 U263312 (.o(n250032),
	.a(n250053),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[435]),
	.d(FE_OFN270_n250035));
   oa22s01 U263313 (.o(n250033),
	.a(n250053),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[434]),
	.d(FE_OFN270_n250035));
   oa22s01 U263314 (.o(n250034),
	.a(n250053),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[433]),
	.d(FE_OFN270_n250035));
   oa22s01 U263315 (.o(n250036),
	.a(n250053),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[432]),
	.d(FE_OFN270_n250035));
   oa22s01 U263316 (.o(n250038),
	.a(n250053),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[430]),
	.d(FE_OFN270_n250035));
   oa22s01 U263317 (.o(n250039),
	.a(n250053),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[429]),
	.d(FE_OFN270_n250035));
   oa22s01 U263318 (.o(n250040),
	.a(n250053),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[428]),
	.d(FE_OFN270_n250035));
   oa22s01 U263319 (.o(n250042),
	.a(n250053),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[426]),
	.d(FE_OFN270_n250035));
   oa22s01 U263320 (.o(n250043),
	.a(n250053),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[425]),
	.d(FE_OFN270_n250035));
   oa22s01 U263321 (.o(n250044),
	.a(n250053),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[424]),
	.d(FE_OFN270_n250035));
   oa22s01 U263322 (.o(n250045),
	.a(n250053),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[423]),
	.d(FE_OFN270_n250035));
   oa22s01 U263323 (.o(n250047),
	.a(n250053),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[422]),
	.d(FE_OFN270_n250035));
   oa22s01 U263324 (.o(n250056),
	.a(n250089),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[415]),
	.d(FE_OFN404_n250071));
   oa22s01 U263325 (.o(n250057),
	.a(n250089),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[414]),
	.d(FE_OFN404_n250071));
   oa22s01 U263326 (.o(n250058),
	.a(n250089),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[413]),
	.d(n250071));
   oa22s01 U263327 (.o(n250059),
	.a(n250089),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[412]),
	.d(FE_OFN404_n250071));
   oa22s01 U263328 (.o(n250060),
	.a(n250089),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[411]),
	.d(FE_OFN404_n250071));
   oa22s01 U263329 (.o(n250061),
	.a(n250089),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[410]),
	.d(FE_OFN404_n250071));
   oa22s01 U263330 (.o(n250062),
	.a(n250089),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[409]),
	.d(FE_OFN404_n250071));
   oa22s01 U263331 (.o(n250063),
	.a(n250089),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[408]),
	.d(n250071));
   oa22s01 U263332 (.o(n250064),
	.a(n250089),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[407]),
	.d(n250071));
   oa22s01 U263333 (.o(n250065),
	.a(n250089),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[406]),
	.d(FE_OFN404_n250071));
   oa22s01 U263334 (.o(n250066),
	.a(n250089),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[405]),
	.d(FE_OFN404_n250071));
   oa22s01 U263335 (.o(n250067),
	.a(n250089),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[404]),
	.d(FE_OFN404_n250071));
   oa22s01 U263336 (.o(n250068),
	.a(n250089),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[403]),
	.d(FE_OFN404_n250071));
   oa22s01 U263337 (.o(n250069),
	.a(n250089),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[402]),
	.d(FE_OFN404_n250071));
   oa22s01 U263338 (.o(n250072),
	.a(n250089),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[400]),
	.d(FE_OFN404_n250071));
   oa22s01 U263339 (.o(n250073),
	.a(n250089),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[399]),
	.d(FE_OFN404_n250071));
   oa22s01 U263340 (.o(n250074),
	.a(n250089),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[398]),
	.d(FE_OFN404_n250071));
   oa22s01 U263341 (.o(n250076),
	.a(n250089),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[396]),
	.d(FE_OFN404_n250071));
   oa22s01 U263342 (.o(n250077),
	.a(n250089),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[395]),
	.d(FE_OFN404_n250071));
   oa22s01 U263343 (.o(n250078),
	.a(n250089),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[394]),
	.d(FE_OFN404_n250071));
   oa22s01 U263344 (.o(n250079),
	.a(n250089),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[393]),
	.d(FE_OFN404_n250071));
   oa22s01 U263345 (.o(n250080),
	.a(n250089),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[392]),
	.d(FE_OFN404_n250071));
   oa22s01 U263346 (.o(n250081),
	.a(n250089),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[391]),
	.d(FE_OFN404_n250071));
   oa22s01 U263347 (.o(n250083),
	.a(n250089),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[390]),
	.d(FE_OFN404_n250071));
   oa22s01 U263348 (.o(n250092),
	.a(n250126),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[383]),
	.d(FE_OFN192_n250107));
   oa22s01 U263349 (.o(n250094),
	.a(n250126),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[381]),
	.d(FE_OFN192_n250107));
   oa22s01 U263350 (.o(n250095),
	.a(n250126),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[380]),
	.d(FE_OFN192_n250107));
   oa22s01 U263351 (.o(n250096),
	.a(n250126),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[379]),
	.d(FE_OFN192_n250107));
   oa22s01 U263352 (.o(n250097),
	.a(n250126),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[378]),
	.d(FE_OFN193_n250107));
   oa22s01 U263353 (.o(n250098),
	.a(n250126),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[377]),
	.d(FE_OFN193_n250107));
   oa22s01 U263354 (.o(n250099),
	.a(n250126),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[376]),
	.d(FE_OFN192_n250107));
   oa22s01 U263355 (.o(n250100),
	.a(n250126),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[375]),
	.d(FE_OFN192_n250107));
   oa22s01 U263356 (.o(n250101),
	.a(n250126),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[374]),
	.d(FE_OFN193_n250107));
   oa22s01 U263357 (.o(n250102),
	.a(n250126),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[373]),
	.d(FE_OFN193_n250107));
   oa22s01 U263358 (.o(n250103),
	.a(n250126),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[372]),
	.d(FE_OFN193_n250107));
   oa22s01 U263359 (.o(n250105),
	.a(n250126),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[370]),
	.d(FE_OFN193_n250107));
   oa22s01 U263360 (.o(n250106),
	.a(n250126),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[369]),
	.d(FE_OFN193_n250107));
   oa22s01 U263361 (.o(n250108),
	.a(n250126),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[368]),
	.d(FE_OFN193_n250107));
   oa22s01 U263362 (.o(n250109),
	.a(n250126),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[367]),
	.d(FE_OFN192_n250107));
   oa22s01 U263363 (.o(n250110),
	.a(n250126),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[366]),
	.d(FE_OFN192_n250107));
   oa22s01 U263364 (.o(n250111),
	.a(n250126),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[365]),
	.d(FE_OFN192_n250107));
   oa22s01 U263365 (.o(n250112),
	.a(n250126),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[364]),
	.d(FE_OFN193_n250107));
   oa22s01 U263366 (.o(n250113),
	.a(n250126),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[363]),
	.d(FE_OFN193_n250107));
   oa22s01 U263367 (.o(n250114),
	.a(n250126),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[362]),
	.d(FE_OFN192_n250107));
   oa22s01 U263368 (.o(n250115),
	.a(n250126),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[361]),
	.d(FE_OFN192_n250107));
   oa22s01 U263369 (.o(n250116),
	.a(n250126),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[360]),
	.d(FE_OFN193_n250107));
   oa22s01 U263370 (.o(n250117),
	.a(n250126),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[359]),
	.d(FE_OFN192_n250107));
   oa22s01 U263371 (.o(n250119),
	.a(n250126),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[358]),
	.d(FE_OFN192_n250107));
   oa22s01 U263372 (.o(n250134),
	.a(n250162),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[346]),
	.d(FE_OFN272_n250144));
   oa22s01 U263373 (.o(n250136),
	.a(n250162),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[344]),
	.d(n250144));
   oa22s01 U263374 (.o(n250138),
	.a(FE_OFN406_n250162),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[342]),
	.d(FE_OFN272_n250144));
   oa22s01 U263375 (.o(n250140),
	.a(n250162),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[340]),
	.d(FE_OFN272_n250144));
   oa22s01 U263376 (.o(n250142),
	.a(n250162),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[338]),
	.d(FE_OFN272_n250144));
   oa22s01 U263377 (.o(n250146),
	.a(n250162),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[335]),
	.d(FE_OFN272_n250144));
   oa22s01 U263378 (.o(n250147),
	.a(n250162),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[334]),
	.d(FE_OFN272_n250144));
   oa22s01 U263379 (.o(n250153),
	.a(FE_OFN406_n250162),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[328]),
	.d(FE_OFN272_n250144));
   oa22s01 U263380 (.o(n250154),
	.a(FE_OFN406_n250162),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[327]),
	.d(FE_OFN272_n250144));
   oa22s01 U263381 (.o(n250165),
	.a(n250198),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[319]),
	.d(FE_OFN274_n250180));
   oa22s01 U263382 (.o(n250166),
	.a(n250198),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[318]),
	.d(FE_OFN274_n250180));
   oa22s01 U263383 (.o(n250167),
	.a(n250198),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[317]),
	.d(FE_OFN274_n250180));
   oa22s01 U263384 (.o(n250168),
	.a(n250198),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[316]),
	.d(FE_OFN274_n250180));
   oa22s01 U263385 (.o(n250169),
	.a(n250198),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[315]),
	.d(FE_OFN274_n250180));
   oa22s01 U263386 (.o(n250170),
	.a(n250198),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[314]),
	.d(FE_OFN274_n250180));
   oa22s01 U263387 (.o(n250171),
	.a(n250198),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[313]),
	.d(FE_OFN274_n250180));
   oa22s01 U263388 (.o(n250172),
	.a(n250198),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[312]),
	.d(FE_OFN274_n250180));
   oa22s01 U263389 (.o(n250174),
	.a(n250198),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[310]),
	.d(FE_OFN274_n250180));
   oa22s01 U263390 (.o(n250175),
	.a(n250198),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[309]),
	.d(FE_OFN274_n250180));
   oa22s01 U263391 (.o(n250176),
	.a(n250198),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[308]),
	.d(FE_OFN274_n250180));
   oa22s01 U263392 (.o(n250177),
	.a(n250198),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[307]),
	.d(FE_OFN274_n250180));
   oa22s01 U263393 (.o(n250178),
	.a(n250198),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[306]),
	.d(FE_OFN274_n250180));
   oa22s01 U263394 (.o(n250179),
	.a(n250198),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[305]),
	.d(FE_OFN274_n250180));
   oa22s01 U263395 (.o(n250181),
	.a(n250198),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[304]),
	.d(FE_OFN274_n250180));
   oa22s01 U263396 (.o(n250182),
	.a(n250198),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[303]),
	.d(FE_OFN274_n250180));
   oa22s01 U263397 (.o(n250183),
	.a(n250198),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[302]),
	.d(FE_OFN274_n250180));
   oa22s01 U263398 (.o(n250184),
	.a(n250198),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[301]),
	.d(FE_OFN274_n250180));
   oa22s01 U263399 (.o(n250185),
	.a(n250198),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[300]),
	.d(FE_OFN274_n250180));
   oa22s01 U263400 (.o(n250186),
	.a(n250198),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[299]),
	.d(FE_OFN274_n250180));
   oa22s01 U263401 (.o(n250187),
	.a(n250198),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[298]),
	.d(FE_OFN274_n250180));
   oa22s01 U263402 (.o(n250188),
	.a(n250198),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[297]),
	.d(FE_OFN274_n250180));
   oa22s01 U263403 (.o(n250190),
	.a(n250198),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[295]),
	.d(FE_OFN274_n250180));
   oa22s01 U263404 (.o(n250192),
	.a(n250198),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[294]),
	.d(FE_OFN274_n250180));
   oa22s01 U263405 (.o(n250239),
	.a(n250272),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[255]),
	.d(FE_OFN278_n250254));
   oa22s01 U263406 (.o(n250240),
	.a(n250272),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[254]),
	.d(FE_OFN278_n250254));
   oa22s01 U263407 (.o(n250241),
	.a(n250272),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[253]),
	.d(FE_OFN278_n250254));
   oa22s01 U263408 (.o(n250242),
	.a(n250272),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[252]),
	.d(FE_OFN278_n250254));
   oa22s01 U263409 (.o(n250244),
	.a(n250272),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[250]),
	.d(FE_OFN278_n250254));
   oa22s01 U263410 (.o(n250245),
	.a(n250272),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[249]),
	.d(FE_OFN278_n250254));
   oa22s01 U263411 (.o(n250246),
	.a(n250272),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[248]),
	.d(FE_OFN278_n250254));
   oa22s01 U263412 (.o(n250247),
	.a(n250272),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[247]),
	.d(FE_OFN278_n250254));
   oa22s01 U263413 (.o(n250248),
	.a(n250272),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[246]),
	.d(FE_OFN278_n250254));
   oa22s01 U263414 (.o(n250249),
	.a(n250272),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[245]),
	.d(FE_OFN278_n250254));
   oa22s01 U263415 (.o(n250250),
	.a(n250272),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[244]),
	.d(FE_OFN278_n250254));
   oa22s01 U263416 (.o(n250251),
	.a(n250272),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[243]),
	.d(FE_OFN278_n250254));
   oa22s01 U263417 (.o(n250252),
	.a(n250272),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[242]),
	.d(FE_OFN278_n250254));
   oa22s01 U263418 (.o(n250253),
	.a(n250272),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[241]),
	.d(FE_OFN278_n250254));
   oa22s01 U263419 (.o(n250255),
	.a(n250272),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[240]),
	.d(FE_OFN278_n250254));
   oa22s01 U263420 (.o(n250256),
	.a(n250272),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[239]),
	.d(FE_OFN278_n250254));
   oa22s01 U263421 (.o(n250257),
	.a(n250272),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[238]),
	.d(FE_OFN278_n250254));
   oa22s01 U263422 (.o(n250258),
	.a(n250272),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[237]),
	.d(FE_OFN278_n250254));
   oa22s01 U263423 (.o(n250260),
	.a(n250272),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[235]),
	.d(FE_OFN278_n250254));
   oa22s01 U263424 (.o(n250261),
	.a(n250272),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[234]),
	.d(FE_OFN278_n250254));
   oa22s01 U263425 (.o(n250262),
	.a(n250272),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[233]),
	.d(FE_OFN278_n250254));
   oa22s01 U263426 (.o(n250263),
	.a(n250272),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[232]),
	.d(FE_OFN278_n250254));
   oa22s01 U263427 (.o(n250264),
	.a(n250272),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[231]),
	.d(FE_OFN278_n250254));
   oa22s01 U263428 (.o(n250266),
	.a(n250272),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[230]),
	.d(FE_OFN278_n250254));
   oa22s01 U263429 (.o(n250274),
	.a(n250307),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[223]),
	.d(FE_OFN408_n250289));
   oa22s01 U263430 (.o(n250275),
	.a(n250307),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[222]),
	.d(FE_OFN408_n250289));
   oa22s01 U263431 (.o(n250277),
	.a(n250307),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[220]),
	.d(FE_OFN408_n250289));
   oa22s01 U263432 (.o(n250278),
	.a(n250307),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[219]),
	.d(FE_OFN408_n250289));
   oa22s01 U263433 (.o(n250279),
	.a(n250307),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[218]),
	.d(FE_OFN408_n250289));
   oa22s01 U263434 (.o(n250280),
	.a(n250307),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[217]),
	.d(FE_OFN408_n250289));
   oa22s01 U263435 (.o(n250281),
	.a(n250307),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[216]),
	.d(FE_OFN408_n250289));
   oa22s01 U263436 (.o(n250282),
	.a(n250307),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[215]),
	.d(FE_OFN408_n250289));
   oa22s01 U263437 (.o(n250283),
	.a(n250307),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[214]),
	.d(FE_OFN408_n250289));
   oa22s01 U263438 (.o(n250284),
	.a(n250307),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[213]),
	.d(FE_OFN408_n250289));
   oa22s01 U263439 (.o(n250285),
	.a(n250307),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[212]),
	.d(FE_OFN408_n250289));
   oa22s01 U263440 (.o(n250286),
	.a(n250307),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[211]),
	.d(FE_OFN408_n250289));
   oa22s01 U263441 (.o(n250287),
	.a(n250307),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[210]),
	.d(FE_OFN408_n250289));
   oa22s01 U263442 (.o(n250288),
	.a(n250307),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[209]),
	.d(FE_OFN408_n250289));
   oa22s01 U263443 (.o(n250290),
	.a(n250307),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[208]),
	.d(FE_OFN408_n250289));
   oa22s01 U263444 (.o(n250291),
	.a(n250307),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[207]),
	.d(FE_OFN408_n250289));
   oa22s01 U263445 (.o(n250293),
	.a(n250307),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[205]),
	.d(FE_OFN408_n250289));
   oa22s01 U263446 (.o(n250294),
	.a(n250307),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[204]),
	.d(FE_OFN408_n250289));
   oa22s01 U263447 (.o(n250295),
	.a(n250307),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[203]),
	.d(FE_OFN408_n250289));
   oa22s01 U263448 (.o(n250297),
	.a(n250307),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[201]),
	.d(FE_OFN408_n250289));
   oa22s01 U263449 (.o(n250298),
	.a(n250307),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[200]),
	.d(FE_OFN408_n250289));
   oa22s01 U263450 (.o(n250299),
	.a(n250307),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[199]),
	.d(FE_OFN408_n250289));
   oa22s01 U263451 (.o(n250301),
	.a(n250307),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[198]),
	.d(FE_OFN408_n250289));
   oa22s01 U263452 (.o(n250310),
	.a(n250343),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[190]),
	.d(FE_OFN280_n250324));
   oa22s01 U263453 (.o(n250311),
	.a(n250343),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[189]),
	.d(FE_OFN280_n250324));
   oa22s01 U263454 (.o(n250312),
	.a(n250343),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[188]),
	.d(FE_OFN280_n250324));
   oa22s01 U263455 (.o(n250313),
	.a(n250343),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[187]),
	.d(FE_OFN280_n250324));
   oa22s01 U263456 (.o(n250314),
	.a(n250343),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[186]),
	.d(FE_OFN280_n250324));
   oa22s01 U263457 (.o(n250315),
	.a(n250343),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[185]),
	.d(FE_OFN280_n250324));
   oa22s01 U263458 (.o(n250316),
	.a(n250343),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[184]),
	.d(FE_OFN280_n250324));
   oa22s01 U263459 (.o(n250317),
	.a(n250343),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[183]),
	.d(FE_OFN280_n250324));
   oa22s01 U263460 (.o(n250318),
	.a(n250343),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[182]),
	.d(FE_OFN280_n250324));
   oa22s01 U263461 (.o(n250319),
	.a(n250343),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[181]),
	.d(FE_OFN280_n250324));
   oa22s01 U263462 (.o(n250320),
	.a(n250343),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[180]),
	.d(FE_OFN280_n250324));
   oa22s01 U263463 (.o(n250321),
	.a(n250343),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[179]),
	.d(FE_OFN280_n250324));
   oa22s01 U263464 (.o(n250322),
	.a(n250343),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[178]),
	.d(FE_OFN280_n250324));
   oa22s01 U263465 (.o(n250323),
	.a(n250343),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[177]),
	.d(FE_OFN280_n250324));
   oa22s01 U263466 (.o(n250326),
	.a(n250343),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[175]),
	.d(FE_OFN280_n250324));
   oa22s01 U263467 (.o(n250327),
	.a(n250343),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[174]),
	.d(FE_OFN280_n250324));
   oa22s01 U263468 (.o(n250328),
	.a(n250343),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[173]),
	.d(FE_OFN280_n250324));
   oa22s01 U263469 (.o(n250330),
	.a(n250343),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[171]),
	.d(FE_OFN280_n250324));
   oa22s01 U263470 (.o(n250331),
	.a(n250343),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[170]),
	.d(FE_OFN280_n250324));
   oa22s01 U263471 (.o(n250332),
	.a(n250343),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[169]),
	.d(FE_OFN280_n250324));
   oa22s01 U263472 (.o(n250333),
	.a(n250343),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[168]),
	.d(FE_OFN280_n250324));
   oa22s01 U263473 (.o(n250334),
	.a(n250343),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[167]),
	.d(FE_OFN280_n250324));
   oa22s01 U263474 (.o(n250336),
	.a(n250343),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[166]),
	.d(FE_OFN280_n250324));
   oa22s01 U263475 (.o(n250345),
	.a(n250378),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[159]),
	.d(FE_OFN410_n250360));
   oa22s01 U263476 (.o(n250346),
	.a(n250378),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[158]),
	.d(FE_OFN410_n250360));
   oa22s01 U263477 (.o(n250348),
	.a(n250378),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[156]),
	.d(FE_OFN410_n250360));
   oa22s01 U263478 (.o(n250349),
	.a(n250378),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[155]),
	.d(FE_OFN410_n250360));
   oa22s01 U263479 (.o(n250350),
	.a(n250378),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[154]),
	.d(FE_OFN410_n250360));
   oa22s01 U263480 (.o(n250351),
	.a(n250378),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[153]),
	.d(FE_OFN410_n250360));
   oa22s01 U263481 (.o(n250352),
	.a(n250378),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[152]),
	.d(FE_OFN410_n250360));
   oa22s01 U263482 (.o(n250353),
	.a(n250378),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[151]),
	.d(FE_OFN410_n250360));
   oa22s01 U263483 (.o(n250354),
	.a(n250378),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[150]),
	.d(FE_OFN410_n250360));
   oa22s01 U263484 (.o(n250355),
	.a(n250378),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[149]),
	.d(FE_OFN410_n250360));
   oa22s01 U263485 (.o(n250356),
	.a(n250378),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[148]),
	.d(FE_OFN410_n250360));
   oa22s01 U263486 (.o(n250357),
	.a(n250378),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[147]),
	.d(FE_OFN410_n250360));
   oa22s01 U263487 (.o(n250359),
	.a(n250378),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[145]),
	.d(FE_OFN410_n250360));
   oa22s01 U263488 (.o(n250361),
	.a(n250378),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[144]),
	.d(FE_OFN410_n250360));
   oa22s01 U263489 (.o(n250362),
	.a(n250378),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[143]),
	.d(FE_OFN410_n250360));
   oa22s01 U263490 (.o(n250363),
	.a(n250378),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[142]),
	.d(FE_OFN410_n250360));
   oa22s01 U263491 (.o(n250364),
	.a(n250378),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[141]),
	.d(FE_OFN410_n250360));
   oa22s01 U263492 (.o(n250365),
	.a(n250378),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[140]),
	.d(FE_OFN410_n250360));
   oa22s01 U263493 (.o(n250366),
	.a(n250378),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[139]),
	.d(FE_OFN410_n250360));
   oa22s01 U263494 (.o(n250367),
	.a(n250378),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[138]),
	.d(FE_OFN410_n250360));
   oa22s01 U263495 (.o(n250368),
	.a(n250378),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[137]),
	.d(FE_OFN410_n250360));
   oa22s01 U263496 (.o(n250369),
	.a(n250378),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[136]),
	.d(FE_OFN410_n250360));
   oa22s01 U263497 (.o(n250370),
	.a(n250378),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[135]),
	.d(FE_OFN410_n250360));
   oa22s01 U263498 (.o(n250372),
	.a(n250378),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[134]),
	.d(FE_OFN410_n250360));
   oa22s01 U263499 (.o(n250381),
	.a(n250413),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[126]),
	.d(FE_OFN195_n250395));
   oa22s01 U263500 (.o(n250382),
	.a(n250413),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[125]),
	.d(FE_OFN195_n250395));
   oa22s01 U263501 (.o(n250383),
	.a(n250413),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[124]),
	.d(FE_OFN195_n250395));
   oa22s01 U263502 (.o(n250384),
	.a(n250413),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[123]),
	.d(FE_OFN195_n250395));
   oa22s01 U263503 (.o(n250385),
	.a(n250413),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[122]),
	.d(FE_OFN195_n250395));
   oa22s01 U263504 (.o(n250386),
	.a(n250413),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[121]),
	.d(FE_OFN195_n250395));
   oa22s01 U263505 (.o(n250387),
	.a(n250413),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[120]),
	.d(FE_OFN195_n250395));
   oa22s01 U263506 (.o(n250388),
	.a(n250413),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[119]),
	.d(FE_OFN195_n250395));
   oa22s01 U263507 (.o(n250389),
	.a(n250413),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[118]),
	.d(FE_OFN195_n250395));
   oa22s01 U263508 (.o(n250390),
	.a(n250413),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[117]),
	.d(FE_OFN195_n250395));
   oa22s01 U263509 (.o(n250392),
	.a(n250413),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[115]),
	.d(FE_OFN195_n250395));
   oa22s01 U263510 (.o(n250393),
	.a(n250413),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[114]),
	.d(FE_OFN195_n250395));
   oa22s01 U263511 (.o(n250394),
	.a(n250413),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[113]),
	.d(FE_OFN195_n250395));
   oa22s01 U263512 (.o(n250396),
	.a(n250413),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[112]),
	.d(FE_OFN195_n250395));
   oa22s01 U263513 (.o(n250397),
	.a(n250413),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[111]),
	.d(FE_OFN195_n250395));
   oa22s01 U263514 (.o(n250398),
	.a(n250413),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[110]),
	.d(FE_OFN195_n250395));
   oa22s01 U263515 (.o(n250399),
	.a(n250413),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[109]),
	.d(FE_OFN195_n250395));
   oa22s01 U263516 (.o(n250400),
	.a(n250413),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[108]),
	.d(FE_OFN195_n250395));
   oa22s01 U263517 (.o(n250401),
	.a(n250413),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[107]),
	.d(FE_OFN195_n250395));
   oa22s01 U263518 (.o(n250402),
	.a(n250413),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[106]),
	.d(FE_OFN195_n250395));
   oa22s01 U263519 (.o(n250403),
	.a(n250413),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[105]),
	.d(FE_OFN195_n250395));
   oa22s01 U263520 (.o(n250404),
	.a(n250413),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[104]),
	.d(FE_OFN195_n250395));
   oa22s01 U263521 (.o(n250405),
	.a(n250413),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[103]),
	.d(FE_OFN195_n250395));
   oa22s01 U263522 (.o(n250407),
	.a(n250413),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[102]),
	.d(FE_OFN195_n250395));
   oa22s01 U263523 (.o(n250451),
	.a(n250484),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[63]),
	.d(FE_OFN284_n250466));
   oa22s01 U263524 (.o(n250452),
	.a(n250484),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[62]),
	.d(FE_OFN284_n250466));
   oa22s01 U263525 (.o(n250453),
	.a(n250484),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[61]),
	.d(FE_OFN284_n250466));
   oa22s01 U263526 (.o(n250454),
	.a(n250484),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[60]),
	.d(FE_OFN284_n250466));
   oa22s01 U263527 (.o(n250455),
	.a(n250484),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[59]),
	.d(FE_OFN284_n250466));
   oa22s01 U263528 (.o(n250456),
	.a(n250484),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[58]),
	.d(FE_OFN284_n250466));
   oa22s01 U263529 (.o(n250457),
	.a(n250484),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[57]),
	.d(FE_OFN284_n250466));
   oa22s01 U263530 (.o(n250459),
	.a(n250484),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[55]),
	.d(FE_OFN284_n250466));
   oa22s01 U263531 (.o(n250460),
	.a(n250484),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[54]),
	.d(FE_OFN284_n250466));
   oa22s01 U263532 (.o(n250461),
	.a(n250484),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[53]),
	.d(FE_OFN284_n250466));
   oa22s01 U263533 (.o(n250462),
	.a(n250484),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[52]),
	.d(FE_OFN284_n250466));
   oa22s01 U263534 (.o(n250463),
	.a(n250484),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[51]),
	.d(FE_OFN284_n250466));
   oa22s01 U263535 (.o(n250464),
	.a(n250484),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[50]),
	.d(FE_OFN284_n250466));
   oa22s01 U263536 (.o(n250465),
	.a(n250484),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[49]),
	.d(FE_OFN284_n250466));
   oa22s01 U263537 (.o(n250467),
	.a(n250484),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[48]),
	.d(FE_OFN284_n250466));
   oa22s01 U263538 (.o(n250468),
	.a(n250484),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[47]),
	.d(n250466));
   oa22s01 U263539 (.o(n250469),
	.a(n250484),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[46]),
	.d(FE_OFN284_n250466));
   oa22s01 U263540 (.o(n250470),
	.a(n250484),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[45]),
	.d(n250466));
   oa22s01 U263541 (.o(n250471),
	.a(n250484),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[44]),
	.d(FE_OFN284_n250466));
   oa22s01 U263542 (.o(n250472),
	.a(n250484),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[43]),
	.d(FE_OFN284_n250466));
   oa22s01 U263543 (.o(n250473),
	.a(n250484),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[42]),
	.d(n250466));
   oa22s01 U263544 (.o(n250475),
	.a(n250484),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[40]),
	.d(FE_OFN284_n250466));
   oa22s01 U263545 (.o(n250476),
	.a(n250484),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[39]),
	.d(n250466));
   oa22s01 U263546 (.o(n250478),
	.a(n250484),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[38]),
	.d(FE_OFN284_n250466));
   oa22s01 U263547 (.o(n250487),
	.a(n250520),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[31]),
	.d(n250502));
   oa22s01 U263548 (.o(n250488),
	.a(n250520),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[30]),
	.d(FE_OFN286_n250502));
   oa22s01 U263549 (.o(n250489),
	.a(n250520),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[29]),
	.d(n250502));
   oa22s01 U263550 (.o(n250490),
	.a(n250520),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[28]),
	.d(n250502));
   oa22s01 U263551 (.o(n250491),
	.a(n250520),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[27]),
	.d(n250502));
   oa22s01 U263552 (.o(n250493),
	.a(n250520),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[25]),
	.d(FE_OFN286_n250502));
   oa22s01 U263553 (.o(n250494),
	.a(n250520),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[24]),
	.d(n250502));
   oa22s01 U263554 (.o(n250495),
	.a(n250520),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[23]),
	.d(n250502));
   oa22s01 U263555 (.o(n250496),
	.a(n250520),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[22]),
	.d(FE_OFN286_n250502));
   oa22s01 U263556 (.o(n250497),
	.a(n250520),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[21]),
	.d(FE_OFN286_n250502));
   oa22s01 U263557 (.o(n250498),
	.a(n250520),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[20]),
	.d(FE_OFN286_n250502));
   oa22s01 U263558 (.o(n250499),
	.a(n250520),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[19]),
	.d(FE_OFN286_n250502));
   oa22s01 U263559 (.o(n250500),
	.a(n250520),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[18]),
	.d(FE_OFN286_n250502));
   oa22s01 U263560 (.o(n250501),
	.a(n250520),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[17]),
	.d(FE_OFN286_n250502));
   oa22s01 U263561 (.o(n250503),
	.a(n250520),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[16]),
	.d(FE_OFN286_n250502));
   oa22s01 U263562 (.o(n250504),
	.a(n250520),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[15]),
	.d(n250502));
   oa22s01 U263563 (.o(n250505),
	.a(n250520),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[14]),
	.d(n250502));
   oa22s01 U263564 (.o(n250506),
	.a(n250520),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[13]),
	.d(n250502));
   oa22s01 U263565 (.o(n250507),
	.a(n250520),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[12]),
	.d(FE_OFN286_n250502));
   oa22s01 U263566 (.o(n250509),
	.a(n250520),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[10]),
	.d(n250502));
   oa22s01 U263567 (.o(n250510),
	.a(n250520),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[9]),
	.d(n250502));
   oa22s01 U263568 (.o(n250511),
	.a(n250520),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[8]),
	.d(FE_OFN286_n250502));
   oa22s01 U263569 (.o(n250512),
	.a(n250520),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[7]),
	.d(n250502));
   oa22s01 U263570 (.o(n250514),
	.a(n250520),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[6]),
	.d(n250502));
   oa22s01 U263571 (.o(n250522),
	.a(n250556),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1023]),
	.d(FE_OFN288_n250540));
   oa22s01 U263572 (.o(n250523),
	.a(n250556),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1022]),
	.d(FE_OFN288_n250540));
   oa22s01 U263573 (.o(n250524),
	.a(n250556),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1021]),
	.d(FE_OFN288_n250540));
   oa22s01 U263574 (.o(n250526),
	.a(n250556),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1019]),
	.d(FE_OFN288_n250540));
   oa22s01 U263575 (.o(n250527),
	.a(n250556),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1018]),
	.d(FE_OFN288_n250540));
   oa22s01 U263576 (.o(n250528),
	.a(n250556),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1017]),
	.d(FE_OFN288_n250540));
   oa22s01 U263577 (.o(n250529),
	.a(n250556),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1016]),
	.d(FE_OFN288_n250540));
   oa22s01 U263578 (.o(n250530),
	.a(n250556),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1015]),
	.d(FE_OFN288_n250540));
   oa22s01 U263579 (.o(n250531),
	.a(n250556),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1014]),
	.d(FE_OFN288_n250540));
   oa22s01 U263580 (.o(n250532),
	.a(n250556),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1013]),
	.d(FE_OFN288_n250540));
   oa22s01 U263581 (.o(n250533),
	.a(n250556),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1012]),
	.d(FE_OFN288_n250540));
   oa22s01 U263582 (.o(n250534),
	.a(n250556),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1011]),
	.d(FE_OFN288_n250540));
   oa22s01 U263583 (.o(n250535),
	.a(n250556),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1010]),
	.d(FE_OFN288_n250540));
   oa22s01 U263584 (.o(n250536),
	.a(n250556),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1009]),
	.d(FE_OFN288_n250540));
   oa22s01 U263585 (.o(n250537),
	.a(n250556),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1008]),
	.d(FE_OFN288_n250540));
   oa22s01 U263586 (.o(n250538),
	.a(n250556),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1007]),
	.d(FE_OFN288_n250540));
   oa22s01 U263587 (.o(n250539),
	.a(n250556),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1006]),
	.d(FE_OFN288_n250540));
   oa22s01 U263588 (.o(n250542),
	.a(n250556),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1004]),
	.d(FE_OFN288_n250540));
   oa22s01 U263589 (.o(n250543),
	.a(n250556),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1003]),
	.d(FE_OFN288_n250540));
   oa22s01 U263590 (.o(n250544),
	.a(n250556),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1002]),
	.d(FE_OFN288_n250540));
   oa22s01 U263591 (.o(n250546),
	.a(n250556),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1000]),
	.d(FE_OFN288_n250540));
   oa22s01 U263592 (.o(n250547),
	.a(n250556),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[999]),
	.d(FE_OFN288_n250540));
   oa22s01 U263593 (.o(n250549),
	.a(n250556),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[998]),
	.d(FE_OFN288_n250540));
   oa22s01 U263594 (.o(n250558),
	.a(n250591),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[991]),
	.d(FE_OFN412_n250576));
   oa22s01 U263595 (.o(n250560),
	.a(n250591),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[989]),
	.d(FE_OFN412_n250576));
   oa22s01 U263596 (.o(n250561),
	.a(n250591),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[988]),
	.d(FE_OFN412_n250576));
   oa22s01 U263597 (.o(n250562),
	.a(n250591),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[987]),
	.d(FE_OFN412_n250576));
   oa22s01 U263598 (.o(n250563),
	.a(n250591),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[986]),
	.d(FE_OFN412_n250576));
   oa22s01 U263599 (.o(n250564),
	.a(n250591),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[985]),
	.d(FE_OFN412_n250576));
   oa22s01 U263600 (.o(n250565),
	.a(n250591),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[984]),
	.d(FE_OFN412_n250576));
   oa22s01 U263601 (.o(n250566),
	.a(n250591),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[983]),
	.d(FE_OFN412_n250576));
   oa22s01 U263602 (.o(n250567),
	.a(n250591),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[982]),
	.d(FE_OFN412_n250576));
   oa22s01 U263603 (.o(n250568),
	.a(n250591),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[981]),
	.d(FE_OFN412_n250576));
   oa22s01 U263604 (.o(n250569),
	.a(n250591),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[980]),
	.d(FE_OFN412_n250576));
   oa22s01 U263605 (.o(n250570),
	.a(n250591),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[979]),
	.d(FE_OFN412_n250576));
   oa22s01 U263606 (.o(n250571),
	.a(n250591),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[978]),
	.d(FE_OFN412_n250576));
   oa22s01 U263607 (.o(n250572),
	.a(n250591),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[977]),
	.d(FE_OFN412_n250576));
   oa22s01 U263608 (.o(n250573),
	.a(n250591),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[976]),
	.d(FE_OFN412_n250576));
   oa22s01 U263609 (.o(n250575),
	.a(n250591),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[974]),
	.d(FE_OFN412_n250576));
   oa22s01 U263610 (.o(n250577),
	.a(n250591),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[973]),
	.d(FE_OFN412_n250576));
   oa22s01 U263611 (.o(n250578),
	.a(n250591),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[972]),
	.d(FE_OFN412_n250576));
   oa22s01 U263612 (.o(n250580),
	.a(n250591),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[970]),
	.d(FE_OFN412_n250576));
   oa22s01 U263613 (.o(n250581),
	.a(n250591),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[969]),
	.d(FE_OFN412_n250576));
   oa22s01 U263614 (.o(n250582),
	.a(n250591),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[968]),
	.d(FE_OFN412_n250576));
   oa22s01 U263615 (.o(n250583),
	.a(n250591),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[967]),
	.d(FE_OFN412_n250576));
   oa22s01 U263616 (.o(n250585),
	.a(n250591),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[966]),
	.d(FE_OFN412_n250576));
   oa22s01 U263617 (.o(n250593),
	.a(n250626),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[959]),
	.d(FE_OFN290_n250611));
   oa22s01 U263618 (.o(n250594),
	.a(n250626),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[958]),
	.d(FE_OFN290_n250611));
   oa22s01 U263619 (.o(n250595),
	.a(n250626),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[957]),
	.d(FE_OFN290_n250611));
   oa22s01 U263620 (.o(n250597),
	.a(n250626),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[955]),
	.d(FE_OFN290_n250611));
   oa22s01 U263621 (.o(n250598),
	.a(n250626),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[954]),
	.d(FE_OFN290_n250611));
   oa22s01 U263622 (.o(n250599),
	.a(n250626),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[953]),
	.d(FE_OFN290_n250611));
   oa22s01 U263623 (.o(n250600),
	.a(n250626),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[952]),
	.d(FE_OFN290_n250611));
   oa22s01 U263624 (.o(n250601),
	.a(n250626),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[951]),
	.d(FE_OFN290_n250611));
   oa22s01 U263625 (.o(n250602),
	.a(n250626),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[950]),
	.d(FE_OFN290_n250611));
   oa22s01 U263626 (.o(n250603),
	.a(n250626),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[949]),
	.d(FE_OFN290_n250611));
   oa22s01 U263627 (.o(n250604),
	.a(n250626),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[948]),
	.d(FE_OFN290_n250611));
   oa22s01 U263628 (.o(n250605),
	.a(n250626),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[947]),
	.d(FE_OFN290_n250611));
   oa22s01 U263629 (.o(n250606),
	.a(n250626),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[946]),
	.d(FE_OFN290_n250611));
   oa22s01 U263630 (.o(n250608),
	.a(n250626),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[944]),
	.d(FE_OFN290_n250611));
   oa22s01 U263631 (.o(n250609),
	.a(n250626),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[943]),
	.d(FE_OFN290_n250611));
   oa22s01 U263632 (.o(n250610),
	.a(n250626),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[942]),
	.d(FE_OFN290_n250611));
   oa22s01 U263633 (.o(n250612),
	.a(n250626),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[941]),
	.d(FE_OFN290_n250611));
   oa22s01 U263634 (.o(n250613),
	.a(n250626),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[940]),
	.d(FE_OFN290_n250611));
   oa22s01 U263635 (.o(n250614),
	.a(n250626),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[939]),
	.d(FE_OFN290_n250611));
   oa22s01 U263636 (.o(n250615),
	.a(n250626),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[938]),
	.d(FE_OFN290_n250611));
   oa22s01 U263637 (.o(n250616),
	.a(n250626),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[937]),
	.d(FE_OFN290_n250611));
   oa22s01 U263638 (.o(n250617),
	.a(n250626),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[936]),
	.d(FE_OFN290_n250611));
   oa22s01 U263639 (.o(n250618),
	.a(n250626),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[935]),
	.d(FE_OFN290_n250611));
   oa22s01 U263640 (.o(n250620),
	.a(n250626),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[934]),
	.d(FE_OFN290_n250611));
   oa22s01 U263641 (.o(n250628),
	.a(n250662),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[927]),
	.d(FE_OFN414_n250646));
   oa22s01 U263642 (.o(n250630),
	.a(n250662),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[925]),
	.d(FE_OFN414_n250646));
   oa22s01 U263643 (.o(n250631),
	.a(n250662),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[924]),
	.d(FE_OFN414_n250646));
   oa22s01 U263644 (.o(n250632),
	.a(n250662),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[923]),
	.d(FE_OFN414_n250646));
   oa22s01 U263645 (.o(n250633),
	.a(n250662),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[922]),
	.d(FE_OFN414_n250646));
   oa22s01 U263646 (.o(n250634),
	.a(n250662),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[921]),
	.d(FE_OFN414_n250646));
   oa22s01 U263647 (.o(n250635),
	.a(n250662),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[920]),
	.d(FE_OFN414_n250646));
   oa22s01 U263648 (.o(n250636),
	.a(n250662),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[919]),
	.d(FE_OFN414_n250646));
   oa22s01 U263649 (.o(n250637),
	.a(n250662),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[918]),
	.d(FE_OFN414_n250646));
   oa22s01 U263650 (.o(n250638),
	.a(n250662),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[917]),
	.d(FE_OFN414_n250646));
   oa22s01 U263651 (.o(n250639),
	.a(n250662),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[916]),
	.d(FE_OFN414_n250646));
   oa22s01 U263652 (.o(n250641),
	.a(n250662),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[914]),
	.d(FE_OFN414_n250646));
   oa22s01 U263653 (.o(n250642),
	.a(n250662),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[913]),
	.d(FE_OFN414_n250646));
   oa22s01 U263654 (.o(n250643),
	.a(n250662),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[912]),
	.d(FE_OFN414_n250646));
   oa22s01 U263655 (.o(n250644),
	.a(n250662),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[911]),
	.d(FE_OFN414_n250646));
   oa22s01 U263656 (.o(n250645),
	.a(n250662),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[910]),
	.d(FE_OFN414_n250646));
   oa22s01 U263657 (.o(n250647),
	.a(n250662),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[909]),
	.d(FE_OFN414_n250646));
   oa22s01 U263658 (.o(n250648),
	.a(n250662),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[908]),
	.d(FE_OFN414_n250646));
   oa22s01 U263659 (.o(n250649),
	.a(n250662),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[907]),
	.d(FE_OFN414_n250646));
   oa22s01 U263660 (.o(n250650),
	.a(n250662),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[906]),
	.d(FE_OFN414_n250646));
   oa22s01 U263661 (.o(n250651),
	.a(n250662),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[905]),
	.d(FE_OFN414_n250646));
   oa22s01 U263662 (.o(n250652),
	.a(n250662),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[904]),
	.d(FE_OFN414_n250646));
   oa22s01 U263663 (.o(n250653),
	.a(n250662),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[903]),
	.d(FE_OFN414_n250646));
   oa22s01 U263664 (.o(n250655),
	.a(n250662),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[902]),
	.d(FE_OFN414_n250646));
   oa22s01 U263665 (.o(n250664),
	.a(n250697),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[895]),
	.d(n250682));
   oa22s01 U263666 (.o(n250665),
	.a(n250697),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[894]),
	.d(FE_OFN198_n250682));
   oa22s01 U263667 (.o(n250666),
	.a(n250697),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[893]),
	.d(FE_OFN197_n250682));
   oa22s01 U263668 (.o(n250667),
	.a(n250697),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[892]),
	.d(n250682));
   oa22s01 U263669 (.o(n250668),
	.a(n250697),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[891]),
	.d(FE_OFN197_n250682));
   oa22s01 U263670 (.o(n250669),
	.a(n250697),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[890]),
	.d(FE_OFN198_n250682));
   oa22s01 U263671 (.o(n250670),
	.a(n250697),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[889]),
	.d(FE_OFN198_n250682));
   oa22s01 U263672 (.o(n250671),
	.a(n250697),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[888]),
	.d(FE_OFN197_n250682));
   oa22s01 U263673 (.o(n250672),
	.a(n250697),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[887]),
	.d(n250682));
   oa22s01 U263674 (.o(n250673),
	.a(n250697),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[886]),
	.d(FE_OFN198_n250682));
   oa22s01 U263675 (.o(n250675),
	.a(n250697),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[884]),
	.d(FE_OFN198_n250682));
   oa22s01 U263676 (.o(n250676),
	.a(n250697),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[883]),
	.d(FE_OFN198_n250682));
   oa22s01 U263677 (.o(n250677),
	.a(n250697),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[882]),
	.d(FE_OFN198_n250682));
   oa22s01 U263678 (.o(n250678),
	.a(n250697),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[881]),
	.d(FE_OFN198_n250682));
   oa22s01 U263679 (.o(n250679),
	.a(n250697),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[880]),
	.d(FE_OFN198_n250682));
   oa22s01 U263680 (.o(n250680),
	.a(n250697),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[879]),
	.d(FE_OFN197_n250682));
   oa22s01 U263681 (.o(n250681),
	.a(n250697),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[878]),
	.d(n250682));
   oa22s01 U263682 (.o(n250683),
	.a(n250697),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[877]),
	.d(n250682));
   oa22s01 U263683 (.o(n250684),
	.a(n250697),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[876]),
	.d(FE_OFN198_n250682));
   oa22s01 U263684 (.o(n250685),
	.a(n250697),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[875]),
	.d(FE_OFN198_n250682));
   oa22s01 U263685 (.o(n250686),
	.a(n250697),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[874]),
	.d(FE_OFN198_n250682));
   oa22s01 U263686 (.o(n250687),
	.a(n250697),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[873]),
	.d(FE_OFN197_n250682));
   oa22s01 U263687 (.o(n250688),
	.a(n250697),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[872]),
	.d(FE_OFN198_n250682));
   oa22s01 U263688 (.o(n250689),
	.a(n250697),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[871]),
	.d(FE_OFN198_n250682));
   oa22s01 U263689 (.o(n250699),
	.a(n250732),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[863]),
	.d(FE_OFN563_n250717));
   oa22s01 U263690 (.o(n250700),
	.a(n250732),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[862]),
	.d(FE_OFN563_n250717));
   oa22s01 U263691 (.o(n250701),
	.a(n250732),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[861]),
	.d(FE_OFN292_n250717));
   oa22s01 U263692 (.o(n250702),
	.a(n250732),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[860]),
	.d(FE_OFN292_n250717));
   oa22s01 U263693 (.o(n250703),
	.a(n250732),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[859]),
	.d(FE_OFN292_n250717));
   oa22s01 U263694 (.o(n250704),
	.a(n250732),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[858]),
	.d(FE_OFN292_n250717));
   oa22s01 U263695 (.o(n250706),
	.a(n250732),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[856]),
	.d(FE_OFN292_n250717));
   oa22s01 U263696 (.o(n250708),
	.a(n250732),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[854]),
	.d(FE_OFN563_n250717));
   oa22s01 U263697 (.o(n250710),
	.a(n250732),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[852]),
	.d(FE_OFN292_n250717));
   oa22s01 U263698 (.o(n250712),
	.a(n250732),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[850]),
	.d(FE_OFN563_n250717));
   oa22s01 U263699 (.o(n250715),
	.a(n250732),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[847]),
	.d(FE_OFN292_n250717));
   oa22s01 U263700 (.o(n250716),
	.a(n250732),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[846]),
	.d(FE_OFN292_n250717));
   oa22s01 U263701 (.o(n250719),
	.a(n250732),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[844]),
	.d(FE_OFN563_n250717));
   oa22s01 U263702 (.o(n250720),
	.a(n250732),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[843]),
	.d(FE_OFN563_n250717));
   oa22s01 U263703 (.o(n250721),
	.a(n250732),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[842]),
	.d(FE_OFN292_n250717));
   oa22s01 U263704 (.o(n250722),
	.a(n250732),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[841]),
	.d(FE_OFN292_n250717));
   oa22s01 U263705 (.o(n250724),
	.a(n250732),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[839]),
	.d(FE_OFN563_n250717));
   oa22s01 U263706 (.o(n250726),
	.a(n250732),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[838]),
	.d(FE_OFN292_n250717));
   oa22s01 U263707 (.o(n250734),
	.a(n250768),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[831]),
	.d(FE_OFN294_n250752));
   oa22s01 U263708 (.o(n250735),
	.a(n250768),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[830]),
	.d(FE_OFN294_n250752));
   oa22s01 U263709 (.o(n250736),
	.a(n250768),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[829]),
	.d(FE_OFN294_n250752));
   oa22s01 U263710 (.o(n250737),
	.a(n250768),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[828]),
	.d(FE_OFN294_n250752));
   oa22s01 U263711 (.o(n250738),
	.a(n250768),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[827]),
	.d(FE_OFN294_n250752));
   oa22s01 U263712 (.o(n250739),
	.a(n250768),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[826]),
	.d(FE_OFN294_n250752));
   oa22s01 U263713 (.o(n250741),
	.a(n250768),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[824]),
	.d(FE_OFN294_n250752));
   oa22s01 U263714 (.o(n250742),
	.a(n250768),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[823]),
	.d(FE_OFN294_n250752));
   oa22s01 U263715 (.o(n250743),
	.a(n250768),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[822]),
	.d(FE_OFN294_n250752));
   oa22s01 U263716 (.o(n250744),
	.a(n250768),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[821]),
	.d(FE_OFN294_n250752));
   oa22s01 U263717 (.o(n250745),
	.a(n250768),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[820]),
	.d(FE_OFN294_n250752));
   oa22s01 U263718 (.o(n250746),
	.a(n250768),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[819]),
	.d(FE_OFN294_n250752));
   oa22s01 U263719 (.o(n250747),
	.a(n250768),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[818]),
	.d(FE_OFN294_n250752));
   oa22s01 U263720 (.o(n250748),
	.a(n250768),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[817]),
	.d(FE_OFN294_n250752));
   oa22s01 U263721 (.o(n250749),
	.a(n250768),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[816]),
	.d(FE_OFN294_n250752));
   oa22s01 U263722 (.o(n250750),
	.a(n250768),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[815]),
	.d(FE_OFN294_n250752));
   oa22s01 U263723 (.o(n250751),
	.a(n250768),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[814]),
	.d(FE_OFN294_n250752));
   oa22s01 U263724 (.o(n250753),
	.a(n250768),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[813]),
	.d(FE_OFN294_n250752));
   oa22s01 U263725 (.o(n250754),
	.a(n250768),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[812]),
	.d(FE_OFN294_n250752));
   oa22s01 U263726 (.o(n250755),
	.a(n250768),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[811]),
	.d(FE_OFN294_n250752));
   oa22s01 U263727 (.o(n250757),
	.a(n250768),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[809]),
	.d(FE_OFN294_n250752));
   oa22s01 U263728 (.o(n250758),
	.a(n250768),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[808]),
	.d(FE_OFN294_n250752));
   oa22s01 U263729 (.o(n250759),
	.a(n250768),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[807]),
	.d(FE_OFN294_n250752));
   oa22s01 U263730 (.o(n250761),
	.a(n250768),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[806]),
	.d(FE_OFN294_n250752));
   oa22s01 U263731 (.o(n250771),
	.a(n250804),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[799]),
	.d(FE_OFN296_n250789));
   oa22s01 U263732 (.o(n250772),
	.a(n250804),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[798]),
	.d(FE_OFN296_n250789));
   oa22s01 U263733 (.o(n250773),
	.a(n250804),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[797]),
	.d(FE_OFN296_n250789));
   oa22s01 U263734 (.o(n250774),
	.a(n250804),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[796]),
	.d(FE_OFN296_n250789));
   oa22s01 U263735 (.o(n250776),
	.a(n250804),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[794]),
	.d(FE_OFN296_n250789));
   oa22s01 U263736 (.o(n250777),
	.a(n250804),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[793]),
	.d(FE_OFN296_n250789));
   oa22s01 U263737 (.o(n250778),
	.a(n250804),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[792]),
	.d(FE_OFN296_n250789));
   oa22s01 U263738 (.o(n250779),
	.a(n250804),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[791]),
	.d(FE_OFN296_n250789));
   oa22s01 U263739 (.o(n250780),
	.a(n250804),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[790]),
	.d(FE_OFN296_n250789));
   oa22s01 U263740 (.o(n250781),
	.a(n250804),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[789]),
	.d(FE_OFN296_n250789));
   oa22s01 U263741 (.o(n250782),
	.a(n250804),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[788]),
	.d(FE_OFN296_n250789));
   oa22s01 U263742 (.o(n250783),
	.a(n250804),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[787]),
	.d(FE_OFN296_n250789));
   oa22s01 U263743 (.o(n250784),
	.a(n250804),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[786]),
	.d(FE_OFN296_n250789));
   oa22s01 U263744 (.o(n250785),
	.a(n250804),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[785]),
	.d(FE_OFN296_n250789));
   oa22s01 U263745 (.o(n250786),
	.a(n250804),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[784]),
	.d(FE_OFN296_n250789));
   oa22s01 U263746 (.o(n250787),
	.a(n250804),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[783]),
	.d(FE_OFN296_n250789));
   oa22s01 U263747 (.o(n250788),
	.a(n250804),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[782]),
	.d(FE_OFN296_n250789));
   oa22s01 U263748 (.o(n250790),
	.a(n250804),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[781]),
	.d(FE_OFN296_n250789));
   oa22s01 U263749 (.o(n250792),
	.a(n250804),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[779]),
	.d(FE_OFN296_n250789));
   oa22s01 U263750 (.o(n250793),
	.a(n250804),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[778]),
	.d(FE_OFN296_n250789));
   oa22s01 U263751 (.o(n250794),
	.a(n250804),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[777]),
	.d(FE_OFN296_n250789));
   oa22s01 U263752 (.o(n250795),
	.a(n250804),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[776]),
	.d(FE_OFN296_n250789));
   oa22s01 U263753 (.o(n250796),
	.a(n250804),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[775]),
	.d(FE_OFN296_n250789));
   oa22s01 U263754 (.o(n250798),
	.a(n250804),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[774]),
	.d(FE_OFN296_n250789));
   oa22s01 U263755 (.o(n250806),
	.a(n250839),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[767]),
	.d(n250824));
   oa22s01 U263756 (.o(n250807),
	.a(n250839),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[766]),
	.d(FE_OFN298_n250824));
   oa22s01 U263757 (.o(n250809),
	.a(n250839),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[764]),
	.d(FE_OFN298_n250824));
   oa22s01 U263758 (.o(n250810),
	.a(n250839),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[763]),
	.d(FE_OFN298_n250824));
   oa22s01 U263759 (.o(n250811),
	.a(n250839),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[762]),
	.d(FE_OFN298_n250824));
   oa22s01 U263760 (.o(n250812),
	.a(n250839),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[761]),
	.d(FE_OFN298_n250824));
   oa22s01 U263761 (.o(n250813),
	.a(n250839),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[760]),
	.d(FE_OFN298_n250824));
   oa22s01 U263762 (.o(n250814),
	.a(n250839),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[759]),
	.d(FE_OFN298_n250824));
   oa22s01 U263763 (.o(n250815),
	.a(n250839),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[758]),
	.d(n250824));
   oa22s01 U263764 (.o(n250816),
	.a(n250839),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[757]),
	.d(FE_OFN298_n250824));
   oa22s01 U263765 (.o(n250817),
	.a(n250839),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[756]),
	.d(FE_OFN298_n250824));
   oa22s01 U263766 (.o(n250818),
	.a(n250839),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[755]),
	.d(FE_OFN298_n250824));
   oa22s01 U263767 (.o(n250819),
	.a(n250839),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[754]),
	.d(FE_OFN298_n250824));
   oa22s01 U263768 (.o(n250820),
	.a(n250839),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[753]),
	.d(FE_OFN298_n250824));
   oa22s01 U263769 (.o(n250821),
	.a(n250839),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[752]),
	.d(FE_OFN298_n250824));
   oa22s01 U263770 (.o(n250822),
	.a(n250839),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[751]),
	.d(FE_OFN298_n250824));
   oa22s01 U263771 (.o(n250825),
	.a(n250839),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[749]),
	.d(n250824));
   oa22s01 U263772 (.o(n250826),
	.a(n250839),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[748]),
	.d(FE_OFN298_n250824));
   oa22s01 U263773 (.o(n250827),
	.a(n250839),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[747]),
	.d(FE_OFN298_n250824));
   oa22s01 U263774 (.o(n250829),
	.a(n250839),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[745]),
	.d(n250824));
   oa22s01 U263775 (.o(n250830),
	.a(n250839),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[744]),
	.d(FE_OFN298_n250824));
   oa22s01 U263776 (.o(n250831),
	.a(n250839),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[743]),
	.d(FE_OFN298_n250824));
   oa22s01 U263777 (.o(n250833),
	.a(n250839),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[742]),
	.d(FE_OFN298_n250824));
   oa22s01 U263778 (.o(n250842),
	.a(n250875),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[734]),
	.d(FE_OFN416_n250859));
   oa22s01 U263779 (.o(n250843),
	.a(n250875),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[733]),
	.d(FE_OFN416_n250859));
   oa22s01 U263780 (.o(n250844),
	.a(n250875),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[732]),
	.d(FE_OFN416_n250859));
   oa22s01 U263781 (.o(n250845),
	.a(n250875),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[731]),
	.d(FE_OFN416_n250859));
   oa22s01 U263782 (.o(n250846),
	.a(n250875),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[730]),
	.d(FE_OFN416_n250859));
   oa22s01 U263783 (.o(n250847),
	.a(n250875),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[729]),
	.d(FE_OFN416_n250859));
   oa22s01 U263784 (.o(n250848),
	.a(n250875),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[728]),
	.d(FE_OFN416_n250859));
   oa22s01 U263785 (.o(n250849),
	.a(n250875),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[727]),
	.d(FE_OFN416_n250859));
   oa22s01 U263786 (.o(n250850),
	.a(n250875),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[726]),
	.d(FE_OFN416_n250859));
   oa22s01 U263787 (.o(n250851),
	.a(n250875),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[725]),
	.d(FE_OFN416_n250859));
   oa22s01 U263788 (.o(n250852),
	.a(n250875),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[724]),
	.d(FE_OFN416_n250859));
   oa22s01 U263789 (.o(n250853),
	.a(n250875),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[723]),
	.d(FE_OFN416_n250859));
   oa22s01 U263790 (.o(n250854),
	.a(n250875),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[722]),
	.d(FE_OFN416_n250859));
   oa22s01 U263791 (.o(n250855),
	.a(n250875),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[721]),
	.d(FE_OFN416_n250859));
   oa22s01 U263792 (.o(n250857),
	.a(n250875),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[719]),
	.d(FE_OFN416_n250859));
   oa22s01 U263793 (.o(n250858),
	.a(n250875),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[718]),
	.d(FE_OFN416_n250859));
   oa22s01 U263794 (.o(n250860),
	.a(n250875),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[717]),
	.d(FE_OFN416_n250859));
   oa22s01 U263795 (.o(n250862),
	.a(n250875),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[715]),
	.d(FE_OFN416_n250859));
   oa22s01 U263796 (.o(n250863),
	.a(n250875),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[714]),
	.d(FE_OFN416_n250859));
   oa22s01 U263797 (.o(n250864),
	.a(n250875),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[713]),
	.d(FE_OFN416_n250859));
   oa22s01 U263798 (.o(n250865),
	.a(n250875),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[712]),
	.d(FE_OFN416_n250859));
   oa22s01 U263799 (.o(n250866),
	.a(n250875),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[711]),
	.d(FE_OFN416_n250859));
   oa22s01 U263800 (.o(n250868),
	.a(n250875),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[710]),
	.d(FE_OFN416_n250859));
   oa22s01 U263801 (.o(n250877),
	.a(n250910),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[703]),
	.d(FE_OFN300_n250895));
   oa22s01 U263802 (.o(n250878),
	.a(n250910),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[702]),
	.d(FE_OFN300_n250895));
   oa22s01 U263803 (.o(n250880),
	.a(n250910),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[700]),
	.d(FE_OFN300_n250895));
   oa22s01 U263804 (.o(n250881),
	.a(n250910),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[699]),
	.d(FE_OFN300_n250895));
   oa22s01 U263805 (.o(n250882),
	.a(n250910),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[698]),
	.d(FE_OFN300_n250895));
   oa22s01 U263806 (.o(n250883),
	.a(n250910),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[697]),
	.d(FE_OFN300_n250895));
   oa22s01 U263807 (.o(n250884),
	.a(n250910),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[696]),
	.d(FE_OFN300_n250895));
   oa22s01 U263808 (.o(n250885),
	.a(n250910),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[695]),
	.d(FE_OFN300_n250895));
   oa22s01 U263809 (.o(n250886),
	.a(n250910),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[694]),
	.d(FE_OFN300_n250895));
   oa22s01 U263810 (.o(n250887),
	.a(n250910),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[693]),
	.d(FE_OFN300_n250895));
   oa22s01 U263811 (.o(n250888),
	.a(n250910),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[692]),
	.d(FE_OFN300_n250895));
   oa22s01 U263812 (.o(n250889),
	.a(n250910),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[691]),
	.d(FE_OFN300_n250895));
   oa22s01 U263813 (.o(n250891),
	.a(n250910),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[689]),
	.d(FE_OFN300_n250895));
   oa22s01 U263814 (.o(n250892),
	.a(n250910),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[688]),
	.d(FE_OFN300_n250895));
   oa22s01 U263815 (.o(n250893),
	.a(n250910),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[687]),
	.d(FE_OFN300_n250895));
   oa22s01 U263816 (.o(n250894),
	.a(n250910),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[686]),
	.d(FE_OFN300_n250895));
   oa22s01 U263817 (.o(n250896),
	.a(n250910),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[685]),
	.d(FE_OFN300_n250895));
   oa22s01 U263818 (.o(n250897),
	.a(n250910),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[684]),
	.d(FE_OFN300_n250895));
   oa22s01 U263819 (.o(n250898),
	.a(n250910),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[683]),
	.d(FE_OFN300_n250895));
   oa22s01 U263820 (.o(n250899),
	.a(n250910),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[682]),
	.d(FE_OFN300_n250895));
   oa22s01 U263821 (.o(n250900),
	.a(n250910),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[681]),
	.d(FE_OFN300_n250895));
   oa22s01 U263822 (.o(n250901),
	.a(n250910),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[680]),
	.d(FE_OFN300_n250895));
   oa22s01 U263823 (.o(n250902),
	.a(n250910),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[679]),
	.d(FE_OFN300_n250895));
   oa22s01 U263824 (.o(n250904),
	.a(n250910),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[678]),
	.d(FE_OFN300_n250895));
   oa22s01 U263825 (.o(n250913),
	.a(n250945),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[670]),
	.d(FE_OFN418_n250930));
   oa22s01 U263826 (.o(n250914),
	.a(n250945),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[669]),
	.d(FE_OFN418_n250930));
   oa22s01 U263827 (.o(n250915),
	.a(n250945),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[668]),
	.d(FE_OFN418_n250930));
   oa22s01 U263828 (.o(n250916),
	.a(n250945),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[667]),
	.d(FE_OFN418_n250930));
   oa22s01 U263829 (.o(n250917),
	.a(n250945),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[666]),
	.d(FE_OFN418_n250930));
   oa22s01 U263830 (.o(n250918),
	.a(n250945),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[665]),
	.d(FE_OFN418_n250930));
   oa22s01 U263831 (.o(n250919),
	.a(n250945),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[664]),
	.d(FE_OFN418_n250930));
   oa22s01 U263832 (.o(n250920),
	.a(n250945),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[663]),
	.d(FE_OFN418_n250930));
   oa22s01 U263833 (.o(n250921),
	.a(n250945),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[662]),
	.d(FE_OFN418_n250930));
   oa22s01 U263834 (.o(n250922),
	.a(n250945),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[661]),
	.d(FE_OFN418_n250930));
   oa22s01 U263835 (.o(n250924),
	.a(n250945),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[659]),
	.d(FE_OFN418_n250930));
   oa22s01 U263836 (.o(n250925),
	.a(n250945),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[658]),
	.d(FE_OFN418_n250930));
   oa22s01 U263837 (.o(n250926),
	.a(n250945),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[657]),
	.d(FE_OFN418_n250930));
   oa22s01 U263838 (.o(n250927),
	.a(n250945),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[656]),
	.d(FE_OFN418_n250930));
   oa22s01 U263839 (.o(n250928),
	.a(n250945),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[655]),
	.d(FE_OFN418_n250930));
   oa22s01 U263840 (.o(n250929),
	.a(n250945),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[654]),
	.d(FE_OFN418_n250930));
   oa22s01 U263841 (.o(n250931),
	.a(n250945),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[653]),
	.d(FE_OFN418_n250930));
   oa22s01 U263842 (.o(n250932),
	.a(n250945),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[652]),
	.d(FE_OFN418_n250930));
   oa22s01 U263843 (.o(n250933),
	.a(n250945),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[651]),
	.d(FE_OFN418_n250930));
   oa22s01 U263844 (.o(n250934),
	.a(n250945),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[650]),
	.d(FE_OFN418_n250930));
   oa22s01 U263845 (.o(n250935),
	.a(n250945),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[649]),
	.d(FE_OFN418_n250930));
   oa22s01 U263846 (.o(n250936),
	.a(n250945),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[648]),
	.d(FE_OFN418_n250930));
   oa22s01 U263847 (.o(n250937),
	.a(n250945),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[647]),
	.d(FE_OFN418_n250930));
   oa22s01 U263848 (.o(n250939),
	.a(n250945),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[646]),
	.d(FE_OFN418_n250930));
   oa22s01 U263849 (.o(n250947),
	.a(n250981),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[639]),
	.d(FE_OFN200_n250965));
   oa22s01 U263850 (.o(n250948),
	.a(n250981),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[638]),
	.d(FE_OFN200_n250965));
   oa22s01 U263851 (.o(n250949),
	.a(n250981),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[637]),
	.d(FE_OFN200_n250965));
   oa22s01 U263852 (.o(n250950),
	.a(n250981),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[636]),
	.d(FE_OFN200_n250965));
   oa22s01 U263853 (.o(n250951),
	.a(n250981),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[635]),
	.d(FE_OFN200_n250965));
   oa22s01 U263854 (.o(n250952),
	.a(n250981),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[634]),
	.d(FE_OFN200_n250965));
   oa22s01 U263855 (.o(n250953),
	.a(n250981),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[633]),
	.d(FE_OFN200_n250965));
   oa22s01 U263856 (.o(n250954),
	.a(n250981),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[632]),
	.d(FE_OFN200_n250965));
   oa22s01 U263857 (.o(n250955),
	.a(n250981),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[631]),
	.d(FE_OFN200_n250965));
   oa22s01 U263858 (.o(n250957),
	.a(n250981),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[629]),
	.d(FE_OFN200_n250965));
   oa22s01 U263859 (.o(n250958),
	.a(n250981),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[628]),
	.d(FE_OFN200_n250965));
   oa22s01 U263860 (.o(n250959),
	.a(n250981),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[627]),
	.d(FE_OFN200_n250965));
   oa22s01 U263861 (.o(n250960),
	.a(n250981),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[626]),
	.d(FE_OFN200_n250965));
   oa22s01 U263862 (.o(n250961),
	.a(n250981),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[625]),
	.d(FE_OFN200_n250965));
   oa22s01 U263863 (.o(n250962),
	.a(n250981),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[624]),
	.d(FE_OFN200_n250965));
   oa22s01 U263864 (.o(n250963),
	.a(n250981),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[623]),
	.d(FE_OFN200_n250965));
   oa22s01 U263865 (.o(n250964),
	.a(n250981),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[622]),
	.d(FE_OFN200_n250965));
   oa22s01 U263866 (.o(n250966),
	.a(n250981),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[621]),
	.d(FE_OFN200_n250965));
   oa22s01 U263867 (.o(n250967),
	.a(n250981),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[620]),
	.d(FE_OFN200_n250965));
   oa22s01 U263868 (.o(n250968),
	.a(n250981),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[619]),
	.d(FE_OFN200_n250965));
   oa22s01 U263869 (.o(n250969),
	.a(n250981),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[618]),
	.d(FE_OFN200_n250965));
   oa22s01 U263870 (.o(n250970),
	.a(n250981),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[617]),
	.d(FE_OFN200_n250965));
   oa22s01 U263871 (.o(n250971),
	.a(n250981),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[616]),
	.d(FE_OFN200_n250965));
   oa22s01 U263872 (.o(n250974),
	.a(n250981),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[614]),
	.d(FE_OFN200_n250965));
   oa22s01 U263873 (.o(n250988),
	.a(n251016),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[602]),
	.d(FE_OFN302_n251001));
   oa22s01 U263874 (.o(n250992),
	.a(n251016),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[598]),
	.d(FE_OFN302_n251001));
   oa22s01 U263875 (.o(n250994),
	.a(n251016),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[596]),
	.d(FE_OFN302_n251001));
   oa22s01 U263876 (.o(n250996),
	.a(n251016),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[594]),
	.d(FE_OFN302_n251001));
   oa22s01 U263877 (.o(n250999),
	.a(n251016),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[591]),
	.d(FE_OFN302_n251001));
   oa22s01 U263878 (.o(n251000),
	.a(n251016),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[590]),
	.d(FE_OFN302_n251001));
   oa22s01 U263879 (.o(n251007),
	.a(n251016),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[584]),
	.d(FE_OFN302_n251001));
   oa22s01 U263880 (.o(n251008),
	.a(n251016),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[583]),
	.d(FE_OFN302_n251001));
   oa22s01 U263881 (.o(n251010),
	.a(n251016),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[582]),
	.d(FE_OFN302_n251001));
   oa22s01 U263882 (.o(n251018),
	.a(n251051),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[575]),
	.d(FE_OFN304_n251036));
   oa22s01 U263883 (.o(n251019),
	.a(n251051),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[574]),
	.d(FE_OFN304_n251036));
   oa22s01 U263884 (.o(n251020),
	.a(n251051),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[573]),
	.d(FE_OFN304_n251036));
   oa22s01 U263885 (.o(n251021),
	.a(n251051),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[572]),
	.d(FE_OFN304_n251036));
   oa22s01 U263886 (.o(n251022),
	.a(n251051),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[571]),
	.d(FE_OFN304_n251036));
   oa22s01 U263887 (.o(n251024),
	.a(n251051),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[569]),
	.d(FE_OFN304_n251036));
   oa22s01 U263888 (.o(n251025),
	.a(n251051),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[568]),
	.d(FE_OFN304_n251036));
   oa22s01 U263889 (.o(n251026),
	.a(n251051),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[567]),
	.d(FE_OFN304_n251036));
   oa22s01 U263890 (.o(n251027),
	.a(n251051),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[566]),
	.d(FE_OFN304_n251036));
   oa22s01 U263891 (.o(n251028),
	.a(n251051),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[565]),
	.d(FE_OFN304_n251036));
   oa22s01 U263892 (.o(n251029),
	.a(n251051),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[564]),
	.d(FE_OFN304_n251036));
   oa22s01 U263893 (.o(n251030),
	.a(n251051),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[563]),
	.d(FE_OFN304_n251036));
   oa22s01 U263894 (.o(n251031),
	.a(n251051),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[562]),
	.d(FE_OFN304_n251036));
   oa22s01 U263895 (.o(n251032),
	.a(n251051),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[561]),
	.d(FE_OFN304_n251036));
   oa22s01 U263896 (.o(n251033),
	.a(n251051),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[560]),
	.d(FE_OFN304_n251036));
   oa22s01 U263897 (.o(n251034),
	.a(n251051),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[559]),
	.d(FE_OFN304_n251036));
   oa22s01 U263898 (.o(n251035),
	.a(n251051),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[558]),
	.d(FE_OFN304_n251036));
   oa22s01 U263899 (.o(n251037),
	.a(n251051),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[557]),
	.d(FE_OFN304_n251036));
   oa22s01 U263900 (.o(n251038),
	.a(n251051),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[556]),
	.d(FE_OFN304_n251036));
   oa22s01 U263901 (.o(n251040),
	.a(n251051),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[554]),
	.d(FE_OFN304_n251036));
   oa22s01 U263902 (.o(n251041),
	.a(n251051),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[553]),
	.d(FE_OFN304_n251036));
   oa22s01 U263903 (.o(n251042),
	.a(n251051),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[552]),
	.d(FE_OFN304_n251036));
   oa22s01 U263904 (.o(n251043),
	.a(n251051),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[551]),
	.d(FE_OFN304_n251036));
   oa22s01 U263905 (.o(n251045),
	.a(n251051),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[550]),
	.d(FE_OFN304_n251036));
   oa22s01 U263906 (.o(n251054),
	.a(n251088),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[543]),
	.d(FE_OFN307_n251072));
   oa22s01 U263907 (.o(n251055),
	.a(n251088),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[542]),
	.d(FE_OFN307_n251072));
   oa22s01 U263908 (.o(n251056),
	.a(n251088),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[541]),
	.d(FE_OFN306_n251072));
   oa22s01 U263909 (.o(n251058),
	.a(n251088),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[539]),
	.d(FE_OFN306_n251072));
   oa22s01 U263910 (.o(n251059),
	.a(n251088),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[538]),
	.d(FE_OFN307_n251072));
   oa22s01 U263911 (.o(n251060),
	.a(n251088),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[537]),
	.d(FE_OFN307_n251072));
   oa22s01 U263912 (.o(n251061),
	.a(n251088),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[536]),
	.d(FE_OFN306_n251072));
   oa22s01 U263913 (.o(n251062),
	.a(n251088),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[535]),
	.d(FE_OFN306_n251072));
   oa22s01 U263914 (.o(n251063),
	.a(n251088),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[534]),
	.d(FE_OFN307_n251072));
   oa22s01 U263915 (.o(n251064),
	.a(n251088),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[533]),
	.d(FE_OFN307_n251072));
   oa22s01 U263916 (.o(n251065),
	.a(n251088),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[532]),
	.d(FE_OFN307_n251072));
   oa22s01 U263917 (.o(n251066),
	.a(n251088),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[531]),
	.d(FE_OFN307_n251072));
   oa22s01 U263918 (.o(n251067),
	.a(n251088),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[530]),
	.d(FE_OFN307_n251072));
   oa22s01 U263919 (.o(n251068),
	.a(n251088),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[529]),
	.d(FE_OFN307_n251072));
   oa22s01 U263920 (.o(n251069),
	.a(n251088),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[528]),
	.d(FE_OFN307_n251072));
   oa22s01 U263921 (.o(n251070),
	.a(n251088),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[527]),
	.d(FE_OFN306_n251072));
   oa22s01 U263922 (.o(n251071),
	.a(n251088),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[526]),
	.d(FE_OFN306_n251072));
   oa22s01 U263923 (.o(n251074),
	.a(n251088),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[524]),
	.d(FE_OFN307_n251072));
   oa22s01 U263924 (.o(n251075),
	.a(n251088),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[523]),
	.d(FE_OFN307_n251072));
   oa22s01 U263925 (.o(n251076),
	.a(n251088),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[522]),
	.d(FE_OFN306_n251072));
   oa22s01 U263926 (.o(n251078),
	.a(n251088),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[520]),
	.d(FE_OFN307_n251072));
   oa22s01 U263927 (.o(n251079),
	.a(n251088),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[519]),
	.d(FE_OFN306_n251072));
   oa22s01 U263928 (.o(n251081),
	.a(n251088),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[518]),
	.d(FE_OFN306_n251072));
   oa22s01 U263929 (.o(n251090),
	.a(n251123),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1535]),
	.d(FE_OFN309_n251105));
   oa22s01 U263930 (.o(n251092),
	.a(n251123),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1533]),
	.d(FE_OFN309_n251105));
   oa22s01 U263931 (.o(n251093),
	.a(n251123),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1532]),
	.d(FE_OFN309_n251105));
   oa22s01 U263932 (.o(n251094),
	.a(n251123),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1531]),
	.d(FE_OFN309_n251105));
   oa22s01 U263933 (.o(n251095),
	.a(n251123),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1530]),
	.d(n251105));
   oa22s01 U263934 (.o(n251096),
	.a(n251123),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1529]),
	.d(FE_OFN309_n251105));
   oa22s01 U263935 (.o(n251097),
	.a(n251123),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1528]),
	.d(FE_OFN309_n251105));
   oa22s01 U263936 (.o(n251098),
	.a(n251123),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1527]),
	.d(FE_OFN309_n251105));
   oa22s01 U263937 (.o(n251099),
	.a(n251123),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1526]),
	.d(FE_OFN309_n251105));
   oa22s01 U263938 (.o(n251100),
	.a(n251123),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1525]),
	.d(FE_OFN309_n251105));
   oa22s01 U263939 (.o(n251101),
	.a(n251123),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1524]),
	.d(FE_OFN309_n251105));
   oa22s01 U263940 (.o(n251102),
	.a(n251123),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1523]),
	.d(FE_OFN309_n251105));
   oa22s01 U263941 (.o(n251103),
	.a(n251123),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1522]),
	.d(n251105));
   oa22s01 U263942 (.o(n251104),
	.a(n251123),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1521]),
	.d(FE_OFN309_n251105));
   oa22s01 U263943 (.o(n251106),
	.a(n251123),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1520]),
	.d(FE_OFN309_n251105));
   oa22s01 U263944 (.o(n251108),
	.a(n251123),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1518]),
	.d(FE_OFN309_n251105));
   oa22s01 U263945 (.o(n251109),
	.a(n251123),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1517]),
	.d(FE_OFN309_n251105));
   oa22s01 U263946 (.o(n251110),
	.a(n251123),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1516]),
	.d(n251105));
   oa22s01 U263947 (.o(n251112),
	.a(n251123),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1514]),
	.d(FE_OFN309_n251105));
   oa22s01 U263948 (.o(n251113),
	.a(n251123),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1513]),
	.d(FE_OFN309_n251105));
   oa22s01 U263949 (.o(n251114),
	.a(n251123),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1512]),
	.d(FE_OFN309_n251105));
   oa22s01 U263950 (.o(n251115),
	.a(n251123),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1511]),
	.d(FE_OFN309_n251105));
   oa22s01 U263951 (.o(n251117),
	.a(n251123),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1510]),
	.d(FE_OFN309_n251105));
   oa22s01 U263952 (.o(n251125),
	.a(n251158),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1503]),
	.d(FE_OFN420_n251140));
   oa22s01 U263953 (.o(n251126),
	.a(n251158),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1502]),
	.d(FE_OFN420_n251140));
   oa22s01 U263954 (.o(n251127),
	.a(n251158),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1501]),
	.d(FE_OFN420_n251140));
   oa22s01 U263955 (.o(n251128),
	.a(n251158),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1500]),
	.d(FE_OFN420_n251140));
   oa22s01 U263956 (.o(n251129),
	.a(n251158),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1499]),
	.d(FE_OFN420_n251140));
   oa22s01 U263957 (.o(n251130),
	.a(n251158),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1498]),
	.d(FE_OFN420_n251140));
   oa22s01 U263958 (.o(n251131),
	.a(n251158),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1497]),
	.d(FE_OFN420_n251140));
   oa22s01 U263959 (.o(n251132),
	.a(n251158),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1496]),
	.d(FE_OFN420_n251140));
   oa22s01 U263960 (.o(n251133),
	.a(n251158),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1495]),
	.d(FE_OFN420_n251140));
   oa22s01 U263961 (.o(n251134),
	.a(n251158),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1494]),
	.d(FE_OFN420_n251140));
   oa22s01 U263962 (.o(n251135),
	.a(n251158),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1493]),
	.d(FE_OFN420_n251140));
   oa22s01 U263963 (.o(n251136),
	.a(n251158),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1492]),
	.d(FE_OFN420_n251140));
   oa22s01 U263964 (.o(n251137),
	.a(n251158),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1491]),
	.d(FE_OFN420_n251140));
   oa22s01 U263965 (.o(n251138),
	.a(n251158),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1490]),
	.d(FE_OFN420_n251140));
   oa22s01 U263966 (.o(n251141),
	.a(n251158),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1488]),
	.d(FE_OFN420_n251140));
   oa22s01 U263967 (.o(n251142),
	.a(n251158),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1487]),
	.d(FE_OFN420_n251140));
   oa22s01 U263968 (.o(n251143),
	.a(n251158),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1486]),
	.d(FE_OFN420_n251140));
   oa22s01 U263969 (.o(n251145),
	.a(n251158),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1484]),
	.d(FE_OFN420_n251140));
   oa22s01 U263970 (.o(n251146),
	.a(n251158),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1483]),
	.d(FE_OFN420_n251140));
   oa22s01 U263971 (.o(n251147),
	.a(n251158),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1482]),
	.d(FE_OFN420_n251140));
   oa22s01 U263972 (.o(n251148),
	.a(n251158),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1481]),
	.d(FE_OFN420_n251140));
   oa22s01 U263973 (.o(n251149),
	.a(n251158),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1480]),
	.d(FE_OFN420_n251140));
   oa22s01 U263974 (.o(n251150),
	.a(n251158),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1479]),
	.d(FE_OFN420_n251140));
   oa22s01 U263975 (.o(n251152),
	.a(n251158),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1478]),
	.d(FE_OFN420_n251140));
   oa22s01 U263976 (.o(n251160),
	.a(n251194),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1471]),
	.d(FE_OFN311_n251175));
   oa22s01 U263977 (.o(n251162),
	.a(n251194),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1469]),
	.d(FE_OFN311_n251175));
   oa22s01 U263978 (.o(n251163),
	.a(n251194),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1468]),
	.d(FE_OFN311_n251175));
   oa22s01 U263979 (.o(n251164),
	.a(n251194),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1467]),
	.d(FE_OFN311_n251175));
   oa22s01 U263980 (.o(n251165),
	.a(n251194),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1466]),
	.d(FE_OFN311_n251175));
   oa22s01 U263981 (.o(n251166),
	.a(n251194),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1465]),
	.d(FE_OFN311_n251175));
   oa22s01 U263982 (.o(n251167),
	.a(n251194),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1464]),
	.d(FE_OFN311_n251175));
   oa22s01 U263983 (.o(n251168),
	.a(n251194),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1463]),
	.d(FE_OFN311_n251175));
   oa22s01 U263984 (.o(n251169),
	.a(n251194),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1462]),
	.d(FE_OFN311_n251175));
   oa22s01 U263985 (.o(n251170),
	.a(n251194),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1461]),
	.d(FE_OFN311_n251175));
   oa22s01 U263986 (.o(n251171),
	.a(n251194),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1460]),
	.d(FE_OFN311_n251175));
   oa22s01 U263987 (.o(n251173),
	.a(n251194),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1458]),
	.d(FE_OFN311_n251175));
   oa22s01 U263988 (.o(n251174),
	.a(n251194),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1457]),
	.d(FE_OFN311_n251175));
   oa22s01 U263989 (.o(n251176),
	.a(n251194),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1456]),
	.d(FE_OFN311_n251175));
   oa22s01 U263990 (.o(n251177),
	.a(n251194),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1455]),
	.d(FE_OFN311_n251175));
   oa22s01 U263991 (.o(n251178),
	.a(n251194),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1454]),
	.d(FE_OFN311_n251175));
   oa22s01 U263992 (.o(n251179),
	.a(n251194),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1453]),
	.d(FE_OFN311_n251175));
   oa22s01 U263993 (.o(n251180),
	.a(n251194),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1452]),
	.d(FE_OFN311_n251175));
   oa22s01 U263994 (.o(n251181),
	.a(n251194),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1451]),
	.d(FE_OFN311_n251175));
   oa22s01 U263995 (.o(n251182),
	.a(n251194),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1450]),
	.d(FE_OFN311_n251175));
   oa22s01 U263996 (.o(n251183),
	.a(n251194),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1449]),
	.d(FE_OFN311_n251175));
   oa22s01 U263997 (.o(n251184),
	.a(n251194),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1448]),
	.d(FE_OFN311_n251175));
   oa22s01 U263998 (.o(n251185),
	.a(n251194),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1447]),
	.d(FE_OFN311_n251175));
   oa22s01 U263999 (.o(n251187),
	.a(n251194),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1446]),
	.d(FE_OFN311_n251175));
   oa22s01 U264000 (.o(n251231),
	.a(n251264),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1407]),
	.d(FE_OFN202_n251246));
   oa22s01 U264001 (.o(n251232),
	.a(n251264),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1406]),
	.d(FE_OFN202_n251246));
   oa22s01 U264002 (.o(n251233),
	.a(n251264),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1405]),
	.d(FE_OFN202_n251246));
   oa22s01 U264003 (.o(n251234),
	.a(n251264),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1404]),
	.d(FE_OFN202_n251246));
   oa22s01 U264004 (.o(n251235),
	.a(n251264),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1403]),
	.d(FE_OFN202_n251246));
   oa22s01 U264005 (.o(n251236),
	.a(n251264),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1402]),
	.d(FE_OFN202_n251246));
   oa22s01 U264006 (.o(n251237),
	.a(n251264),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1401]),
	.d(FE_OFN202_n251246));
   oa22s01 U264007 (.o(n251238),
	.a(n251264),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1400]),
	.d(FE_OFN202_n251246));
   oa22s01 U264008 (.o(n251240),
	.a(n251264),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1398]),
	.d(FE_OFN202_n251246));
   oa22s01 U264009 (.o(n251241),
	.a(n251264),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1397]),
	.d(FE_OFN202_n251246));
   oa22s01 U264010 (.o(n251242),
	.a(n251264),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1396]),
	.d(FE_OFN202_n251246));
   oa22s01 U264011 (.o(n251243),
	.a(n251264),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1395]),
	.d(FE_OFN202_n251246));
   oa22s01 U264012 (.o(n251244),
	.a(n251264),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1394]),
	.d(FE_OFN202_n251246));
   oa22s01 U264013 (.o(n251245),
	.a(n251264),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1393]),
	.d(FE_OFN202_n251246));
   oa22s01 U264014 (.o(n251247),
	.a(n251264),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1392]),
	.d(FE_OFN202_n251246));
   oa22s01 U264015 (.o(n251248),
	.a(n251264),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1391]),
	.d(FE_OFN202_n251246));
   oa22s01 U264016 (.o(n251249),
	.a(n251264),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1390]),
	.d(FE_OFN202_n251246));
   oa22s01 U264017 (.o(n251250),
	.a(n251264),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1389]),
	.d(FE_OFN202_n251246));
   oa22s01 U264018 (.o(n251251),
	.a(n251264),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1388]),
	.d(FE_OFN202_n251246));
   oa22s01 U264019 (.o(n251252),
	.a(n251264),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1387]),
	.d(FE_OFN202_n251246));
   oa22s01 U264020 (.o(n251253),
	.a(n251264),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1386]),
	.d(FE_OFN202_n251246));
   oa22s01 U264021 (.o(n251254),
	.a(n251264),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1385]),
	.d(FE_OFN202_n251246));
   oa22s01 U264022 (.o(n251256),
	.a(n251264),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1383]),
	.d(FE_OFN202_n251246));
   oa22s01 U264023 (.o(n251258),
	.a(n251264),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1382]),
	.d(FE_OFN202_n251246));
   oa22s01 U264024 (.o(n251302),
	.a(n251335),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1343]),
	.d(FE_OFN316_n251317));
   oa22s01 U264025 (.o(n251303),
	.a(n251335),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1342]),
	.d(FE_OFN316_n251317));
   oa22s01 U264026 (.o(n251304),
	.a(n251335),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1341]),
	.d(FE_OFN316_n251317));
   oa22s01 U264027 (.o(n251305),
	.a(n251335),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1340]),
	.d(FE_OFN316_n251317));
   oa22s01 U264028 (.o(n251307),
	.a(n251335),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1338]),
	.d(FE_OFN316_n251317));
   oa22s01 U264029 (.o(n251308),
	.a(n251335),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1337]),
	.d(FE_OFN316_n251317));
   oa22s01 U264030 (.o(n251309),
	.a(n251335),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1336]),
	.d(FE_OFN316_n251317));
   oa22s01 U264031 (.o(n251310),
	.a(n251335),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1335]),
	.d(FE_OFN316_n251317));
   oa22s01 U264032 (.o(n251311),
	.a(n251335),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1334]),
	.d(FE_OFN316_n251317));
   oa22s01 U264033 (.o(n251312),
	.a(n251335),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1333]),
	.d(FE_OFN316_n251317));
   oa22s01 U264034 (.o(n251313),
	.a(n251335),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1332]),
	.d(FE_OFN316_n251317));
   oa22s01 U264035 (.o(n251314),
	.a(n251335),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1331]),
	.d(FE_OFN316_n251317));
   oa22s01 U264036 (.o(n251315),
	.a(n251335),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1330]),
	.d(FE_OFN316_n251317));
   oa22s01 U264037 (.o(n251316),
	.a(n251335),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1329]),
	.d(FE_OFN316_n251317));
   oa22s01 U264038 (.o(n251318),
	.a(n251335),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1328]),
	.d(FE_OFN316_n251317));
   oa22s01 U264039 (.o(n251319),
	.a(n251335),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1327]),
	.d(FE_OFN316_n251317));
   oa22s01 U264040 (.o(n251320),
	.a(n251335),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1326]),
	.d(FE_OFN316_n251317));
   oa22s01 U264041 (.o(n251321),
	.a(n251335),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1325]),
	.d(FE_OFN316_n251317));
   oa22s01 U264042 (.o(n251323),
	.a(n251335),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1323]),
	.d(FE_OFN316_n251317));
   oa22s01 U264043 (.o(n251324),
	.a(n251335),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1322]),
	.d(FE_OFN316_n251317));
   oa22s01 U264044 (.o(n251325),
	.a(n251335),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1321]),
	.d(FE_OFN316_n251317));
   oa22s01 U264045 (.o(n251326),
	.a(n251335),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1320]),
	.d(FE_OFN316_n251317));
   oa22s01 U264046 (.o(n251327),
	.a(n251335),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1319]),
	.d(FE_OFN316_n251317));
   oa22s01 U264047 (.o(n251329),
	.a(n251335),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1318]),
	.d(FE_OFN316_n251317));
   oa22s01 U264048 (.o(n251338),
	.a(n251371),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1311]),
	.d(FE_OFN318_n251353));
   oa22s01 U264049 (.o(n251339),
	.a(n251371),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1310]),
	.d(FE_OFN318_n251353));
   oa22s01 U264050 (.o(n251341),
	.a(n251371),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1308]),
	.d(FE_OFN318_n251353));
   oa22s01 U264051 (.o(n251342),
	.a(n251371),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1307]),
	.d(FE_OFN318_n251353));
   oa22s01 U264052 (.o(n251343),
	.a(n251371),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1306]),
	.d(FE_OFN318_n251353));
   oa22s01 U264053 (.o(n251344),
	.a(n251371),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1305]),
	.d(FE_OFN318_n251353));
   oa22s01 U264054 (.o(n251345),
	.a(n251371),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1304]),
	.d(FE_OFN318_n251353));
   oa22s01 U264055 (.o(n251346),
	.a(n251371),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1303]),
	.d(FE_OFN318_n251353));
   oa22s01 U264056 (.o(n251347),
	.a(n251371),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1302]),
	.d(FE_OFN318_n251353));
   oa22s01 U264057 (.o(n251348),
	.a(n251371),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1301]),
	.d(FE_OFN318_n251353));
   oa22s01 U264058 (.o(n251349),
	.a(n251371),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1300]),
	.d(FE_OFN318_n251353));
   oa22s01 U264059 (.o(n251350),
	.a(n251371),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1299]),
	.d(FE_OFN318_n251353));
   oa22s01 U264060 (.o(n251351),
	.a(n251371),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1298]),
	.d(FE_OFN318_n251353));
   oa22s01 U264061 (.o(n251352),
	.a(n251371),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1297]),
	.d(FE_OFN318_n251353));
   oa22s01 U264062 (.o(n251354),
	.a(n251371),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1296]),
	.d(FE_OFN318_n251353));
   oa22s01 U264063 (.o(n251355),
	.a(n251371),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1295]),
	.d(FE_OFN318_n251353));
   oa22s01 U264064 (.o(n251357),
	.a(n251371),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1293]),
	.d(FE_OFN318_n251353));
   oa22s01 U264065 (.o(n251358),
	.a(n251371),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1292]),
	.d(FE_OFN318_n251353));
   oa22s01 U264066 (.o(n251359),
	.a(n251371),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1291]),
	.d(FE_OFN318_n251353));
   oa22s01 U264067 (.o(n251361),
	.a(n251371),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1289]),
	.d(FE_OFN318_n251353));
   oa22s01 U264068 (.o(n251362),
	.a(n251371),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1288]),
	.d(FE_OFN318_n251353));
   oa22s01 U264069 (.o(n251363),
	.a(n251371),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1287]),
	.d(FE_OFN318_n251353));
   oa22s01 U264070 (.o(n251365),
	.a(n251371),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1286]),
	.d(FE_OFN318_n251353));
   oa22s01 U264071 (.o(n251374),
	.a(n251407),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1278]),
	.d(FE_OFN320_n251388));
   oa22s01 U264072 (.o(n251375),
	.a(n251407),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1277]),
	.d(FE_OFN320_n251388));
   oa22s01 U264073 (.o(n251376),
	.a(n251407),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1276]),
	.d(FE_OFN320_n251388));
   oa22s01 U264074 (.o(n251377),
	.a(n251407),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1275]),
	.d(FE_OFN320_n251388));
   oa22s01 U264075 (.o(n251378),
	.a(n251407),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1274]),
	.d(FE_OFN320_n251388));
   oa22s01 U264076 (.o(n251379),
	.a(n251407),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1273]),
	.d(FE_OFN320_n251388));
   oa22s01 U264077 (.o(n251380),
	.a(n251407),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1272]),
	.d(FE_OFN320_n251388));
   oa22s01 U264078 (.o(n251381),
	.a(n251407),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1271]),
	.d(FE_OFN320_n251388));
   oa22s01 U264079 (.o(n251382),
	.a(n251407),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1270]),
	.d(FE_OFN320_n251388));
   oa22s01 U264080 (.o(n251383),
	.a(n251407),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1269]),
	.d(FE_OFN320_n251388));
   oa22s01 U264081 (.o(n251384),
	.a(n251407),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1268]),
	.d(FE_OFN320_n251388));
   oa22s01 U264082 (.o(n251385),
	.a(n251407),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1267]),
	.d(FE_OFN320_n251388));
   oa22s01 U264083 (.o(n251386),
	.a(n251407),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1266]),
	.d(FE_OFN320_n251388));
   oa22s01 U264084 (.o(n251387),
	.a(n251407),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1265]),
	.d(FE_OFN320_n251388));
   oa22s01 U264085 (.o(n251390),
	.a(n251407),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1263]),
	.d(FE_OFN320_n251388));
   oa22s01 U264086 (.o(n251391),
	.a(n251407),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1262]),
	.d(FE_OFN320_n251388));
   oa22s01 U264087 (.o(n251392),
	.a(n251407),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1261]),
	.d(FE_OFN320_n251388));
   oa22s01 U264088 (.o(n251394),
	.a(n251407),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1259]),
	.d(FE_OFN320_n251388));
   oa22s01 U264089 (.o(n251395),
	.a(n251407),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1258]),
	.d(FE_OFN320_n251388));
   oa22s01 U264090 (.o(n251396),
	.a(n251407),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1257]),
	.d(FE_OFN320_n251388));
   oa22s01 U264091 (.o(n251397),
	.a(n251407),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1256]),
	.d(FE_OFN320_n251388));
   oa22s01 U264092 (.o(n251398),
	.a(n251407),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1255]),
	.d(FE_OFN320_n251388));
   oa22s01 U264093 (.o(n251400),
	.a(n251407),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1254]),
	.d(FE_OFN320_n251388));
   oa22s01 U264094 (.o(n251409),
	.a(n251442),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1247]),
	.d(FE_OFN426_n251424));
   oa22s01 U264095 (.o(n251410),
	.a(n251442),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1246]),
	.d(FE_OFN426_n251424));
   oa22s01 U264096 (.o(n251412),
	.a(n251442),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1244]),
	.d(FE_OFN426_n251424));
   oa22s01 U264097 (.o(n251413),
	.a(n251442),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1243]),
	.d(FE_OFN426_n251424));
   oa22s01 U264098 (.o(n251414),
	.a(n251442),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1242]),
	.d(FE_OFN426_n251424));
   oa22s01 U264099 (.o(n251415),
	.a(n251442),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1241]),
	.d(FE_OFN426_n251424));
   oa22s01 U264100 (.o(n251416),
	.a(n251442),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1240]),
	.d(FE_OFN426_n251424));
   oa22s01 U264101 (.o(n251417),
	.a(n251442),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1239]),
	.d(FE_OFN426_n251424));
   oa22s01 U264102 (.o(n251418),
	.a(n251442),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1238]),
	.d(FE_OFN426_n251424));
   oa22s01 U264103 (.o(n251419),
	.a(n251442),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1237]),
	.d(FE_OFN426_n251424));
   oa22s01 U264104 (.o(n251420),
	.a(n251442),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1236]),
	.d(FE_OFN426_n251424));
   oa22s01 U264105 (.o(n251421),
	.a(n251442),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1235]),
	.d(FE_OFN426_n251424));
   oa22s01 U264106 (.o(n251423),
	.a(n251442),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1233]),
	.d(FE_OFN426_n251424));
   oa22s01 U264107 (.o(n251425),
	.a(n251442),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1232]),
	.d(FE_OFN426_n251424));
   oa22s01 U264108 (.o(n251426),
	.a(n251442),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1231]),
	.d(FE_OFN426_n251424));
   oa22s01 U264109 (.o(n251427),
	.a(n251442),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1230]),
	.d(FE_OFN426_n251424));
   oa22s01 U264110 (.o(n251428),
	.a(n251442),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1229]),
	.d(FE_OFN426_n251424));
   oa22s01 U264111 (.o(n251429),
	.a(n251442),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1228]),
	.d(FE_OFN426_n251424));
   oa22s01 U264112 (.o(n251430),
	.a(n251442),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1227]),
	.d(FE_OFN426_n251424));
   oa22s01 U264113 (.o(n251431),
	.a(n251442),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1226]),
	.d(FE_OFN426_n251424));
   oa22s01 U264114 (.o(n251432),
	.a(n251442),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1225]),
	.d(FE_OFN426_n251424));
   oa22s01 U264115 (.o(n251433),
	.a(n251442),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1224]),
	.d(FE_OFN426_n251424));
   oa22s01 U264116 (.o(n251434),
	.a(n251442),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1223]),
	.d(FE_OFN426_n251424));
   oa22s01 U264117 (.o(n251436),
	.a(n251442),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1222]),
	.d(FE_OFN426_n251424));
   oa22s01 U264118 (.o(n251445),
	.a(n251477),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1214]),
	.d(FE_OFN322_n251459));
   oa22s01 U264119 (.o(n251446),
	.a(n251477),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1213]),
	.d(FE_OFN322_n251459));
   oa22s01 U264120 (.o(n251447),
	.a(n251477),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1212]),
	.d(FE_OFN322_n251459));
   oa22s01 U264121 (.o(n251448),
	.a(n251477),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1211]),
	.d(FE_OFN322_n251459));
   oa22s01 U264122 (.o(n251449),
	.a(n251477),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1210]),
	.d(FE_OFN322_n251459));
   oa22s01 U264123 (.o(n251450),
	.a(n251477),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1209]),
	.d(FE_OFN322_n251459));
   oa22s01 U264124 (.o(n251451),
	.a(n251477),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1208]),
	.d(FE_OFN322_n251459));
   oa22s01 U264125 (.o(n251452),
	.a(n251477),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1207]),
	.d(FE_OFN322_n251459));
   oa22s01 U264126 (.o(n251453),
	.a(n251477),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1206]),
	.d(FE_OFN322_n251459));
   oa22s01 U264127 (.o(n251454),
	.a(n251477),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1205]),
	.d(FE_OFN322_n251459));
   oa22s01 U264128 (.o(n251456),
	.a(n251477),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1203]),
	.d(FE_OFN322_n251459));
   oa22s01 U264129 (.o(n251457),
	.a(n251477),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1202]),
	.d(FE_OFN322_n251459));
   oa22s01 U264130 (.o(n251458),
	.a(n251477),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1201]),
	.d(FE_OFN322_n251459));
   oa22s01 U264131 (.o(n251460),
	.a(n251477),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1200]),
	.d(FE_OFN322_n251459));
   oa22s01 U264132 (.o(n251461),
	.a(n251477),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1199]),
	.d(FE_OFN322_n251459));
   oa22s01 U264133 (.o(n251462),
	.a(n251477),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1198]),
	.d(FE_OFN322_n251459));
   oa22s01 U264134 (.o(n251463),
	.a(n251477),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1197]),
	.d(FE_OFN322_n251459));
   oa22s01 U264135 (.o(n251464),
	.a(n251477),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1196]),
	.d(FE_OFN322_n251459));
   oa22s01 U264136 (.o(n251465),
	.a(n251477),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1195]),
	.d(FE_OFN322_n251459));
   oa22s01 U264137 (.o(n251466),
	.a(n251477),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1194]),
	.d(FE_OFN322_n251459));
   oa22s01 U264138 (.o(n251467),
	.a(n251477),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1193]),
	.d(FE_OFN322_n251459));
   oa22s01 U264139 (.o(n251468),
	.a(n251477),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1192]),
	.d(FE_OFN322_n251459));
   oa22s01 U264140 (.o(n251469),
	.a(n251477),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1191]),
	.d(FE_OFN322_n251459));
   oa22s01 U264141 (.o(n251471),
	.a(n251477),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1190]),
	.d(FE_OFN322_n251459));
   oa22s01 U264142 (.o(n251515),
	.a(n251548),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1151]),
	.d(FE_OFN204_n251530));
   oa22s01 U264143 (.o(n251516),
	.a(n251548),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1150]),
	.d(FE_OFN204_n251530));
   oa22s01 U264144 (.o(n251517),
	.a(n251548),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1149]),
	.d(FE_OFN204_n251530));
   oa22s01 U264145 (.o(n251518),
	.a(n251548),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1148]),
	.d(FE_OFN204_n251530));
   oa22s01 U264146 (.o(n251519),
	.a(n251548),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1147]),
	.d(FE_OFN204_n251530));
   oa22s01 U264147 (.o(n251520),
	.a(n251548),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1146]),
	.d(FE_OFN204_n251530));
   oa22s01 U264148 (.o(n251521),
	.a(n251548),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1145]),
	.d(FE_OFN204_n251530));
   oa22s01 U264149 (.o(n251523),
	.a(n251548),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1143]),
	.d(FE_OFN204_n251530));
   oa22s01 U264150 (.o(n251524),
	.a(n251548),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1142]),
	.d(FE_OFN204_n251530));
   oa22s01 U264151 (.o(n251525),
	.a(n251548),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1141]),
	.d(FE_OFN204_n251530));
   oa22s01 U264152 (.o(n251526),
	.a(n251548),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1140]),
	.d(FE_OFN204_n251530));
   oa22s01 U264153 (.o(n251527),
	.a(n251548),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1139]),
	.d(FE_OFN204_n251530));
   oa22s01 U264154 (.o(n251528),
	.a(n251548),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1138]),
	.d(FE_OFN204_n251530));
   oa22s01 U264155 (.o(n251529),
	.a(n251548),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1137]),
	.d(FE_OFN204_n251530));
   oa22s01 U264156 (.o(n251531),
	.a(n251548),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1136]),
	.d(FE_OFN204_n251530));
   oa22s01 U264157 (.o(n251532),
	.a(n251548),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1135]),
	.d(FE_OFN204_n251530));
   oa22s01 U264158 (.o(n251533),
	.a(n251548),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1134]),
	.d(FE_OFN204_n251530));
   oa22s01 U264159 (.o(n251534),
	.a(n251548),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1133]),
	.d(FE_OFN204_n251530));
   oa22s01 U264160 (.o(n251535),
	.a(n251548),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1132]),
	.d(FE_OFN204_n251530));
   oa22s01 U264161 (.o(n251536),
	.a(n251548),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1131]),
	.d(FE_OFN204_n251530));
   oa22s01 U264162 (.o(n251537),
	.a(n251548),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1130]),
	.d(FE_OFN204_n251530));
   oa22s01 U264163 (.o(n251539),
	.a(n251548),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1128]),
	.d(FE_OFN204_n251530));
   oa22s01 U264164 (.o(n251540),
	.a(n251548),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1127]),
	.d(FE_OFN204_n251530));
   oa22s01 U264165 (.o(n251542),
	.a(n251548),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1126]),
	.d(FE_OFN204_n251530));
   oa22s01 U264166 (.o(n251557),
	.a(n251583),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1112]),
	.d(FE_OFN324_n251565));
   oa22s01 U264167 (.o(n251559),
	.a(n251583),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1110]),
	.d(FE_OFN325_n251565));
   oa22s01 U264168 (.o(n251561),
	.a(n251583),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1108]),
	.d(FE_OFN325_n251565));
   oa22s01 U264169 (.o(n251563),
	.a(n251583),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1106]),
	.d(FE_OFN325_n251565));
   oa22s01 U264170 (.o(n251567),
	.a(n251583),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1103]),
	.d(FE_OFN324_n251565));
   oa22s01 U264171 (.o(n251568),
	.a(n251583),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1102]),
	.d(FE_OFN324_n251565));
   oa22s01 U264172 (.o(n251574),
	.a(n251583),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1096]),
	.d(FE_OFN325_n251565));
   oa22s01 U264173 (.o(n251575),
	.a(n251583),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1095]),
	.d(FE_OFN325_n251565));
   oa22s01 U264174 (.o(n251577),
	.a(n251583),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1094]),
	.d(FE_OFN324_n251565));
   oa22s01 U264175 (.o(n251585),
	.a(n251619),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1087]),
	.d(FE_OFN327_n251600));
   oa22s01 U264176 (.o(n251586),
	.a(n251619),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1086]),
	.d(FE_OFN327_n251600));
   oa22s01 U264177 (.o(n251587),
	.a(n251619),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1085]),
	.d(FE_OFN327_n251600));
   oa22s01 U264178 (.o(n251589),
	.a(n251619),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1083]),
	.d(FE_OFN327_n251600));
   oa22s01 U264179 (.o(n251590),
	.a(n251619),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1082]),
	.d(FE_OFN327_n251600));
   oa22s01 U264180 (.o(n251591),
	.a(n251619),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1081]),
	.d(FE_OFN327_n251600));
   oa22s01 U264181 (.o(n251592),
	.a(n251619),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1080]),
	.d(FE_OFN327_n251600));
   oa22s01 U264182 (.o(n251593),
	.a(n251619),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1079]),
	.d(FE_OFN327_n251600));
   oa22s01 U264183 (.o(n251594),
	.a(n251619),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1078]),
	.d(FE_OFN327_n251600));
   oa22s01 U264184 (.o(n251595),
	.a(n251619),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1077]),
	.d(FE_OFN327_n251600));
   oa22s01 U264185 (.o(n251596),
	.a(n251619),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1076]),
	.d(FE_OFN327_n251600));
   oa22s01 U264186 (.o(n251597),
	.a(n251619),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1075]),
	.d(FE_OFN327_n251600));
   oa22s01 U264187 (.o(n251598),
	.a(n251619),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1074]),
	.d(FE_OFN327_n251600));
   oa22s01 U264188 (.o(n251599),
	.a(n251619),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1073]),
	.d(FE_OFN327_n251600));
   oa22s01 U264189 (.o(n251601),
	.a(n251619),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1072]),
	.d(FE_OFN327_n251600));
   oa22s01 U264190 (.o(n251602),
	.a(n251619),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1071]),
	.d(FE_OFN327_n251600));
   oa22s01 U264191 (.o(n251603),
	.a(n251619),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1070]),
	.d(FE_OFN327_n251600));
   oa22s01 U264192 (.o(n251605),
	.a(n251619),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1068]),
	.d(FE_OFN327_n251600));
   oa22s01 U264193 (.o(n251606),
	.a(n251619),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1067]),
	.d(FE_OFN327_n251600));
   oa22s01 U264194 (.o(n251607),
	.a(n251619),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1066]),
	.d(FE_OFN327_n251600));
   oa22s01 U264195 (.o(n251609),
	.a(n251619),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1064]),
	.d(FE_OFN327_n251600));
   oa22s01 U264196 (.o(n251610),
	.a(n251619),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1063]),
	.d(FE_OFN327_n251600));
   oa22s01 U264197 (.o(n251612),
	.a(n251619),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1062]),
	.d(FE_OFN327_n251600));
   oa22s01 U264198 (.o(n251622),
	.a(n251655),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1055]),
	.d(FE_OFN329_n251637));
   oa22s01 U264199 (.o(n251624),
	.a(n251655),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1053]),
	.d(FE_OFN329_n251637));
   oa22s01 U264200 (.o(n251625),
	.a(n251655),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1052]),
	.d(FE_OFN329_n251637));
   oa22s01 U264201 (.o(n251626),
	.a(n251655),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1051]),
	.d(FE_OFN329_n251637));
   oa22s01 U264202 (.o(n251627),
	.a(n251655),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1050]),
	.d(FE_OFN329_n251637));
   oa22s01 U264203 (.o(n251628),
	.a(n251655),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1049]),
	.d(FE_OFN329_n251637));
   oa22s01 U264204 (.o(n251629),
	.a(n251655),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1048]),
	.d(FE_OFN329_n251637));
   oa22s01 U264205 (.o(n251630),
	.a(n251655),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1047]),
	.d(FE_OFN329_n251637));
   oa22s01 U264206 (.o(n251631),
	.a(n251655),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1046]),
	.d(FE_OFN329_n251637));
   oa22s01 U264207 (.o(n251632),
	.a(n251655),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1045]),
	.d(FE_OFN329_n251637));
   oa22s01 U264208 (.o(n251633),
	.a(n251655),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1044]),
	.d(FE_OFN329_n251637));
   oa22s01 U264209 (.o(n251634),
	.a(n251655),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1043]),
	.d(FE_OFN329_n251637));
   oa22s01 U264210 (.o(n251635),
	.a(n251655),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1042]),
	.d(FE_OFN329_n251637));
   oa22s01 U264211 (.o(n251636),
	.a(n251655),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1041]),
	.d(FE_OFN329_n251637));
   oa22s01 U264212 (.o(n251638),
	.a(n251655),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1040]),
	.d(FE_OFN329_n251637));
   oa22s01 U264213 (.o(n251640),
	.a(n251655),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1038]),
	.d(FE_OFN329_n251637));
   oa22s01 U264214 (.o(n251641),
	.a(n251655),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1037]),
	.d(FE_OFN329_n251637));
   oa22s01 U264215 (.o(n251642),
	.a(n251655),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1036]),
	.d(FE_OFN329_n251637));
   oa22s01 U264216 (.o(n251644),
	.a(n251655),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1034]),
	.d(FE_OFN329_n251637));
   oa22s01 U264217 (.o(n251645),
	.a(n251655),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1033]),
	.d(FE_OFN329_n251637));
   oa22s01 U264218 (.o(n251646),
	.a(n251655),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1032]),
	.d(FE_OFN329_n251637));
   oa22s01 U264219 (.o(n251647),
	.a(n251655),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1031]),
	.d(FE_OFN329_n251637));
   oa22s01 U264220 (.o(n251649),
	.a(n251655),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1030]),
	.d(FE_OFN329_n251637));
   oa22s01 U264221 (.o(n251657),
	.a(n251690),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[2047]),
	.d(FE_OFN331_n251675));
   oa22s01 U264222 (.o(n251658),
	.a(n251690),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[2046]),
	.d(FE_OFN331_n251675));
   oa22s01 U264223 (.o(n251659),
	.a(n251690),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[2045]),
	.d(FE_OFN331_n251675));
   oa22s01 U264224 (.o(n251661),
	.a(n251690),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[2043]),
	.d(FE_OFN331_n251675));
   oa22s01 U264225 (.o(n251662),
	.a(n251690),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[2042]),
	.d(FE_OFN331_n251675));
   oa22s01 U264226 (.o(n251663),
	.a(n251690),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[2041]),
	.d(FE_OFN331_n251675));
   oa22s01 U264227 (.o(n251664),
	.a(n251690),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[2040]),
	.d(FE_OFN331_n251675));
   oa22s01 U264228 (.o(n251665),
	.a(n251690),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[2039]),
	.d(FE_OFN331_n251675));
   oa22s01 U264229 (.o(n251666),
	.a(n251690),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[2038]),
	.d(FE_OFN331_n251675));
   oa22s01 U264230 (.o(n251667),
	.a(n251690),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[2037]),
	.d(FE_OFN331_n251675));
   oa22s01 U264231 (.o(n251668),
	.a(n251690),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[2036]),
	.d(FE_OFN331_n251675));
   oa22s01 U264232 (.o(n251669),
	.a(n251690),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[2035]),
	.d(FE_OFN331_n251675));
   oa22s01 U264233 (.o(n251670),
	.a(n251690),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[2034]),
	.d(FE_OFN331_n251675));
   oa22s01 U264234 (.o(n251672),
	.a(n251690),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[2032]),
	.d(FE_OFN331_n251675));
   oa22s01 U264235 (.o(n251673),
	.a(n251690),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[2031]),
	.d(FE_OFN331_n251675));
   oa22s01 U264236 (.o(n251674),
	.a(n251690),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[2030]),
	.d(FE_OFN331_n251675));
   oa22s01 U264237 (.o(n251676),
	.a(n251690),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[2029]),
	.d(FE_OFN331_n251675));
   oa22s01 U264238 (.o(n251677),
	.a(n251690),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[2028]),
	.d(FE_OFN331_n251675));
   oa22s01 U264239 (.o(n251678),
	.a(n251690),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[2027]),
	.d(FE_OFN331_n251675));
   oa22s01 U264240 (.o(n251679),
	.a(n251690),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[2026]),
	.d(FE_OFN331_n251675));
   oa22s01 U264241 (.o(n251680),
	.a(n251690),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[2025]),
	.d(FE_OFN331_n251675));
   oa22s01 U264242 (.o(n251681),
	.a(n251690),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[2024]),
	.d(FE_OFN331_n251675));
   oa22s01 U264243 (.o(n251682),
	.a(n251690),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[2023]),
	.d(FE_OFN331_n251675));
   oa22s01 U264244 (.o(n251684),
	.a(n251690),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[2022]),
	.d(FE_OFN331_n251675));
   oa22s01 U264245 (.o(n251692),
	.a(n251726),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[2015]),
	.d(n251710));
   oa22s01 U264246 (.o(n251694),
	.a(n251726),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[2013]),
	.d(FE_OFN430_n251710));
   oa22s01 U264247 (.o(n251695),
	.a(n251726),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[2012]),
	.d(FE_OFN430_n251710));
   oa22s01 U264248 (.o(n251696),
	.a(n251726),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[2011]),
	.d(FE_OFN430_n251710));
   oa22s01 U264249 (.o(n251697),
	.a(n251726),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[2010]),
	.d(FE_OFN430_n251710));
   oa22s01 U264250 (.o(n251698),
	.a(n251726),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[2009]),
	.d(n251710));
   oa22s01 U264251 (.o(n251699),
	.a(n251726),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[2008]),
	.d(FE_OFN430_n251710));
   oa22s01 U264252 (.o(n251700),
	.a(n251726),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[2007]),
	.d(FE_OFN430_n251710));
   oa22s01 U264253 (.o(n251701),
	.a(n251726),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[2006]),
	.d(FE_OFN430_n251710));
   oa22s01 U264254 (.o(n251702),
	.a(n251726),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[2005]),
	.d(FE_OFN430_n251710));
   oa22s01 U264255 (.o(n251703),
	.a(n251726),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[2004]),
	.d(FE_OFN430_n251710));
   oa22s01 U264256 (.o(n251705),
	.a(n251726),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[2002]),
	.d(FE_OFN430_n251710));
   oa22s01 U264257 (.o(n251706),
	.a(n251726),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[2001]),
	.d(FE_OFN430_n251710));
   oa22s01 U264258 (.o(n251707),
	.a(n251726),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[2000]),
	.d(FE_OFN430_n251710));
   oa22s01 U264259 (.o(n251708),
	.a(n251726),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1999]),
	.d(FE_OFN430_n251710));
   oa22s01 U264260 (.o(n251709),
	.a(n251726),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1998]),
	.d(FE_OFN430_n251710));
   oa22s01 U264261 (.o(n251711),
	.a(n251726),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1997]),
	.d(FE_OFN430_n251710));
   oa22s01 U264262 (.o(n251712),
	.a(n251726),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1996]),
	.d(FE_OFN430_n251710));
   oa22s01 U264263 (.o(n251713),
	.a(n251726),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1995]),
	.d(FE_OFN430_n251710));
   oa22s01 U264264 (.o(n251714),
	.a(n251726),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1994]),
	.d(n251710));
   oa22s01 U264265 (.o(n251715),
	.a(n251726),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1993]),
	.d(FE_OFN430_n251710));
   oa22s01 U264266 (.o(n251716),
	.a(n251726),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1992]),
	.d(n251710));
   oa22s01 U264267 (.o(n251717),
	.a(n251726),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1991]),
	.d(FE_OFN430_n251710));
   oa22s01 U264268 (.o(n251719),
	.a(n251726),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1990]),
	.d(FE_OFN430_n251710));
   oa22s01 U264269 (.o(n251728),
	.a(n251761),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1983]),
	.d(n251746));
   oa22s01 U264270 (.o(n251729),
	.a(n251761),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1982]),
	.d(FE_OFN333_n251746));
   oa22s01 U264271 (.o(n251730),
	.a(n251761),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1981]),
	.d(FE_OFN333_n251746));
   oa22s01 U264272 (.o(n251731),
	.a(n251761),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1980]),
	.d(FE_OFN333_n251746));
   oa22s01 U264273 (.o(n251732),
	.a(n251761),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1979]),
	.d(FE_OFN333_n251746));
   oa22s01 U264274 (.o(n251733),
	.a(n251761),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1978]),
	.d(FE_OFN333_n251746));
   oa22s01 U264275 (.o(n251734),
	.a(n251761),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1977]),
	.d(FE_OFN333_n251746));
   oa22s01 U264276 (.o(n251735),
	.a(n251761),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1976]),
	.d(FE_OFN333_n251746));
   oa22s01 U264277 (.o(n251736),
	.a(n251761),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1975]),
	.d(FE_OFN333_n251746));
   oa22s01 U264278 (.o(n251737),
	.a(n251761),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1974]),
	.d(FE_OFN333_n251746));
   oa22s01 U264279 (.o(n251739),
	.a(n251761),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1972]),
	.d(FE_OFN333_n251746));
   oa22s01 U264280 (.o(n251740),
	.a(n251761),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1971]),
	.d(FE_OFN333_n251746));
   oa22s01 U264281 (.o(n251741),
	.a(n251761),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1970]),
	.d(FE_OFN333_n251746));
   oa22s01 U264282 (.o(n251742),
	.a(n251761),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1969]),
	.d(FE_OFN333_n251746));
   oa22s01 U264283 (.o(n251743),
	.a(n251761),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1968]),
	.d(FE_OFN333_n251746));
   oa22s01 U264284 (.o(n251744),
	.a(n251761),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1967]),
	.d(FE_OFN333_n251746));
   oa22s01 U264285 (.o(n251745),
	.a(n251761),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1966]),
	.d(FE_OFN333_n251746));
   oa22s01 U264286 (.o(n251747),
	.a(n251761),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1965]),
	.d(FE_OFN333_n251746));
   oa22s01 U264287 (.o(n251748),
	.a(n251761),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1964]),
	.d(FE_OFN333_n251746));
   oa22s01 U264288 (.o(n251749),
	.a(n251761),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1963]),
	.d(FE_OFN333_n251746));
   oa22s01 U264289 (.o(n251750),
	.a(n251761),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1962]),
	.d(FE_OFN333_n251746));
   oa22s01 U264290 (.o(n251751),
	.a(n251761),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1961]),
	.d(FE_OFN333_n251746));
   oa22s01 U264291 (.o(n251752),
	.a(n251761),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1960]),
	.d(FE_OFN333_n251746));
   oa22s01 U264292 (.o(n251753),
	.a(n251761),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1959]),
	.d(FE_OFN333_n251746));
   oa22s01 U264293 (.o(n251763),
	.a(n251796),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1951]),
	.d(FE_OFN432_n251781));
   oa22s01 U264294 (.o(n251764),
	.a(n251796),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1950]),
	.d(FE_OFN432_n251781));
   oa22s01 U264295 (.o(n251765),
	.a(n251796),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1949]),
	.d(FE_OFN432_n251781));
   oa22s01 U264296 (.o(n251766),
	.a(n251796),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1948]),
	.d(FE_OFN432_n251781));
   oa22s01 U264297 (.o(n251767),
	.a(n251796),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1947]),
	.d(FE_OFN432_n251781));
   oa22s01 U264298 (.o(n251768),
	.a(n251796),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1946]),
	.d(FE_OFN432_n251781));
   oa22s01 U264299 (.o(n251769),
	.a(n251796),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1945]),
	.d(FE_OFN432_n251781));
   oa22s01 U264300 (.o(n251770),
	.a(n251796),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1944]),
	.d(FE_OFN432_n251781));
   oa22s01 U264301 (.o(n251772),
	.a(n251796),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1942]),
	.d(FE_OFN432_n251781));
   oa22s01 U264302 (.o(n251773),
	.a(n251796),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1941]),
	.d(FE_OFN432_n251781));
   oa22s01 U264303 (.o(n251774),
	.a(n251796),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1940]),
	.d(FE_OFN432_n251781));
   oa22s01 U264304 (.o(n251775),
	.a(n251796),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1939]),
	.d(FE_OFN432_n251781));
   oa22s01 U264305 (.o(n251776),
	.a(n251796),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1938]),
	.d(FE_OFN432_n251781));
   oa22s01 U264306 (.o(n251777),
	.a(n251796),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1937]),
	.d(FE_OFN432_n251781));
   oa22s01 U264307 (.o(n251778),
	.a(n251796),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1936]),
	.d(FE_OFN432_n251781));
   oa22s01 U264308 (.o(n251779),
	.a(n251796),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1935]),
	.d(FE_OFN432_n251781));
   oa22s01 U264309 (.o(n251780),
	.a(n251796),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1934]),
	.d(FE_OFN432_n251781));
   oa22s01 U264310 (.o(n251782),
	.a(n251796),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1933]),
	.d(FE_OFN432_n251781));
   oa22s01 U264311 (.o(n251783),
	.a(n251796),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1932]),
	.d(FE_OFN432_n251781));
   oa22s01 U264312 (.o(n251784),
	.a(n251796),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1931]),
	.d(FE_OFN432_n251781));
   oa22s01 U264313 (.o(n251785),
	.a(n251796),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1930]),
	.d(FE_OFN432_n251781));
   oa22s01 U264314 (.o(n251786),
	.a(n251796),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1929]),
	.d(FE_OFN432_n251781));
   oa22s01 U264315 (.o(n251788),
	.a(n251796),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1927]),
	.d(FE_OFN432_n251781));
   oa22s01 U264316 (.o(n251790),
	.a(n251796),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1926]),
	.d(FE_OFN432_n251781));
   oa22s01 U264317 (.o(n251798),
	.a(n251832),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1919]),
	.d(FE_OFN206_n251816));
   oa22s01 U264318 (.o(n251799),
	.a(n251832),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1918]),
	.d(FE_OFN206_n251816));
   oa22s01 U264319 (.o(n251800),
	.a(n251832),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1917]),
	.d(FE_OFN206_n251816));
   oa22s01 U264320 (.o(n251801),
	.a(n251832),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1916]),
	.d(FE_OFN206_n251816));
   oa22s01 U264321 (.o(n251802),
	.a(n251832),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1915]),
	.d(FE_OFN206_n251816));
   oa22s01 U264322 (.o(n251803),
	.a(n251832),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1914]),
	.d(FE_OFN206_n251816));
   oa22s01 U264323 (.o(n251805),
	.a(n251832),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1912]),
	.d(FE_OFN206_n251816));
   oa22s01 U264324 (.o(n251806),
	.a(n251832),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1911]),
	.d(FE_OFN206_n251816));
   oa22s01 U264325 (.o(n251807),
	.a(n251832),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1910]),
	.d(FE_OFN206_n251816));
   oa22s01 U264326 (.o(n251808),
	.a(n251832),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1909]),
	.d(FE_OFN206_n251816));
   oa22s01 U264327 (.o(n251809),
	.a(n251832),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1908]),
	.d(FE_OFN206_n251816));
   oa22s01 U264328 (.o(n251810),
	.a(n251832),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1907]),
	.d(FE_OFN206_n251816));
   oa22s01 U264329 (.o(n251811),
	.a(n251832),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1906]),
	.d(FE_OFN206_n251816));
   oa22s01 U264330 (.o(n251812),
	.a(n251832),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1905]),
	.d(FE_OFN206_n251816));
   oa22s01 U264331 (.o(n251813),
	.a(n251832),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1904]),
	.d(FE_OFN206_n251816));
   oa22s01 U264332 (.o(n251814),
	.a(n251832),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1903]),
	.d(FE_OFN206_n251816));
   oa22s01 U264333 (.o(n251815),
	.a(n251832),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1902]),
	.d(FE_OFN206_n251816));
   oa22s01 U264334 (.o(n251817),
	.a(n251832),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1901]),
	.d(FE_OFN206_n251816));
   oa22s01 U264335 (.o(n251818),
	.a(n251832),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1900]),
	.d(FE_OFN206_n251816));
   oa22s01 U264336 (.o(n251819),
	.a(n251832),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1899]),
	.d(FE_OFN206_n251816));
   oa22s01 U264337 (.o(n251821),
	.a(n251832),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1897]),
	.d(FE_OFN206_n251816));
   oa22s01 U264338 (.o(n251822),
	.a(n251832),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1896]),
	.d(FE_OFN206_n251816));
   oa22s01 U264339 (.o(n251823),
	.a(n251832),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1895]),
	.d(FE_OFN206_n251816));
   oa22s01 U264340 (.o(n251825),
	.a(n251832),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1894]),
	.d(FE_OFN206_n251816));
   oa22s01 U264341 (.o(n251834),
	.a(n251867),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1887]),
	.d(FE_OFN335_n251852));
   oa22s01 U264342 (.o(n251835),
	.a(n251867),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1886]),
	.d(FE_OFN335_n251852));
   oa22s01 U264343 (.o(n251836),
	.a(n251867),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1885]),
	.d(FE_OFN561_n251852));
   oa22s01 U264344 (.o(n251837),
	.a(n251867),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1884]),
	.d(FE_OFN560_n251852));
   oa22s01 U264345 (.o(n251839),
	.a(n251867),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1882]),
	.d(FE_OFN335_n251852));
   oa22s01 U264346 (.o(n251840),
	.a(n251867),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1881]),
	.d(FE_OFN335_n251852));
   oa22s01 U264347 (.o(n251841),
	.a(n251867),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1880]),
	.d(FE_OFN560_n251852));
   oa22s01 U264348 (.o(n251842),
	.a(n251867),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1879]),
	.d(FE_OFN561_n251852));
   oa22s01 U264349 (.o(n251843),
	.a(n251867),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1878]),
	.d(FE_OFN335_n251852));
   oa22s01 U264350 (.o(n251844),
	.a(n251867),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1877]),
	.d(FE_OFN335_n251852));
   oa22s01 U264351 (.o(n251845),
	.a(n251867),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1876]),
	.d(FE_OFN335_n251852));
   oa22s01 U264352 (.o(n251846),
	.a(n251867),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1875]),
	.d(FE_OFN335_n251852));
   oa22s01 U264353 (.o(n251847),
	.a(n251867),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1874]),
	.d(FE_OFN335_n251852));
   oa22s01 U264354 (.o(n251848),
	.a(n251867),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1873]),
	.d(FE_OFN335_n251852));
   oa22s01 U264355 (.o(n251849),
	.a(n251867),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1872]),
	.d(FE_OFN335_n251852));
   oa22s01 U264356 (.o(n251850),
	.a(n251867),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1871]),
	.d(FE_OFN561_n251852));
   oa22s01 U264357 (.o(n251851),
	.a(n251867),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1870]),
	.d(FE_OFN561_n251852));
   oa22s01 U264358 (.o(n251853),
	.a(n251867),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1869]),
	.d(FE_OFN561_n251852));
   oa22s01 U264359 (.o(n251855),
	.a(n251867),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1867]),
	.d(FE_OFN335_n251852));
   oa22s01 U264360 (.o(n251856),
	.a(n251867),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1866]),
	.d(FE_OFN561_n251852));
   oa22s01 U264361 (.o(n251857),
	.a(n251867),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1865]),
	.d(FE_OFN561_n251852));
   oa22s01 U264362 (.o(n251858),
	.a(n251867),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1864]),
	.d(FE_OFN335_n251852));
   oa22s01 U264363 (.o(n251859),
	.a(n251867),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1863]),
	.d(FE_OFN335_n251852));
   oa22s01 U264364 (.o(n251861),
	.a(n251867),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1862]),
	.d(FE_OFN561_n251852));
   oa22s01 U264365 (.o(n251869),
	.a(n251902),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1855]),
	.d(FE_OFN337_n251887));
   oa22s01 U264366 (.o(n251870),
	.a(n251902),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1854]),
	.d(FE_OFN337_n251887));
   oa22s01 U264367 (.o(n251872),
	.a(n251902),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1852]),
	.d(n251887));
   oa22s01 U264368 (.o(n251873),
	.a(n251902),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1851]),
	.d(FE_OFN337_n251887));
   oa22s01 U264369 (.o(n251874),
	.a(n251902),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1850]),
	.d(FE_OFN337_n251887));
   oa22s01 U264370 (.o(n251875),
	.a(n251902),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1849]),
	.d(FE_OFN337_n251887));
   oa22s01 U264371 (.o(n251876),
	.a(n251902),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1848]),
	.d(FE_OFN337_n251887));
   oa22s01 U264372 (.o(n251877),
	.a(n251902),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1847]),
	.d(FE_OFN337_n251887));
   oa22s01 U264373 (.o(n251878),
	.a(n251902),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1846]),
	.d(FE_OFN337_n251887));
   oa22s01 U264374 (.o(n251879),
	.a(n251902),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1845]),
	.d(FE_OFN337_n251887));
   oa22s01 U264375 (.o(n251880),
	.a(n251902),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1844]),
	.d(FE_OFN337_n251887));
   oa22s01 U264376 (.o(n251881),
	.a(n251902),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1843]),
	.d(FE_OFN337_n251887));
   oa22s01 U264377 (.o(n251882),
	.a(n251902),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1842]),
	.d(FE_OFN337_n251887));
   oa22s01 U264378 (.o(n251883),
	.a(n251902),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1841]),
	.d(FE_OFN337_n251887));
   oa22s01 U264379 (.o(n251884),
	.a(n251902),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1840]),
	.d(FE_OFN337_n251887));
   oa22s01 U264380 (.o(n251885),
	.a(n251902),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1839]),
	.d(n251887));
   oa22s01 U264381 (.o(n251888),
	.a(n251902),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1837]),
	.d(n251887));
   oa22s01 U264382 (.o(n251889),
	.a(n251902),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1836]),
	.d(FE_OFN337_n251887));
   oa22s01 U264383 (.o(n251890),
	.a(n251902),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1835]),
	.d(FE_OFN337_n251887));
   oa22s01 U264384 (.o(n251892),
	.a(n251902),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1833]),
	.d(n251887));
   oa22s01 U264385 (.o(n251893),
	.a(n251902),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1832]),
	.d(FE_OFN337_n251887));
   oa22s01 U264386 (.o(n251894),
	.a(n251902),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1831]),
	.d(n251887));
   oa22s01 U264387 (.o(n251896),
	.a(n251902),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1830]),
	.d(FE_OFN337_n251887));
   oa22s01 U264388 (.o(n251906),
	.a(n251939),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1822]),
	.d(FE_OFN339_n251923));
   oa22s01 U264389 (.o(n251907),
	.a(n251939),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1821]),
	.d(FE_OFN339_n251923));
   oa22s01 U264390 (.o(n251908),
	.a(n251939),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1820]),
	.d(FE_OFN339_n251923));
   oa22s01 U264391 (.o(n251909),
	.a(n251939),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1819]),
	.d(FE_OFN339_n251923));
   oa22s01 U264392 (.o(n251910),
	.a(n251939),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1818]),
	.d(FE_OFN339_n251923));
   oa22s01 U264393 (.o(n251911),
	.a(n251939),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1817]),
	.d(FE_OFN339_n251923));
   oa22s01 U264394 (.o(n251912),
	.a(n251939),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1816]),
	.d(FE_OFN339_n251923));
   oa22s01 U264395 (.o(n251913),
	.a(n251939),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1815]),
	.d(FE_OFN339_n251923));
   oa22s01 U264396 (.o(n251914),
	.a(n251939),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1814]),
	.d(FE_OFN339_n251923));
   oa22s01 U264397 (.o(n251915),
	.a(n251939),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1813]),
	.d(FE_OFN339_n251923));
   oa22s01 U264398 (.o(n251916),
	.a(n251939),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1812]),
	.d(FE_OFN339_n251923));
   oa22s01 U264399 (.o(n251917),
	.a(n251939),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1811]),
	.d(FE_OFN339_n251923));
   oa22s01 U264400 (.o(n251918),
	.a(n251939),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1810]),
	.d(FE_OFN339_n251923));
   oa22s01 U264401 (.o(n251919),
	.a(n251939),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1809]),
	.d(FE_OFN339_n251923));
   oa22s01 U264402 (.o(n251921),
	.a(n251939),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1807]),
	.d(FE_OFN339_n251923));
   oa22s01 U264403 (.o(n251922),
	.a(n251939),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1806]),
	.d(FE_OFN339_n251923));
   oa22s01 U264404 (.o(n251924),
	.a(n251939),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1805]),
	.d(FE_OFN339_n251923));
   oa22s01 U264405 (.o(n251926),
	.a(n251939),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1803]),
	.d(FE_OFN339_n251923));
   oa22s01 U264406 (.o(n251927),
	.a(n251939),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1802]),
	.d(FE_OFN339_n251923));
   oa22s01 U264407 (.o(n251928),
	.a(n251939),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1801]),
	.d(FE_OFN339_n251923));
   oa22s01 U264408 (.o(n251929),
	.a(n251939),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1800]),
	.d(FE_OFN339_n251923));
   oa22s01 U264409 (.o(n251930),
	.a(n251939),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1799]),
	.d(FE_OFN339_n251923));
   oa22s01 U264410 (.o(n251932),
	.a(n251939),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1798]),
	.d(FE_OFN339_n251923));
   oa22s01 U264411 (.o(n251942),
	.a(n251975),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1791]),
	.d(FE_OFN341_n251960));
   oa22s01 U264412 (.o(n251943),
	.a(n251975),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1790]),
	.d(FE_OFN341_n251960));
   oa22s01 U264413 (.o(n251945),
	.a(n251975),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1788]),
	.d(FE_OFN341_n251960));
   oa22s01 U264414 (.o(n251946),
	.a(n251975),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1787]),
	.d(FE_OFN341_n251960));
   oa22s01 U264415 (.o(n251947),
	.a(n251975),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1786]),
	.d(FE_OFN341_n251960));
   oa22s01 U264416 (.o(n251948),
	.a(n251975),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1785]),
	.d(FE_OFN341_n251960));
   oa22s01 U264417 (.o(n251949),
	.a(n251975),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1784]),
	.d(FE_OFN341_n251960));
   oa22s01 U264418 (.o(n251950),
	.a(n251975),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1783]),
	.d(FE_OFN341_n251960));
   oa22s01 U264419 (.o(n251951),
	.a(n251975),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1782]),
	.d(FE_OFN341_n251960));
   oa22s01 U264420 (.o(n251952),
	.a(n251975),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1781]),
	.d(FE_OFN341_n251960));
   oa22s01 U264421 (.o(n251953),
	.a(n251975),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1780]),
	.d(FE_OFN341_n251960));
   oa22s01 U264422 (.o(n251954),
	.a(n251975),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1779]),
	.d(FE_OFN341_n251960));
   oa22s01 U264423 (.o(n251956),
	.a(n251975),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1777]),
	.d(FE_OFN341_n251960));
   oa22s01 U264424 (.o(n251957),
	.a(n251975),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1776]),
	.d(FE_OFN341_n251960));
   oa22s01 U264425 (.o(n251958),
	.a(n251975),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1775]),
	.d(FE_OFN341_n251960));
   oa22s01 U264426 (.o(n251959),
	.a(n251975),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1774]),
	.d(FE_OFN341_n251960));
   oa22s01 U264427 (.o(n251961),
	.a(n251975),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1773]),
	.d(FE_OFN341_n251960));
   oa22s01 U264428 (.o(n251962),
	.a(n251975),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1772]),
	.d(FE_OFN341_n251960));
   oa22s01 U264429 (.o(n251963),
	.a(n251975),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1771]),
	.d(FE_OFN341_n251960));
   oa22s01 U264430 (.o(n251964),
	.a(n251975),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1770]),
	.d(FE_OFN341_n251960));
   oa22s01 U264431 (.o(n251965),
	.a(n251975),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1769]),
	.d(FE_OFN341_n251960));
   oa22s01 U264432 (.o(n251966),
	.a(n251975),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1768]),
	.d(FE_OFN341_n251960));
   oa22s01 U264433 (.o(n251967),
	.a(n251975),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1767]),
	.d(FE_OFN341_n251960));
   oa22s01 U264434 (.o(n251969),
	.a(n251975),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1766]),
	.d(FE_OFN341_n251960));
   oa22s01 U264435 (.o(n251979),
	.a(n252011),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1758]),
	.d(FE_OFN434_n251996));
   oa22s01 U264436 (.o(n251980),
	.a(n252011),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1757]),
	.d(FE_OFN434_n251996));
   oa22s01 U264437 (.o(n251981),
	.a(n252011),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1756]),
	.d(FE_OFN434_n251996));
   oa22s01 U264438 (.o(n251982),
	.a(n252011),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1755]),
	.d(FE_OFN434_n251996));
   oa22s01 U264439 (.o(n251983),
	.a(n252011),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1754]),
	.d(FE_OFN434_n251996));
   oa22s01 U264440 (.o(n251984),
	.a(n252011),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1753]),
	.d(FE_OFN434_n251996));
   oa22s01 U264441 (.o(n251985),
	.a(n252011),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1752]),
	.d(FE_OFN434_n251996));
   oa22s01 U264442 (.o(n251986),
	.a(n252011),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1751]),
	.d(FE_OFN434_n251996));
   oa22s01 U264443 (.o(n251987),
	.a(n252011),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1750]),
	.d(FE_OFN434_n251996));
   oa22s01 U264444 (.o(n251988),
	.a(n252011),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1749]),
	.d(FE_OFN434_n251996));
   oa22s01 U264445 (.o(n251990),
	.a(n252011),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1747]),
	.d(FE_OFN434_n251996));
   oa22s01 U264446 (.o(n251991),
	.a(n252011),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1746]),
	.d(FE_OFN434_n251996));
   oa22s01 U264447 (.o(n251992),
	.a(n252011),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1745]),
	.d(FE_OFN434_n251996));
   oa22s01 U264448 (.o(n251993),
	.a(n252011),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1744]),
	.d(FE_OFN434_n251996));
   oa22s01 U264449 (.o(n251994),
	.a(n252011),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1743]),
	.d(FE_OFN434_n251996));
   oa22s01 U264450 (.o(n251995),
	.a(n252011),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1742]),
	.d(FE_OFN434_n251996));
   oa22s01 U264451 (.o(n251997),
	.a(n252011),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1741]),
	.d(FE_OFN434_n251996));
   oa22s01 U264452 (.o(n251998),
	.a(n252011),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1740]),
	.d(FE_OFN434_n251996));
   oa22s01 U264453 (.o(n251999),
	.a(n252011),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1739]),
	.d(FE_OFN434_n251996));
   oa22s01 U264454 (.o(n252000),
	.a(n252011),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1738]),
	.d(FE_OFN434_n251996));
   oa22s01 U264455 (.o(n252001),
	.a(n252011),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1737]),
	.d(FE_OFN434_n251996));
   oa22s01 U264456 (.o(n252002),
	.a(n252011),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1736]),
	.d(FE_OFN434_n251996));
   oa22s01 U264457 (.o(n252003),
	.a(n252011),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1735]),
	.d(FE_OFN434_n251996));
   oa22s01 U264458 (.o(n252005),
	.a(n252011),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1734]),
	.d(FE_OFN434_n251996));
   oa22s01 U264459 (.o(n252014),
	.a(n252048),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1727]),
	.d(FE_OFN343_n252032));
   oa22s01 U264460 (.o(n252015),
	.a(n252048),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1726]),
	.d(FE_OFN343_n252032));
   oa22s01 U264461 (.o(n252016),
	.a(n252048),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1725]),
	.d(FE_OFN343_n252032));
   oa22s01 U264462 (.o(n252017),
	.a(n252048),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1724]),
	.d(FE_OFN343_n252032));
   oa22s01 U264463 (.o(n252018),
	.a(n252048),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1723]),
	.d(FE_OFN343_n252032));
   oa22s01 U264464 (.o(n252019),
	.a(n252048),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1722]),
	.d(FE_OFN343_n252032));
   oa22s01 U264465 (.o(n252021),
	.a(n252048),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1720]),
	.d(FE_OFN343_n252032));
   oa22s01 U264466 (.o(n252025),
	.a(n252048),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1716]),
	.d(FE_OFN343_n252032));
   oa22s01 U264467 (.o(n252027),
	.a(n252048),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1714]),
	.d(FE_OFN343_n252032));
   oa22s01 U264468 (.o(n252030),
	.a(n252048),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1711]),
	.d(FE_OFN343_n252032));
   oa22s01 U264469 (.o(n252031),
	.a(n252048),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1710]),
	.d(FE_OFN343_n252032));
   oa22s01 U264470 (.o(n252034),
	.a(n252048),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1708]),
	.d(FE_OFN343_n252032));
   oa22s01 U264471 (.o(n252035),
	.a(n252048),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1707]),
	.d(FE_OFN343_n252032));
   oa22s01 U264472 (.o(n252036),
	.a(n252048),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1706]),
	.d(FE_OFN343_n252032));
   oa22s01 U264473 (.o(n252037),
	.a(n252048),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1705]),
	.d(FE_OFN343_n252032));
   oa22s01 U264474 (.o(n252038),
	.a(n252048),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1704]),
	.d(FE_OFN343_n252032));
   oa22s01 U264475 (.o(n252041),
	.a(n252048),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1702]),
	.d(FE_OFN343_n252032));
   oa22s01 U264476 (.o(n252087),
	.a(n252120),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1663]),
	.d(FE_OFN208_n252105));
   oa22s01 U264477 (.o(n252088),
	.a(n252120),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1662]),
	.d(FE_OFN208_n252105));
   oa22s01 U264478 (.o(n252089),
	.a(n252120),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1661]),
	.d(FE_OFN208_n252105));
   oa22s01 U264479 (.o(n252090),
	.a(n252120),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1660]),
	.d(FE_OFN208_n252105));
   oa22s01 U264480 (.o(n252091),
	.a(n252120),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1659]),
	.d(FE_OFN208_n252105));
   oa22s01 U264481 (.o(n252093),
	.a(n252120),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1657]),
	.d(FE_OFN208_n252105));
   oa22s01 U264482 (.o(n252094),
	.a(n252120),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1656]),
	.d(FE_OFN208_n252105));
   oa22s01 U264483 (.o(n252095),
	.a(n252120),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1655]),
	.d(FE_OFN208_n252105));
   oa22s01 U264484 (.o(n252096),
	.a(n252120),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1654]),
	.d(FE_OFN208_n252105));
   oa22s01 U264485 (.o(n252097),
	.a(n252120),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1653]),
	.d(FE_OFN208_n252105));
   oa22s01 U264486 (.o(n252098),
	.a(n252120),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1652]),
	.d(FE_OFN208_n252105));
   oa22s01 U264487 (.o(n252099),
	.a(n252120),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1651]),
	.d(FE_OFN208_n252105));
   oa22s01 U264488 (.o(n252100),
	.a(n252120),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1650]),
	.d(FE_OFN208_n252105));
   oa22s01 U264489 (.o(n252101),
	.a(n252120),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1649]),
	.d(FE_OFN208_n252105));
   oa22s01 U264490 (.o(n252102),
	.a(n252120),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1648]),
	.d(FE_OFN208_n252105));
   oa22s01 U264491 (.o(n252103),
	.a(n252120),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1647]),
	.d(FE_OFN208_n252105));
   oa22s01 U264492 (.o(n252104),
	.a(n252120),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1646]),
	.d(FE_OFN208_n252105));
   oa22s01 U264493 (.o(n252106),
	.a(n252120),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1645]),
	.d(FE_OFN208_n252105));
   oa22s01 U264494 (.o(n252107),
	.a(n252120),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1644]),
	.d(FE_OFN208_n252105));
   oa22s01 U264495 (.o(n252109),
	.a(n252120),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1642]),
	.d(FE_OFN208_n252105));
   oa22s01 U264496 (.o(n252110),
	.a(n252120),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1641]),
	.d(FE_OFN208_n252105));
   oa22s01 U264497 (.o(n252111),
	.a(n252120),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1640]),
	.d(FE_OFN208_n252105));
   oa22s01 U264498 (.o(n252112),
	.a(n252120),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1639]),
	.d(FE_OFN208_n252105));
   oa22s01 U264499 (.o(n252114),
	.a(n252120),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1638]),
	.d(FE_OFN208_n252105));
   oa22s01 U264500 (.o(n252123),
	.a(n252157),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1631]),
	.d(FE_OFN346_n252141));
   oa22s01 U264501 (.o(n252124),
	.a(n252157),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1630]),
	.d(FE_OFN346_n252141));
   oa22s01 U264502 (.o(n252125),
	.a(n252157),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1629]),
	.d(FE_OFN345_n252141));
   oa22s01 U264503 (.o(n252127),
	.a(n252157),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1627]),
	.d(FE_OFN345_n252141));
   oa22s01 U264504 (.o(n252128),
	.a(n252157),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1626]),
	.d(FE_OFN346_n252141));
   oa22s01 U264505 (.o(n252129),
	.a(n252157),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1625]),
	.d(FE_OFN346_n252141));
   oa22s01 U264506 (.o(n252130),
	.a(n252157),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1624]),
	.d(FE_OFN345_n252141));
   oa22s01 U264507 (.o(n252131),
	.a(n252157),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1623]),
	.d(FE_OFN345_n252141));
   oa22s01 U264508 (.o(n252132),
	.a(n252157),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1622]),
	.d(FE_OFN346_n252141));
   oa22s01 U264509 (.o(n252133),
	.a(n252157),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1621]),
	.d(FE_OFN346_n252141));
   oa22s01 U264510 (.o(n252134),
	.a(n252157),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1620]),
	.d(FE_OFN346_n252141));
   oa22s01 U264511 (.o(n252135),
	.a(n252157),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1619]),
	.d(FE_OFN346_n252141));
   oa22s01 U264512 (.o(n252136),
	.a(n252157),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1618]),
	.d(FE_OFN346_n252141));
   oa22s01 U264513 (.o(n252137),
	.a(n252157),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1617]),
	.d(FE_OFN346_n252141));
   oa22s01 U264514 (.o(n252138),
	.a(n252157),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1616]),
	.d(FE_OFN346_n252141));
   oa22s01 U264515 (.o(n252139),
	.a(n252157),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1615]),
	.d(FE_OFN345_n252141));
   oa22s01 U264516 (.o(n252140),
	.a(n252157),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1614]),
	.d(FE_OFN345_n252141));
   oa22s01 U264517 (.o(n252143),
	.a(n252157),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1612]),
	.d(FE_OFN346_n252141));
   oa22s01 U264518 (.o(n252144),
	.a(n252157),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1611]),
	.d(FE_OFN346_n252141));
   oa22s01 U264519 (.o(n252145),
	.a(n252157),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1610]),
	.d(FE_OFN345_n252141));
   oa22s01 U264520 (.o(n252147),
	.a(n252157),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1608]),
	.d(FE_OFN346_n252141));
   oa22s01 U264521 (.o(n252148),
	.a(n252157),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1607]),
	.d(FE_OFN346_n252141));
   oa22s01 U264522 (.o(n252150),
	.a(n252157),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1606]),
	.d(FE_OFN345_n252141));
   oa22s01 U264523 (.o(n252160),
	.a(n252193),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1599]),
	.d(FE_OFN348_n252178));
   oa22s01 U264524 (.o(n252162),
	.a(n252193),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1597]),
	.d(FE_OFN348_n252178));
   oa22s01 U264525 (.o(n252163),
	.a(n252193),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1596]),
	.d(FE_OFN348_n252178));
   oa22s01 U264526 (.o(n252164),
	.a(n252193),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1595]),
	.d(FE_OFN348_n252178));
   oa22s01 U264527 (.o(n252165),
	.a(n252193),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1594]),
	.d(FE_OFN348_n252178));
   oa22s01 U264528 (.o(n252166),
	.a(n252193),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1593]),
	.d(FE_OFN348_n252178));
   oa22s01 U264529 (.o(n252167),
	.a(n252193),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1592]),
	.d(FE_OFN348_n252178));
   oa22s01 U264530 (.o(n252168),
	.a(n252193),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1591]),
	.d(FE_OFN348_n252178));
   oa22s01 U264531 (.o(n252169),
	.a(n252193),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1590]),
	.d(FE_OFN348_n252178));
   oa22s01 U264532 (.o(n252170),
	.a(n252193),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1589]),
	.d(FE_OFN348_n252178));
   oa22s01 U264533 (.o(n252171),
	.a(n252193),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1588]),
	.d(FE_OFN348_n252178));
   oa22s01 U264534 (.o(n252172),
	.a(n252193),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1587]),
	.d(FE_OFN348_n252178));
   oa22s01 U264535 (.o(n252173),
	.a(n252193),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1586]),
	.d(FE_OFN348_n252178));
   oa22s01 U264536 (.o(n252174),
	.a(n252193),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1585]),
	.d(FE_OFN348_n252178));
   oa22s01 U264537 (.o(n252175),
	.a(n252193),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1584]),
	.d(FE_OFN348_n252178));
   oa22s01 U264538 (.o(n252177),
	.a(n252193),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1582]),
	.d(FE_OFN348_n252178));
   oa22s01 U264539 (.o(n252179),
	.a(n252193),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1581]),
	.d(FE_OFN348_n252178));
   oa22s01 U264540 (.o(n252180),
	.a(n252193),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1580]),
	.d(FE_OFN348_n252178));
   oa22s01 U264541 (.o(n252182),
	.a(n252193),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1578]),
	.d(FE_OFN348_n252178));
   oa22s01 U264542 (.o(n252183),
	.a(n252193),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1577]),
	.d(FE_OFN348_n252178));
   oa22s01 U264543 (.o(n252184),
	.a(n252193),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1576]),
	.d(FE_OFN348_n252178));
   oa22s01 U264544 (.o(n252185),
	.a(n252193),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1575]),
	.d(FE_OFN348_n252178));
   oa22s01 U264545 (.o(n252187),
	.a(n252193),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1574]),
	.d(FE_OFN348_n252178));
   oa22s01 U264546 (.o(n252197),
	.a(n252230),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1567]),
	.d(FE_OFN350_n252215));
   oa22s01 U264547 (.o(n252198),
	.a(n252230),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1566]),
	.d(FE_OFN350_n252215));
   oa22s01 U264548 (.o(n252199),
	.a(n252230),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1565]),
	.d(FE_OFN350_n252215));
   oa22s01 U264549 (.o(n252201),
	.a(n252230),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1563]),
	.d(FE_OFN350_n252215));
   oa22s01 U264550 (.o(n252202),
	.a(n252230),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1562]),
	.d(FE_OFN350_n252215));
   oa22s01 U264551 (.o(n252203),
	.a(n252230),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1561]),
	.d(FE_OFN350_n252215));
   oa22s01 U264552 (.o(n252204),
	.a(n252230),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1560]),
	.d(FE_OFN350_n252215));
   oa22s01 U264553 (.o(n252205),
	.a(n252230),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1559]),
	.d(FE_OFN350_n252215));
   oa22s01 U264554 (.o(n252206),
	.a(n252230),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1558]),
	.d(FE_OFN350_n252215));
   oa22s01 U264555 (.o(n252207),
	.a(n252230),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1557]),
	.d(FE_OFN350_n252215));
   oa22s01 U264556 (.o(n252208),
	.a(n252230),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1556]),
	.d(FE_OFN350_n252215));
   oa22s01 U264557 (.o(n252209),
	.a(n252230),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1555]),
	.d(FE_OFN350_n252215));
   oa22s01 U264558 (.o(n252210),
	.a(n252230),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1554]),
	.d(FE_OFN350_n252215));
   oa22s01 U264559 (.o(n252212),
	.a(n252230),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1552]),
	.d(FE_OFN350_n252215));
   oa22s01 U264560 (.o(n252213),
	.a(n252230),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1551]),
	.d(FE_OFN350_n252215));
   oa22s01 U264561 (.o(n252214),
	.a(n252230),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1550]),
	.d(FE_OFN350_n252215));
   oa22s01 U264562 (.o(n252216),
	.a(n252230),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1549]),
	.d(FE_OFN350_n252215));
   oa22s01 U264563 (.o(n252217),
	.a(n252230),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1548]),
	.d(FE_OFN350_n252215));
   oa22s01 U264564 (.o(n252218),
	.a(n252230),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1547]),
	.d(FE_OFN350_n252215));
   oa22s01 U264565 (.o(n252219),
	.a(n252230),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1546]),
	.d(FE_OFN350_n252215));
   oa22s01 U264566 (.o(n252220),
	.a(n252230),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1545]),
	.d(FE_OFN350_n252215));
   oa22s01 U264567 (.o(n252221),
	.a(n252230),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1544]),
	.d(FE_OFN350_n252215));
   oa22s01 U264568 (.o(n252222),
	.a(n252230),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1543]),
	.d(FE_OFN350_n252215));
   oa22s01 U264569 (.o(n252224),
	.a(n252230),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1542]),
	.d(FE_OFN350_n252215));
   in01f01 U264571 (.o(n249032),
	.a(n249052));
   oa12f01 U264572 (.o(n244991),
	.a(n248998),
	.b(n249077),
	.c(FE_OFN491_regtop_g_a_r_3_));
   ao12f01 U264573 (.o(n248998),
	.a(n249211),
	.b(n248997),
	.c(n249073));
   no02f01 U264574 (.o(n248995),
	.a(n248994),
	.b(n248992));
   oa12f01 U264575 (.o(n244992),
	.a(n248988),
	.b(n249077),
	.c(FE_OFN548_regtop_g_a_r_2_));
   na02f01 U264576 (.o(n244995),
	.a(n249188),
	.b(n249187));
   na02f01 U264577 (.o(n244996),
	.a(n249182),
	.b(n249181));
   no02f01 U264578 (.o(n249182),
	.a(n249179),
	.b(n249178));
   na02f01 U264579 (.o(n244997),
	.a(n249175),
	.b(n249174));
   no02f02 U264580 (.o(n249175),
	.a(n249173),
	.b(n249172));
   na02f01 U264581 (.o(n244998),
	.a(n249169),
	.b(n249168));
   na02f01 U264582 (.o(n244999),
	.a(n249163),
	.b(n249162));
   no02f02 U264583 (.o(n249163),
	.a(n249161),
	.b(n249160));
   na02f01 U264584 (.o(n245000),
	.a(n249158),
	.b(n249157));
   no02f02 U264585 (.o(n249158),
	.a(n249156),
	.b(n249155));
   na02f01 U264586 (.o(n245001),
	.a(n249153),
	.b(n249152));
   no02f02 U264587 (.o(n249153),
	.a(n249151),
	.b(n249150));
   na02f01 U264588 (.o(n245002),
	.a(n249219),
	.b(n249218));
   ao12f01 U264589 (.o(n249219),
	.a(n249217),
	.b(n249252),
	.c(regtop_g_usrd_r[8]));
   oa12f01 U264590 (.o(n249217),
	.a(n249216),
	.b(n249250),
	.c(n252810));
   na02f04 U264591 (.o(n245003),
	.a(n249148),
	.b(n249147));
   ao12f01 U264592 (.o(n249148),
	.a(n249146),
	.b(n249252),
	.c(regtop_g_usrd_r[9]));
   oa12f02 U264593 (.o(n249146),
	.a(n249145),
	.b(n249250),
	.c(n252782));
   na02f02 U264594 (.o(n245004),
	.a(n249233),
	.b(n249232));
   ao12f01 U264595 (.o(n249233),
	.a(n249231),
	.b(n249252),
	.c(regtop_g_usrd_r[10]));
   oa12f01 U264596 (.o(n249231),
	.a(n249230),
	.b(n249250),
	.c(n252786));
   na02f01 U264597 (.o(n245005),
	.a(n249240),
	.b(n249239));
   ao12f01 U264598 (.o(n249240),
	.a(n249238),
	.b(n249252),
	.c(regtop_g_usrd_r[11]));
   oa12f01 U264599 (.o(n249238),
	.a(n249237),
	.b(n249250),
	.c(n252790));
   na02s02 U264600 (.o(n245006),
	.a(n249254),
	.b(n249253));
   ao12f01 U264601 (.o(n249254),
	.a(n249251),
	.b(n249252),
	.c(regtop_g_usrd_r[12]));
   oa12f01 U264602 (.o(n249251),
	.a(n249249),
	.b(n249250),
	.c(n252794));
   na02f01 U264603 (.o(n245007),
	.a(n249202),
	.b(n249201));
   oa12f01 U264604 (.o(n249200),
	.a(n249199),
	.b(n249250),
	.c(n252798));
   ao12f01 U264605 (.o(n249226),
	.a(n249224),
	.b(n249252),
	.c(regtop_g_usrd_r[14]));
   oa12f01 U264606 (.o(n249224),
	.a(n249223),
	.b(n249250),
	.c(n252802));
   na02f02 U264607 (.o(n245009),
	.a(n249209),
	.b(n249208));
   ao12f01 U264608 (.o(n249209),
	.a(n249207),
	.b(n249252),
	.c(regtop_g_usrd_r[15]));
   oa12f01 U264609 (.o(n249207),
	.a(n249206),
	.b(n249250),
	.c(n252806));
   ao12f01 U264610 (.o(n249134),
	.a(n249131),
	.b(regtop_g_paramdata_r[19]),
	.c(n249132));
   na02f01 U264611 (.o(n245013),
	.a(n249094),
	.b(n249093));
   ao12f01 U264612 (.o(n249094),
	.a(n249092),
	.b(regtop_g_paramdata_r[20]),
	.c(n249132));
   na02f01 U264613 (.o(n245014),
	.a(n249105),
	.b(n249104));
   ao12f01 U264614 (.o(n249105),
	.a(n249103),
	.b(regtop_g_paramdata_r[21]),
	.c(n249132));
   na02f01 U264615 (.o(n245015),
	.a(n249125),
	.b(n249124));
   ao12f01 U264616 (.o(n249125),
	.a(n249123),
	.b(regtop_g_paramdata_r[22]),
	.c(n249132));
   na03f01 U264617 (.o(n245016),
	.a(n249085),
	.b(n249084),
	.c(n249083));
   ao22s01 U264618 (.o(n249085),
	.a(n249127),
	.b(regtop_g_atscd_r[22]),
	.c(n249128),
	.d(regtop_g_usrd_r[22]));
   na02f02 U264619 (.o(n249084),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[22]));
   na03f01 U264620 (.o(n245017),
	.a(n249088),
	.b(n249087),
	.c(n249086));
   ao22s01 U264621 (.o(n249088),
	.a(n249127),
	.b(regtop_g_atscd_r[23]),
	.c(n249128),
	.d(regtop_g_usrd_r[23]));
   na02f01 U264622 (.o(n249087),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[23]));
   na03f02 U264623 (.o(n245018),
	.a(n248964),
	.b(n248963),
	.c(n248962));
   na02f01 U264624 (.o(n248962),
	.a(regtop_g_paramdata_r[17]),
	.b(n248980));
   na02f01 U264625 (.o(n248963),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[24]));
   na03f03 U264626 (.o(n245019),
	.a(n248983),
	.b(n248982),
	.c(n248981));
   na02f01 U264627 (.o(n248981),
	.a(regtop_g_paramdata_r[18]),
	.b(n248980));
   na02f01 U264628 (.o(n248982),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[25]));
   na03f04 U264629 (.o(n245020),
	.a(n248976),
	.b(n248975),
	.c(n248974));
   na02f01 U264630 (.o(n248974),
	.a(regtop_g_paramdata_r[19]),
	.b(n248980));
   na02f01 U264631 (.o(n248975),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[26]));
   na03f03 U264632 (.o(n245021),
	.a(n248958),
	.b(n248957),
	.c(n248956));
   na03f03 U264633 (.o(n245022),
	.a(n248967),
	.b(n248966),
	.c(n248965));
   na02f01 U264634 (.o(n248965),
	.a(regtop_g_paramdata_r[21]),
	.b(n248980));
   na03f06 U264635 (.o(n245023),
	.a(n248970),
	.b(n248969),
	.c(n248968));
   na02f01 U264636 (.o(n248968),
	.a(regtop_g_paramdata_r[22]),
	.b(n248980));
   na03f01 U264637 (.o(n245024),
	.a(n248973),
	.b(n248972),
	.c(n248971));
   na02f01 U264638 (.o(n248971),
	.a(regtop_g_paramdata_r[23]),
	.b(n248980));
   na02f01 U264639 (.o(n248960),
	.a(FE_OFN502_n246205),
	.b(regtop_g_wd_r[31]));
   na02f01 U264640 (.o(n245010),
	.a(n249120),
	.b(n249119));
   ao12f01 U264641 (.o(n249120),
	.a(n249118),
	.b(regtop_g_paramdata_r[17]),
	.c(n249132));
   na02f01 U264642 (.o(n245011),
	.a(n249100),
	.b(n249099));
   ao12f01 U264643 (.o(n249100),
	.a(n249098),
	.b(regtop_g_paramdata_r[18]),
	.c(n249132));
   na02f01 U264644 (.o(n186680),
	.a(n252262),
	.b(n252261));
   ao22f01 U264645 (.o(n252262),
	.a(n252269),
	.b(regtop_g_wd_r[17]),
	.c(regtop_g_icfb_r),
	.d(n252259));
   na04f03 U264646 (.o(n252259),
	.a(n252258),
	.b(n252257),
	.c(n252298),
	.d(n252296));
   ao22s01 U264647 (.o(n247601),
	.a(regtop_g_wd_r[0]),
	.b(n247603),
	.c(regtop_g_adb_cpu_r[0]),
	.d(n247602));
   ao22s01 U264648 (.o(n247600),
	.a(regtop_g_wd_r[1]),
	.b(n247603),
	.c(regtop_g_adb_cpu_r[1]),
	.d(n247602));
   ao22s01 U264649 (.o(n247604),
	.a(regtop_g_wd_r[2]),
	.b(n247603),
	.c(regtop_g_adb_cpu_r[2]),
	.d(n247602));
   ao22s01 U264650 (.o(n247598),
	.a(regtop_g_wd_r[3]),
	.b(n247603),
	.c(regtop_g_adb_cpu_r[3]),
	.d(n247602));
   ao22s01 U264651 (.o(n247597),
	.a(regtop_g_wd_r[4]),
	.b(n247603),
	.c(regtop_g_adb_cpu_r[4]),
	.d(n247602));
   ao22s01 U264652 (.o(n247599),
	.a(regtop_g_wd_r[5]),
	.b(n247603),
	.c(regtop_g_adb_cpu_r[5]),
	.d(n247602));
   ao22s01 U264653 (.o(n247596),
	.a(regtop_g_wd_r[6]),
	.b(n247603),
	.c(regtop_g_adb_cpu_r[6]),
	.d(n247602));
   ao22s01 U264654 (.o(n252287),
	.a(n252377),
	.b(regtop_g_tmg_ferr_hit_r),
	.c(n252300),
	.d(regtop_g_fbst_r[9]));
   ao22s01 U264655 (.o(n252303),
	.a(n252302),
	.b(n252301),
	.c(regtop_g_fbst_r[6]),
	.d(n252300));
   ao22s01 U264656 (.o(n246595),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[13]),
	.c(FE_OFN486_n245940),
	.d(regtop_g_hsv_r[0]));
   ao22s01 U264657 (.o(n246590),
	.a(regtop_g_paramdata_r[24]),
	.b(FE_OFN366_n246266),
	.c(FE_OFN486_n245940),
	.d(regtop_g_hsv_r[11]));
   ao22s01 U264658 (.o(n246589),
	.a(regtop_g_paramdata_r[23]),
	.b(FE_OFN366_n246266),
	.c(FE_OFN486_n245940),
	.d(regtop_g_hsv_r[10]));
   ao22s01 U264659 (.o(n246594),
	.a(regtop_g_paramdata_r[22]),
	.b(FE_OFN366_n246266),
	.c(FE_OFN486_n245940),
	.d(regtop_g_hsv_r[9]));
   ao22s01 U264660 (.o(n246588),
	.a(regtop_g_paramdata_r[21]),
	.b(FE_OFN366_n246266),
	.c(FE_OFN486_n245940),
	.d(regtop_g_hsv_r[8]));
   ao22s01 U264661 (.o(n246592),
	.a(regtop_g_paramdata_r[20]),
	.b(FE_OFN366_n246266),
	.c(FE_OFN486_n245940),
	.d(regtop_g_hsv_r[7]));
   ao22s01 U264662 (.o(n246606),
	.a(regtop_g_paramdata_r[19]),
	.b(FE_OFN366_n246266),
	.c(FE_OFN486_n245940),
	.d(regtop_g_hsv_r[6]));
   ao22s01 U264663 (.o(n246603),
	.a(regtop_g_paramdata_r[18]),
	.b(FE_OFN366_n246266),
	.c(FE_OFN486_n245940),
	.d(regtop_g_hsv_r[5]));
   ao22s01 U264664 (.o(n246601),
	.a(regtop_g_paramdata_r[16]),
	.b(FE_OFN366_n246266),
	.c(FE_OFN486_n245940),
	.d(regtop_g_hsv_r[3]));
   ao22s01 U264665 (.o(n246600),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[15]),
	.c(FE_OFN486_n245940),
	.d(regtop_g_hsv_r[2]));
   ao22s01 U264666 (.o(n246598),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[14]),
	.c(FE_OFN486_n245940),
	.d(regtop_g_hsv_r[1]));
   ao22s01 U264667 (.o(n246591),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[5]),
	.c(FE_OFN486_n245940),
	.d(regtop_g_vsv_r[4]));
   ao22s01 U264668 (.o(n246596),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[6]),
	.c(FE_OFN486_n245940),
	.d(regtop_g_vsv_r[5]));
   ao22s01 U264669 (.o(n246586),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[7]),
	.c(FE_OFN486_n245940),
	.d(regtop_g_vsv_r[6]));
   ao22s01 U264670 (.o(n246593),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[8]),
	.c(n245940),
	.d(regtop_g_vsv_r[7]));
   ao22s01 U264671 (.o(n246604),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[9]),
	.c(FE_OFN485_n245940),
	.d(regtop_g_vsv_r[8]));
   ao22s01 U264672 (.o(n246597),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[11]),
	.c(n245940),
	.d(regtop_g_vsv_r[10]));
   ao22s01 U264673 (.o(n246599),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[12]),
	.c(n245940),
	.d(regtop_g_vsv_r[11]));
   ao22f01 U264674 (.o(n246926),
	.a(n246925),
	.b(n246924),
	.c(regtop_g_udb0_r[6]),
	.d(n246923));
   in01s01 U264675 (.o(n246923),
	.a(n246925));
   in01s01 U264676 (.o(n211949),
	.a(n247043));
   ao22f01 U264677 (.o(n247043),
	.a(n247042),
	.b(n247041),
	.c(regtop_g_udb0_r[5]),
	.d(n247040));
   in01s01 U264678 (.o(n211950),
	.a(n247038));
   ao22f01 U264679 (.o(n247038),
	.a(regtop_g_udb0_r[4]),
	.b(n247040),
	.c(n247042),
	.d(n247037));
   oa22f01 U264680 (.o(n211951),
	.a(n247034),
	.b(n246951),
	.c(n246954),
	.d(n246950));
   oa12f01 U264681 (.o(n211952),
	.a(n246906),
	.b(n246907),
	.c(n247034));
   oa22f01 U264682 (.o(n211953),
	.a(n247034),
	.b(n246955),
	.c(n246954),
	.d(n246953));
   oa22f01 U264683 (.o(n211954),
	.a(regtop_g_udb0_r[0]),
	.b(n246954),
	.c(n247034),
	.d(n246948));
   oa12f01 U264684 (.o(n211955),
	.a(n246940),
	.b(n246942),
	.c(n246941));
   ao22f01 U264685 (.o(n246881),
	.a(n246880),
	.b(n246879),
	.c(regtop_g_udb2_r[5]),
	.d(n246939));
   na02f01 U264686 (.o(n211957),
	.a(n246873),
	.b(n246872));
   na03f01 U264687 (.o(n246861),
	.a(n246880),
	.b(n246871),
	.c(n246860));
   ao22f01 U264688 (.o(n246878),
	.a(regtop_g_udb2_r[2]),
	.b(n246877),
	.c(n246876),
	.d(n246875));
   oa22s01 U264689 (.o(n211960),
	.a(n246852),
	.b(n246941),
	.c(n246870),
	.d(n246851));
   oa22s01 U264690 (.o(n211961),
	.a(regtop_g_udb2_r[0]),
	.b(n246941),
	.c(n246870),
	.d(n246062));
   ao22s01 U264691 (.o(n252369),
	.a(n252368),
	.b(n252377),
	.c(regtop_g_nfst_r[6]),
	.d(n252485));
   ao22s01 U264692 (.o(n252373),
	.a(n252377),
	.b(n252372),
	.c(regtop_g_nfst_r[4]),
	.d(n252485));
   oa12s01 U264693 (.o(n211966),
	.a(n246839),
	.b(n246840),
	.c(FE_OFN494_n252377));
   ao22s01 U264694 (.o(n252375),
	.a(n252377),
	.b(n252374),
	.c(n252485),
	.d(regtop_g_nfst_r[1]));
   ao22s01 U264695 (.o(n252378),
	.a(n252377),
	.b(n252376),
	.c(n252485),
	.d(regtop_g_nfst_r[9]));
   oa22s01 U264696 (.o(n252385),
	.a(n252401),
	.b(regtop_g_paramdata_r[10]),
	.c(regtop_g_fcho2_r[1]),
	.d(n252400));
   oa22s01 U264697 (.o(n252386),
	.a(n252401),
	.b(regtop_g_paramdata_r[11]),
	.c(regtop_g_fcho2_r[2]),
	.d(n252400));
   oa22s01 U264698 (.o(n252387),
	.a(n252401),
	.b(regtop_g_paramdata_r[12]),
	.c(regtop_g_fcho2_r[3]),
	.d(n252400));
   oa22s01 U264699 (.o(n252388),
	.a(n252401),
	.b(regtop_g_paramdata_r[13]),
	.c(regtop_g_fcho2_r[4]),
	.d(n252400));
   oa22s01 U264700 (.o(n252389),
	.a(n252401),
	.b(regtop_g_paramdata_r[14]),
	.c(regtop_g_fcho2_r[5]),
	.d(n252400));
   oa22s01 U264701 (.o(n252390),
	.a(n252401),
	.b(regtop_g_paramdata_r[15]),
	.c(regtop_g_fcho2_r[6]),
	.d(n252400));
   oa22s01 U264702 (.o(n252391),
	.a(n252401),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_fcho2_r[7]),
	.d(n252400));
   oa22s01 U264703 (.o(n252392),
	.a(n252401),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_fcho2_r[8]),
	.d(n252400));
   oa22s01 U264704 (.o(n252396),
	.a(n252401),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_fcho2_r[12]),
	.d(n252400));
   oa22s01 U264705 (.o(n252397),
	.a(n252401),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_fcho2_r[13]),
	.d(n252400));
   oa22s01 U264706 (.o(n252398),
	.a(n252401),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_fcho2_r[14]),
	.d(n252400));
   oa22s01 U264707 (.o(n252399),
	.a(n252401),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_fcho2_r[15]),
	.d(n252400));
   oa22s01 U264708 (.o(n252402),
	.a(n252401),
	.b(regtop_g_paramdata_r[9]),
	.c(regtop_g_fcho2_r[0]),
	.d(n252400));
   oa22s01 U264709 (.o(n252406),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[10]),
	.c(regtop_g_fcho0_r[1]),
	.d(n252421));
   oa22s01 U264710 (.o(n252407),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[11]),
	.c(regtop_g_fcho0_r[2]),
	.d(n252421));
   oa22s01 U264711 (.o(n252408),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[12]),
	.c(regtop_g_fcho0_r[3]),
	.d(n252421));
   oa22s01 U264712 (.o(n252409),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[13]),
	.c(regtop_g_fcho0_r[4]),
	.d(n252421));
   oa22s01 U264713 (.o(n252410),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[14]),
	.c(regtop_g_fcho0_r[5]),
	.d(n252421));
   oa22s01 U264714 (.o(n252411),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[15]),
	.c(regtop_g_fcho0_r[6]),
	.d(n252421));
   oa22s01 U264715 (.o(n252412),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_fcho0_r[7]),
	.d(n252421));
   oa22s01 U264716 (.o(n252414),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_fcho0_r[9]),
	.d(n252421));
   oa22s01 U264717 (.o(n252415),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_fcho0_r[10]),
	.d(n252421));
   oa22s01 U264718 (.o(n252416),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_fcho0_r[11]),
	.d(n252421));
   oa22s01 U264719 (.o(n252419),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_fcho0_r[14]),
	.d(n252421));
   oa22s01 U264720 (.o(n252420),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_fcho0_r[15]),
	.d(n252421));
   oa22s01 U264721 (.o(n252423),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[9]),
	.c(regtop_g_fcho0_r[0]),
	.d(n252421));
   oa22s01 U264722 (.o(n252450),
	.a(n252460),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_tr_r[1]),
	.d(n252459));
   oa22s01 U264723 (.o(n252452),
	.a(n252460),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_tr_r[3]),
	.d(n252459));
   oa22s01 U264724 (.o(n252453),
	.a(n252460),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_tr_r[4]),
	.d(n252459));
   oa22s01 U264725 (.o(n252454),
	.a(n252460),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_tr_r[5]),
	.d(n252459));
   oa22s01 U264726 (.o(n252455),
	.a(n252460),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_tr_r[6]),
	.d(n252459));
   oa22s01 U264727 (.o(n252456),
	.a(n252460),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_tr_r[7]),
	.d(n252459));
   oa22s01 U264728 (.o(n252457),
	.a(n252460),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_tr_r[8]),
	.d(n252459));
   oa22s01 U264729 (.o(n252458),
	.a(n252460),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_tr_r[9]),
	.d(n252459));
   oa22s01 U264730 (.o(n252461),
	.a(n252460),
	.b(regtop_g_paramdata_r[15]),
	.c(regtop_g_tr_r[0]),
	.d(n252459));
   in01s01 U264731 (.o(n246931),
	.a(n246933));
   in01s01 U264732 (.o(n212050),
	.a(n247054));
   ao22f01 U264733 (.o(n247054),
	.a(n247053),
	.b(n247052),
	.c(regtop_g_udb1_r[5]),
	.d(n247051));
   in01s01 U264734 (.o(n212051),
	.a(n247049));
   ao22f01 U264735 (.o(n247049),
	.a(regtop_g_udb1_r[4]),
	.b(n247051),
	.c(n247053),
	.d(n247048));
   oa22f01 U264736 (.o(n212052),
	.a(n247045),
	.b(n246958),
	.c(n246963),
	.d(n246957));
   oa12s01 U264737 (.o(n212053),
	.a(n246911),
	.b(n246912),
	.c(n247045));
   oa22f01 U264738 (.o(n212054),
	.a(n247045),
	.b(n246961),
	.c(n246963),
	.d(n246960));
   oa22f01 U264739 (.o(n212055),
	.a(regtop_g_udb1_r[0]),
	.b(n246963),
	.c(n247045),
	.d(n246962));
   oa22s01 U264740 (.o(n252492),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[10]),
	.c(regtop_g_fcho1_r[1]),
	.d(n252507));
   oa22s01 U264741 (.o(n252493),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[11]),
	.c(regtop_g_fcho1_r[2]),
	.d(n252507));
   oa22s01 U264742 (.o(n252494),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[12]),
	.c(regtop_g_fcho1_r[3]),
	.d(n252507));
   oa22s01 U264743 (.o(n252495),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[13]),
	.c(regtop_g_fcho1_r[4]),
	.d(n252507));
   oa22s01 U264744 (.o(n252496),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[14]),
	.c(regtop_g_fcho1_r[5]),
	.d(n252507));
   oa22s01 U264745 (.o(n252497),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[15]),
	.c(regtop_g_fcho1_r[6]),
	.d(n252507));
   oa22s01 U264746 (.o(n252498),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_fcho1_r[7]),
	.d(n252507));
   oa22s01 U264747 (.o(n252499),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_fcho1_r[8]),
	.d(n252507));
   oa22s01 U264748 (.o(n252502),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_fcho1_r[11]),
	.d(n252507));
   oa22s01 U264749 (.o(n252503),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_fcho1_r[12]),
	.d(n252507));
   oa22s01 U264750 (.o(n252505),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_fcho1_r[14]),
	.d(n252507));
   oa22s01 U264751 (.o(n252506),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_fcho1_r[15]),
	.d(n252507));
   oa22s01 U264752 (.o(n252509),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[9]),
	.c(regtop_g_fcho1_r[0]),
	.d(n252507));
   oa22s01 U264753 (.o(n252524),
	.a(n252540),
	.b(regtop_g_paramdata_r[10]),
	.c(regtop_g_vd_r[1]),
	.d(FE_OFN508_n252540));
   oa22s01 U264754 (.o(n252525),
	.a(n252540),
	.b(regtop_g_paramdata_r[11]),
	.c(regtop_g_vd_r[2]),
	.d(FE_OFN508_n252540));
   oa22s01 U264755 (.o(n252527),
	.a(n252540),
	.b(regtop_g_paramdata_r[13]),
	.c(regtop_g_vd_r[4]),
	.d(FE_OFN508_n252540));
   oa22s01 U264756 (.o(n252528),
	.a(n252540),
	.b(regtop_g_paramdata_r[14]),
	.c(regtop_g_vd_r[5]),
	.d(FE_OFN508_n252540));
   oa22s01 U264757 (.o(n252529),
	.a(n252540),
	.b(regtop_g_paramdata_r[15]),
	.c(regtop_g_vd_r[6]),
	.d(FE_OFN508_n252540));
   oa22s01 U264758 (.o(n252530),
	.a(n252540),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_vd_r[7]),
	.d(FE_OFN508_n252540));
   oa22s01 U264759 (.o(n252531),
	.a(n252540),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_vd_r[8]),
	.d(FE_OFN508_n252540));
   oa22s01 U264760 (.o(n252532),
	.a(n252540),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_vd_r[9]),
	.d(FE_OFN508_n252540));
   oa22s01 U264761 (.o(n252533),
	.a(n252540),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_vd_r[10]),
	.d(FE_OFN508_n252540));
   oa22s01 U264762 (.o(n252534),
	.a(n252540),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_vd_r[11]),
	.d(FE_OFN508_n252540));
   oa22s01 U264763 (.o(n252535),
	.a(n252540),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_vd_r[12]),
	.d(FE_OFN508_n252540));
   oa22s01 U264764 (.o(n252536),
	.a(n252540),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_vd_r[13]),
	.d(FE_OFN508_n252540));
   oa22s01 U264765 (.o(n252537),
	.a(n252540),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_vd_r[14]),
	.d(FE_OFN508_n252540));
   oa22s01 U264766 (.o(n252538),
	.a(n252540),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_vd_r[15]),
	.d(FE_OFN508_n252540));
   oa22s01 U264767 (.o(n252541),
	.a(n252540),
	.b(regtop_g_paramdata_r[9]),
	.c(regtop_g_vd_r[0]),
	.d(FE_OFN508_n252540));
   oa22s01 U264768 (.o(n212147),
	.a(n252580),
	.b(n252579),
	.c(n252581),
	.d(n252578));
   ao12s01 U264769 (.o(n252580),
	.a(n252577),
	.b(n252581),
	.c(n252595));
   oa22s01 U264770 (.o(n252614),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[10]),
	.c(regtop_g_fcvo1_r[1]),
	.d(n252629));
   oa22s01 U264771 (.o(n252615),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[11]),
	.c(regtop_g_fcvo1_r[2]),
	.d(n252629));
   oa22s01 U264772 (.o(n252616),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[12]),
	.c(regtop_g_fcvo1_r[3]),
	.d(n252629));
   oa22s01 U264773 (.o(n252617),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[13]),
	.c(regtop_g_fcvo1_r[4]),
	.d(n252629));
   oa22s01 U264774 (.o(n252618),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[14]),
	.c(regtop_g_fcvo1_r[5]),
	.d(n252629));
   oa22s01 U264775 (.o(n252619),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[15]),
	.c(regtop_g_fcvo1_r[6]),
	.d(n252629));
   oa22s01 U264776 (.o(n252620),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_fcvo1_r[7]),
	.d(n252629));
   oa22s01 U264777 (.o(n252621),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_fcvo1_r[8]),
	.d(n252629));
   oa22s01 U264778 (.o(n252622),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_fcvo1_r[9]),
	.d(n252629));
   oa22s01 U264779 (.o(n252623),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_fcvo1_r[10]),
	.d(n252629));
   oa22s01 U264780 (.o(n252624),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_fcvo1_r[11]),
	.d(n252629));
   oa22s01 U264781 (.o(n252625),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_fcvo1_r[12]),
	.d(n252629));
   oa22s01 U264782 (.o(n252626),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_fcvo1_r[13]),
	.d(n252629));
   oa22s01 U264783 (.o(n252628),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_fcvo1_r[15]),
	.d(n252629));
   oa22s01 U264784 (.o(n252631),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[9]),
	.c(regtop_g_fcvo1_r[0]),
	.d(n252629));
   oa12s01 U264785 (.o(n212201),
	.a(n246003),
	.b(n252682),
	.c(n252676));
   oa22s01 U264786 (.o(n252701),
	.a(n252704),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_pct_r[1]),
	.d(n252703));
   oa22s01 U264787 (.o(n252702),
	.a(n252704),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_pct_r[2]),
	.d(n252703));
   oa22s01 U264788 (.o(n252705),
	.a(n252704),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_pct_r[0]),
	.d(n252703));
   oa22s01 U264789 (.o(n252713),
	.a(n252728),
	.b(regtop_g_paramdata_r[11]),
	.c(regtop_g_fcvo0_r[2]),
	.d(n252727));
   oa22s01 U264790 (.o(n252714),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[12]),
	.c(regtop_g_fcvo0_r[3]),
	.d(n252727));
   oa22s01 U264791 (.o(n252715),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[13]),
	.c(regtop_g_fcvo0_r[4]),
	.d(n252727));
   oa22s01 U264792 (.o(n252716),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[14]),
	.c(regtop_g_fcvo0_r[5]),
	.d(n252727));
   oa22s01 U264793 (.o(n252717),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[15]),
	.c(regtop_g_fcvo0_r[6]),
	.d(n252727));
   oa22s01 U264794 (.o(n252718),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_fcvo0_r[7]),
	.d(n252727));
   oa22s01 U264795 (.o(n252719),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_fcvo0_r[8]),
	.d(n252727));
   oa22s01 U264796 (.o(n252720),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_fcvo0_r[9]),
	.d(n252727));
   oa22s01 U264797 (.o(n252721),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_fcvo0_r[10]),
	.d(n252727));
   oa22s01 U264798 (.o(n252722),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_fcvo0_r[11]),
	.d(n252727));
   oa22s01 U264799 (.o(n252723),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_fcvo0_r[12]),
	.d(n252727));
   oa22s01 U264800 (.o(n252724),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_fcvo0_r[13]),
	.d(n252727));
   oa22s01 U264801 (.o(n252725),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_fcvo0_r[14]),
	.d(n252727));
   oa22s01 U264802 (.o(n252726),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_fcvo0_r[15]),
	.d(n252727));
   oa22s01 U264803 (.o(n252732),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[10]),
	.c(regtop_g_fcvo2_r[1]),
	.d(n252747));
   oa22s01 U264804 (.o(n252733),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[11]),
	.c(regtop_g_fcvo2_r[2]),
	.d(n252747));
   oa22s01 U264805 (.o(n252734),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[12]),
	.c(regtop_g_fcvo2_r[3]),
	.d(n252747));
   oa22s01 U264806 (.o(n252735),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[13]),
	.c(regtop_g_fcvo2_r[4]),
	.d(n252747));
   oa22s01 U264807 (.o(n252736),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[14]),
	.c(regtop_g_fcvo2_r[5]),
	.d(n252747));
   oa22s01 U264808 (.o(n252737),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[15]),
	.c(regtop_g_fcvo2_r[6]),
	.d(n252747));
   oa22s01 U264809 (.o(n252738),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_fcvo2_r[7]),
	.d(n252747));
   oa22s01 U264810 (.o(n252739),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_fcvo2_r[8]),
	.d(n252747));
   oa22s01 U264811 (.o(n252740),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_fcvo2_r[9]),
	.d(n252747));
   oa22s01 U264812 (.o(n252741),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_fcvo2_r[10]),
	.d(n252747));
   oa22s01 U264813 (.o(n252742),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_fcvo2_r[11]),
	.d(n252747));
   oa22s01 U264814 (.o(n252743),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_fcvo2_r[12]),
	.d(n252747));
   oa22s01 U264815 (.o(n252744),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_fcvo2_r[13]),
	.d(n252747));
   oa22s01 U264816 (.o(n252745),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_fcvo2_r[14]),
	.d(n252747));
   oa22s01 U264817 (.o(n252749),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[9]),
	.c(regtop_g_fcvo2_r[0]),
	.d(n252747));
   oa12s01 U264818 (.o(n252787),
	.a(n252786),
	.b(n252788),
	.c(n252811));
   oa22s01 U264819 (.o(n246754),
	.a(FE_OFN6_n246618),
	.b(n246753),
	.c(n252656),
	.d(n246773));
   oa22s01 U264820 (.o(n246750),
	.a(FE_OFN6_n246618),
	.b(n246749),
	.c(n252658),
	.d(n246773));
   oa22s01 U264821 (.o(n246775),
	.a(FE_OFN6_n246618),
	.b(n246774),
	.c(n252660),
	.d(n246773));
   oa22s01 U264822 (.o(n246770),
	.a(FE_OFN6_n246618),
	.b(n246769),
	.c(n252662),
	.d(n246773));
   oa22s01 U264823 (.o(n246766),
	.a(FE_OFN6_n246618),
	.b(n246765),
	.c(n252664),
	.d(n246773));
   oa22s01 U264824 (.o(n246758),
	.a(FE_OFN6_n246618),
	.b(n246757),
	.c(n252666),
	.d(n246773));
   oa22s01 U264825 (.o(n246762),
	.a(FE_OFN6_n246618),
	.b(n246761),
	.c(n252778),
	.d(n246773));
   oa22s01 U264826 (.o(n246746),
	.a(FE_OFN6_n246618),
	.b(n246745),
	.c(n252755),
	.d(n246773));
   na02s01 U264827 (.o(n246429),
	.a(g_swrst_r_n),
	.b(n246428));
   na02f01 U264828 (.o(n246059),
	.a(vldtop_vld_syndec_vld_seqhed_state_0_),
	.b(n246058));
   ao22f01 U264829 (.o(n246058),
	.a(n246025),
	.b(n247000),
	.c(n246057),
	.d(n247002));
   oa22s01 U264830 (.o(n243166),
	.a(n249063),
	.b(n249022),
	.c(n249028),
	.d(n246898));
   oa22s01 U264831 (.o(n243167),
	.a(n249026),
	.b(n249022),
	.c(n249028),
	.d(n249021));
   oa22s01 U264832 (.o(n212465),
	.a(n249063),
	.b(n249060),
	.c(n249028),
	.d(n249027));
   oa22s01 U264833 (.o(n252835),
	.a(n252834),
	.b(regtop_g_wd_r[16]),
	.c(g_vs60p_r[0]),
	.d(FE_OFN454_n252863));
   ao22s01 U264834 (.o(n212535),
	.a(FE_OFN454_n252863),
	.b(n252901),
	.c(n252836),
	.d(n252834));
   oa22s01 U264835 (.o(n252837),
	.a(n252834),
	.b(regtop_g_wd_r[21]),
	.c(g_vs60p_r[5]),
	.d(FE_OFN454_n252863));
   oa22s01 U264836 (.o(n252839),
	.a(n252834),
	.b(regtop_g_wd_r[19]),
	.c(g_vs60p_r[3]),
	.d(FE_OFN454_n252863));
   ao22s01 U264837 (.o(n212539),
	.a(FE_OFN454_n252863),
	.b(n252894),
	.c(n252840),
	.d(n252834));
   ao22s01 U264838 (.o(n212540),
	.a(FE_OFN454_n252863),
	.b(n252915),
	.c(n252841),
	.d(n252834));
   oa22s01 U264839 (.o(n252842),
	.a(n252834),
	.b(regtop_g_wd_r[24]),
	.c(g_hs60p_r[0]),
	.d(FE_OFN454_n252863));
   ao22s01 U264840 (.o(n212542),
	.a(FE_OFN454_n252863),
	.b(n252844),
	.c(n252843),
	.d(n252834));
   oa22s01 U264841 (.o(n252845),
	.a(n252834),
	.b(regtop_g_wd_r[29]),
	.c(g_hs60p_r[5]),
	.d(FE_OFN454_n252863));
   oa22s01 U264842 (.o(n252846),
	.a(n252834),
	.b(regtop_g_wd_r[28]),
	.c(g_hs60p_r[4]),
	.d(FE_OFN454_n252863));
   ao22s01 U264843 (.o(n212545),
	.a(FE_OFN454_n252863),
	.b(n252909),
	.c(n252847),
	.d(n252834));
   oa22s01 U264844 (.o(n252848),
	.a(n252834),
	.b(regtop_g_wd_r[26]),
	.c(g_hs60p_r[2]),
	.d(FE_OFN454_n252863));
   oa22s01 U264845 (.o(n252849),
	.a(n252834),
	.b(regtop_g_wd_r[25]),
	.c(g_hs60p_r[1]),
	.d(FE_OFN454_n252863));
   ao22s01 U264846 (.o(n212548),
	.a(FE_OFN454_n252863),
	.b(n252953),
	.c(n252850),
	.d(n252834));
   ao22s01 U264847 (.o(n212549),
	.a(FE_OFN454_n252863),
	.b(n252885),
	.c(n252851),
	.d(n252834));
   oa22s01 U264848 (.o(n252852),
	.a(n252834),
	.b(regtop_g_wd_r[5]),
	.c(g_vsdc_r[5]),
	.d(FE_OFN454_n252863));
   oa22s01 U264849 (.o(n252853),
	.a(n252834),
	.b(regtop_g_wd_r[4]),
	.c(g_vsdc_r[4]),
	.d(FE_OFN454_n252863));
   ao22s01 U264850 (.o(n212552),
	.a(FE_OFN454_n252863),
	.b(n253002),
	.c(n252854),
	.d(n252834));
   oa22s01 U264851 (.o(n252855),
	.a(n252834),
	.b(regtop_g_wd_r[2]),
	.c(g_vsdc_r[2]),
	.d(FE_OFN454_n252863));
   oa22s01 U264852 (.o(n252856),
	.a(n252834),
	.b(regtop_g_wd_r[1]),
	.c(g_vsdc_r[1]),
	.d(FE_OFN454_n252863));
   oa22s01 U264853 (.o(n252857),
	.a(n252834),
	.b(regtop_g_wd_r[9]),
	.c(g_hsdc_r[1]),
	.d(FE_OFN454_n252863));
   oa22s01 U264854 (.o(n252858),
	.a(n252834),
	.b(regtop_g_wd_r[10]),
	.c(g_hsdc_r[2]),
	.d(FE_OFN454_n252863));
   oa22s01 U264855 (.o(n252860),
	.a(n252834),
	.b(regtop_g_wd_r[12]),
	.c(g_hsdc_r[4]),
	.d(FE_OFN454_n252863));
   oa22s01 U264856 (.o(n252861),
	.a(n252834),
	.b(regtop_g_wd_r[13]),
	.c(g_hsdc_r[5]),
	.d(FE_OFN454_n252863));
   oa22s01 U264857 (.o(n252865),
	.a(n252834),
	.b(regtop_g_wd_r[8]),
	.c(g_hsdc_r[0]),
	.d(FE_OFN454_n252863));
   oa22s01 U264858 (.o(n212576),
	.a(n246838),
	.b(n246670),
	.c(n246837),
	.d(n246836));
   ao22s01 U264859 (.o(n246837),
	.a(n246835),
	.b(n246834),
	.c(n246833),
	.d(n246832));
   ao12f01 U264860 (.o(n253071),
	.a(n247161),
	.b(n247162),
	.c(n247126));
   na02f01 U264861 (.o(n212582),
	.a(n247271),
	.b(n247270));
   ao12f01 U264862 (.o(n247271),
	.a(FE_OFN68_n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[31]));
   ao22f01 U264863 (.o(n247270),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[31]),
	.b(n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[31]));
   ao12f01 U264864 (.o(n253072),
	.a(n247165),
	.b(n247166),
	.c(FE_OCPN583_n247126));
   na02f01 U264865 (.o(n212584),
	.a(n247219),
	.b(n247218));
   ao22f01 U264866 (.o(n247218),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[30]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[30]));
   ao12f01 U264867 (.o(n253073),
	.a(n247291),
	.b(n247292),
	.c(n247126));
   na02f01 U264868 (.o(n212586),
	.a(n247168),
	.b(n247167));
   ao22f01 U264869 (.o(n247167),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[29]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[29]));
   ao12f01 U264870 (.o(n253074),
	.a(n247334),
	.b(n247335),
	.c(FE_OCPN583_n247126));
   na02f01 U264871 (.o(n212588),
	.a(n247352),
	.b(n247351));
   ao12f01 U264872 (.o(n247352),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[28]));
   ao22f01 U264873 (.o(n247351),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[28]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[28]));
   ao12f01 U264874 (.o(n253075),
	.a(n247212),
	.b(n247213),
	.c(FE_OCPN583_n247126));
   na02f01 U264875 (.o(n212590),
	.a(n247257),
	.b(n247256));
   ao12f01 U264876 (.o(n247257),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[27]));
   ao12f01 U264877 (.o(n253076),
	.a(n247242),
	.b(n247243),
	.c(FE_OCPN583_n247126));
   ao12f01 U264878 (.o(n247373),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[26]));
   ao22f01 U264879 (.o(n247372),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[26]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[26]));
   ao12f01 U264880 (.o(n253077),
	.a(n247133),
	.b(n247134),
	.c(FE_OFN577_n247126));
   ao12f01 U264881 (.o(n247154),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[25]));
   ao12f01 U264882 (.o(n253078),
	.a(n247370),
	.b(n247371),
	.c(FE_OCPN583_n247126));
   na02f01 U264883 (.o(n212596),
	.a(n247205),
	.b(n247204));
   ao12f01 U264884 (.o(n247205),
	.a(FE_OFN68_n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[24]));
   ao12f01 U264885 (.o(n253079),
	.a(n247295),
	.b(n247296),
	.c(FE_OFN577_n247126));
   na02f01 U264886 (.o(n212598),
	.a(n247305),
	.b(n247304));
   ao12f01 U264887 (.o(n247305),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[23]));
   ao12f01 U264888 (.o(n253080),
	.a(n247278),
	.b(n247279),
	.c(FE_OCPN583_n247126));
   na02f01 U264889 (.o(n212600),
	.a(n247251),
	.b(n247250));
   ao12f01 U264890 (.o(n253081),
	.a(n247129),
	.b(n247130),
	.c(FE_OFN577_n247126));
   na02f01 U264891 (.o(n212602),
	.a(n247188),
	.b(n247187));
   ao12f01 U264892 (.o(n247188),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[21]));
   ao12f01 U264893 (.o(n253082),
	.a(n247175),
	.b(n247176),
	.c(FE_OCPN583_n247126));
   na02f01 U264894 (.o(n212604),
	.a(n247178),
	.b(n247177));
   ao12f01 U264895 (.o(n247178),
	.a(FE_OFN68_n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[20]));
   ao12f01 U264896 (.o(n253083),
	.a(n247366),
	.b(n247367),
	.c(FE_OCPN583_n247126));
   na02f01 U264897 (.o(n212606),
	.a(n247253),
	.b(n247252));
   ao12f01 U264898 (.o(n247253),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[19]));
   ao22f01 U264899 (.o(n247252),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[19]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[19]));
   ao12f01 U264900 (.o(n247209),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[18]));
   ao12f01 U264901 (.o(n253085),
	.a(n247197),
	.b(n247198),
	.c(FE_OCPN583_n247126));
   na02f01 U264902 (.o(n212610),
	.a(n247355),
	.b(n247354));
   ao12f01 U264903 (.o(n253086),
	.a(n247185),
	.b(n247186),
	.c(FE_OCPN583_n247126));
   na02f01 U264904 (.o(n212612),
	.a(n247247),
	.b(n247246));
   ao12f01 U264905 (.o(n253087),
	.a(n247201),
	.b(n247202),
	.c(FE_OFN577_n247126));
   na02f01 U264906 (.o(n212614),
	.a(n247383),
	.b(n247382));
   ao12f01 U264907 (.o(n247383),
	.a(FE_OFN68_n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[15]));
   ao12f01 U264908 (.o(n253088),
	.a(n247318),
	.b(n247319),
	.c(FE_OCPN583_n247126));
   na02f01 U264909 (.o(n212616),
	.a(n247221),
	.b(n247220));
   ao12f01 U264910 (.o(n247221),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[14]));
   ao12f01 U264911 (.o(n253089),
	.a(n247171),
	.b(n247172),
	.c(FE_OCPN583_n247126));
   na02f01 U264912 (.o(n212618),
	.a(n247249),
	.b(n247248));
   ao12f01 U264913 (.o(n253090),
	.a(n247157),
	.b(n247158),
	.c(FE_OCPN583_n247126));
   na02f01 U264914 (.o(n212620),
	.a(n247207),
	.b(n247206));
   ao12f01 U264915 (.o(n247207),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[12]));
   ao12s01 U264916 (.o(n253091),
	.a(n247314),
	.b(n247315),
	.c(FE_OFN577_n247126));
   ao12f01 U264917 (.o(n247263),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[11]));
   ao22f01 U264918 (.o(n247262),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[11]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[11]));
   ao12f01 U264919 (.o(n253092),
	.a(n247224),
	.b(n247225),
	.c(FE_OCPN583_n247126));
   ao22f01 U264920 (.o(n247306),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[10]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[10]));
   ao12f01 U264921 (.o(n253093),
	.a(n247266),
	.b(n247267),
	.c(FE_OCPN583_n247126));
   na02f01 U264922 (.o(n212626),
	.a(n247300),
	.b(n247299));
   ao12f01 U264923 (.o(n247300),
	.a(FE_OFN68_n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[9]));
   ao12f01 U264924 (.o(n253094),
	.a(n247260),
	.b(n247261),
	.c(FE_OCPN583_n247126));
   na02f01 U264925 (.o(n212628),
	.a(n247227),
	.b(n247226));
   ao22f01 U264926 (.o(n247226),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[8]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[8]));
   ao12s01 U264927 (.o(n253095),
	.a(n247216),
	.b(n247217),
	.c(n247126));
   na02f01 U264928 (.o(n212630),
	.a(n247152),
	.b(n247151));
   ao22f01 U264929 (.o(n247151),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[7]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[7]));
   ao12f01 U264930 (.o(n253096),
	.a(n247141),
	.b(n247142),
	.c(FE_OCPN583_n247126));
   na02f01 U264931 (.o(n212632),
	.a(n247337),
	.b(n247336));
   ao12f01 U264932 (.o(n247337),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[6]));
   ao12f01 U264933 (.o(n253097),
	.a(n247230),
	.b(n247231),
	.c(FE_OFN577_n247126));
   na02f01 U264934 (.o(n212634),
	.a(n247329),
	.b(n247328));
   ao22f01 U264935 (.o(n247328),
	.a(FE_OFN14_n247150),
	.b(vldtop_vld_syndec_vld_vlfeed_temporal[5]),
	.c(vldtop_vld_syndec_vld_vlfeed_lower[5]),
	.d(FE_OFN577_n247126));
   ao12f01 U264936 (.o(n253098),
	.a(n247181),
	.b(n247182),
	.c(n247126));
   na02f01 U264937 (.o(n212636),
	.a(n247331),
	.b(n247330));
   ao12f01 U264938 (.o(n247331),
	.a(FE_OFN68_n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[4]));
   na02f01 U264939 (.o(n212638),
	.a(n247302),
	.b(n247301));
   ao12f01 U264940 (.o(n247302),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[3]));
   ao12f01 U264941 (.o(n253100),
	.a(n247310),
	.b(n247311),
	.c(n247126));
   na02f01 U264942 (.o(n212640),
	.a(n247269),
	.b(n247268));
   ao12f01 U264943 (.o(n247269),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[2]));
   ao12f01 U264944 (.o(n253101),
	.a(n247286),
	.b(n247288),
	.c(n247126));
   na02f01 U264945 (.o(n212642),
	.a(n247245),
	.b(n247244));
   ao12f01 U264946 (.o(n253102),
	.a(n247297),
	.b(n247298),
	.c(n247126));
   na02f01 U264947 (.o(n212644),
	.a(n247190),
	.b(n247189));
   no02f01 U264948 (.o(n253039),
	.a(n247285),
	.b(n247284));
   in01s01 U264949 (.o(n247285),
	.a(n247283));
   na03f01 U264950 (.o(n247283),
	.a(g_swrst_r_n),
	.b(n247494),
	.c(n247282));
   no02f01 U264951 (.o(n253043),
	.a(n247281),
	.b(n247280));
   na03f02 U264952 (.o(n247451),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247450));
   no02f01 U264953 (.o(n253045),
	.a(n247449),
	.b(n247448));
   in01s01 U264954 (.o(n247449),
	.a(n247447));
   na03s02 U264955 (.o(n247447),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247446));
   no02s01 U264956 (.o(n253046),
	.a(n247466),
	.b(n247465));
   in01s01 U264957 (.o(n247466),
	.a(n247464));
   na03f01 U264958 (.o(n247464),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247494),
	.c(n247463));
   no02f01 U264959 (.o(n253049),
	.a(n247593),
	.b(n247592));
   in01s01 U264960 (.o(n247593),
	.a(n247590));
   na03s02 U264961 (.o(n247590),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247589));
   na03f01 U264962 (.o(n247460),
	.a(FE_OFN2_g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247459));
   na03s02 U264963 (.o(n247361),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247360));
   no02f01 U264964 (.o(n253057),
	.a(n247341),
	.b(n247340));
   na03s02 U264965 (.o(n247339),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247338));
   no02f01 U264966 (.o(n253059),
	.a(n247445),
	.b(n247444));
   in01s01 U264967 (.o(n247445),
	.a(n247443));
   na03s02 U264968 (.o(n247443),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247442));
   no02f01 U264969 (.o(n253060),
	.a(n247239),
	.b(n247238));
   in01s01 U264970 (.o(n247239),
	.a(n247237));
   na03f01 U264971 (.o(n247237),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247236));
   no02s01 U264972 (.o(n253061),
	.a(n246857),
	.b(n246856));
   in01s01 U264973 (.o(n246857),
	.a(n246855));
   na03f01 U264974 (.o(n246855),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247494),
	.c(n246854));
   in01s01 U264975 (.o(n247458),
	.a(n247456));
   na03s02 U264976 (.o(n247456),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247455));
   no02f01 U264977 (.o(n253066),
	.a(n247482),
	.b(n247481));
   in01s01 U264978 (.o(n247482),
	.a(n247480));
   na03f01 U264979 (.o(n247480),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247494),
	.c(n247479));
   no02f01 U264980 (.o(n253067),
	.a(n247235),
	.b(n247234));
   in01s01 U264981 (.o(n247235),
	.a(n247233));
   na03s02 U264982 (.o(n247233),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247232));
   no02f01 U264983 (.o(n253068),
	.a(n247588),
	.b(n247587));
   in01s01 U264984 (.o(n247588),
	.a(n247586));
   no02f01 U264985 (.o(n253069),
	.a(n247381),
	.b(n247380));
   in01s01 U264986 (.o(n247381),
	.a(n247379));
   no02f01 U264987 (.o(n253070),
	.a(n247377),
	.b(n247376));
   in01s01 U264988 (.o(n247377),
	.a(n247375));
   na03s02 U264989 (.o(n247375),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247374));
   oa22s01 U264990 (.o(n212677),
	.a(n246838),
	.b(n247145),
	.c(n247143),
	.d(n246836));
   oa12s01 U264991 (.o(n212678),
	.a(n246825),
	.b(n247143),
	.c(n247146));
   oa22s01 U264992 (.o(n252902),
	.a(FE_OFN441_n252905),
	.b(regtop_g_wd_r[23]),
	.c(g_pcut_r[7]),
	.d(n252875));
   oa22s01 U264993 (.o(n252951),
	.a(n252954),
	.b(regtop_g_wd_r[1]),
	.c(g_bmod_r),
	.d(n252957));
   oa22s01 U264994 (.o(n252973),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[11]),
	.c(g_field_start_add_r[11]),
	.d(n252995));
   oa22s01 U264995 (.o(n252974),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[12]),
	.c(g_field_start_add_r[12]),
	.d(n252995));
   oa22s01 U264996 (.o(n252975),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[13]),
	.c(g_field_start_add_r[13]),
	.d(n252995));
   oa22s01 U264997 (.o(n252976),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[14]),
	.c(g_field_start_add_r[14]),
	.d(n252995));
   oa22s01 U264998 (.o(n252977),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[15]),
	.c(g_field_start_add_r[15]),
	.d(n252995));
   oa22s01 U264999 (.o(n252978),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[16]),
	.c(g_field_start_add_r[16]),
	.d(n252995));
   oa22s01 U265000 (.o(n252979),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[17]),
	.c(g_field_start_add_r[17]),
	.d(n252995));
   oa22s01 U265001 (.o(n252980),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[18]),
	.c(g_field_start_add_r[18]),
	.d(n252995));
   oa22s01 U265002 (.o(n252981),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[19]),
	.c(g_field_start_add_r[19]),
	.d(n252995));
   ao22s01 U265003 (.o(n212751),
	.a(n252995),
	.b(n252983),
	.c(n252982),
	.d(FE_OFN458_n252996));
   oa22s01 U265004 (.o(n252984),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[21]),
	.c(g_field_start_add_r[21]),
	.d(n252995));
   oa22s01 U265005 (.o(n252985),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[22]),
	.c(g_field_start_add_r[22]),
	.d(n252995));
   oa22s01 U265006 (.o(n252986),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[23]),
	.c(g_field_start_add_r[23]),
	.d(n252995));
   oa22s01 U265007 (.o(n252987),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[24]),
	.c(g_field_start_add_r[24]),
	.d(n252995));
   oa22s01 U265008 (.o(n252988),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[25]),
	.c(g_field_start_add_r[25]),
	.d(n252995));
   oa22s01 U265009 (.o(n252989),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[26]),
	.c(g_field_start_add_r[26]),
	.d(n252995));
   oa22s01 U265010 (.o(n252990),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[27]),
	.c(g_field_start_add_r[27]),
	.d(n252995));
   oa22s01 U265011 (.o(n252991),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[28]),
	.c(g_field_start_add_r[28]),
	.d(n252995));
   oa22s01 U265012 (.o(n252992),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[29]),
	.c(g_field_start_add_r[29]),
	.d(n252995));
   oa22s01 U265013 (.o(n252993),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[30]),
	.c(g_field_start_add_r[30]),
	.d(n252995));
   oa22s01 U265014 (.o(n252994),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[31]),
	.c(g_field_start_add_r[31]),
	.d(n252995));
   oa22s01 U265015 (.o(n252997),
	.a(FE_OFN458_n252996),
	.b(regtop_g_wd_r[10]),
	.c(g_field_start_add_r[10]),
	.d(n252995));
   oa22s01 U265016 (.o(n252999),
	.a(n253012),
	.b(regtop_g_wd_r[1]),
	.c(g_field_offset_r[1]),
	.d(n253011));
   oa22s01 U265017 (.o(n253000),
	.a(n253012),
	.b(regtop_g_wd_r[2]),
	.c(g_field_offset_r[2]),
	.d(n253011));
   oa22s01 U265018 (.o(n253003),
	.a(n253012),
	.b(regtop_g_wd_r[4]),
	.c(g_field_offset_r[4]),
	.d(n253011));
   oa22s01 U265019 (.o(n253006),
	.a(n253012),
	.b(regtop_g_wd_r[7]),
	.c(g_field_offset_r[7]),
	.d(n253011));
   oa22s01 U265020 (.o(n253007),
	.a(n253012),
	.b(regtop_g_wd_r[8]),
	.c(g_field_offset_r[8]),
	.d(n253011));
   oa22s01 U265021 (.o(n253008),
	.a(n253012),
	.b(regtop_g_wd_r[9]),
	.c(g_field_offset_r[9]),
	.d(n253011));
   oa22s01 U265022 (.o(n253009),
	.a(n253012),
	.b(regtop_g_wd_r[10]),
	.c(g_field_offset_r[10]),
	.d(n253011));
   oa22s01 U265023 (.o(n253010),
	.a(n253012),
	.b(regtop_g_wd_r[11]),
	.c(g_field_offset_r[11]),
	.d(n253011));
   oa22s01 U265024 (.o(n253013),
	.a(n253012),
	.b(regtop_g_wd_r[0]),
	.c(g_field_offset_r[0]),
	.d(n253011));
   oa22s01 U265025 (.o(n253016),
	.a(n253029),
	.b(regtop_g_wd_r[1]),
	.c(g_cbcr_offset_r[1]),
	.d(n253028));
   oa22s01 U265026 (.o(n253017),
	.a(n253029),
	.b(regtop_g_wd_r[2]),
	.c(g_cbcr_offset_r[2]),
	.d(n253028));
   oa22s01 U265027 (.o(n253018),
	.a(n253029),
	.b(regtop_g_wd_r[3]),
	.c(g_cbcr_offset_r[3]),
	.d(n253028));
   oa22s01 U265028 (.o(n253019),
	.a(n253029),
	.b(regtop_g_wd_r[4]),
	.c(g_cbcr_offset_r[4]),
	.d(n253028));
   oa22s01 U265029 (.o(n253020),
	.a(n253029),
	.b(regtop_g_wd_r[5]),
	.c(g_cbcr_offset_r[5]),
	.d(n253028));
   oa22s01 U265030 (.o(n253021),
	.a(n253029),
	.b(regtop_g_wd_r[6]),
	.c(g_cbcr_offset_r[6]),
	.d(n253028));
   oa22s01 U265031 (.o(n253024),
	.a(n253029),
	.b(regtop_g_wd_r[8]),
	.c(g_cbcr_offset_r[8]),
	.d(n253028));
   oa22s01 U265032 (.o(n253026),
	.a(n253029),
	.b(regtop_g_wd_r[10]),
	.c(g_cbcr_offset_r[10]),
	.d(n253028));
   oa22s01 U265033 (.o(n253027),
	.a(n253029),
	.b(regtop_g_wd_r[11]),
	.c(g_cbcr_offset_r[11]),
	.d(n253028));
   oa22s01 U265034 (.o(n253030),
	.a(n253029),
	.b(regtop_g_wd_r[0]),
	.c(g_cbcr_offset_r[0]),
	.d(n253028));
   na02f02 U265035 (.o(regtop_w1_hdi00_q[31]),
	.a(n248845),
	.b(n248844));
   no04f02 U265036 (.o(n248845),
	.a(n248823),
	.b(n248822),
	.c(n248821),
	.d(FE_OFN579_n248820));
   no04f06 U265037 (.o(n248844),
	.a(FE_OFN256_n248843),
	.b(n248842),
	.c(n248841),
	.d(n248840));
   na04f01 U265038 (.o(n248820),
	.a(n248819),
	.b(n248818),
	.c(n248817),
	.d(n248816));
   no04f03 U265040 (.o(n248185),
	.a(n248184),
	.b(n248183),
	.c(n248182),
	.d(n248181));
   na04f04 U265041 (.o(n248184),
	.a(n248157),
	.b(n248156),
	.c(n248155),
	.d(n248154));
   no04f04 U265042 (.o(n247583),
	.a(n247582),
	.b(n247581),
	.c(n247580),
	.d(n247579));
   no04f02 U265043 (.o(n247541),
	.a(n247540),
	.b(n247539),
	.c(FE_OFN514_n247538),
	.d(n247537));
   na04f03 U265044 (.o(n247539),
	.a(n247526),
	.b(n247525),
	.c(n247524),
	.d(n247523));
   no04f06 U265045 (.o(n247439),
	.a(n247438),
	.b(n247437),
	.c(n247436),
	.d(n247435));
   no04f04 U265046 (.o(n248425),
	.a(n248390),
	.b(FE_OFN240_n248389),
	.c(n248388),
	.d(n248387));
   no04f04 U265047 (.o(n247864),
	.a(n247863),
	.b(n247862),
	.c(n247861),
	.d(n247860));
   na04f02 U265048 (.o(n247860),
	.a(n247859),
	.b(n247858),
	.c(n247857),
	.d(n247856));
   no04f02 U265049 (.o(n248312),
	.a(n248290),
	.b(n248289),
	.c(n248288),
	.d(n248287));
   no04f02 U265050 (.o(n248311),
	.a(n248310),
	.b(n248309),
	.c(n248308),
	.d(n248307));
   na04f02 U265051 (.o(n248290),
	.a(n248274),
	.b(n248273),
	.c(n248272),
	.d(n248271));
   na04s02 U265052 (.o(n248896),
	.a(n248869),
	.b(n248868),
	.c(n248867),
	.d(n248866));
   na02f02 U265053 (.o(regtop_w1_hdi00_q[20]),
	.a(n248509),
	.b(FE_OFN522_n248508));
   no04f01 U265054 (.o(n248509),
	.a(n248487),
	.b(n248486),
	.c(n248485),
	.d(n248484));
   no04f02 U265055 (.o(n248508),
	.a(n248507),
	.b(n248506),
	.c(n248505),
	.d(n248504));
   na04f03 U265056 (.o(n248486),
	.a(n248475),
	.b(n248474),
	.c(n248473),
	.d(n248472));
   no04f04 U265057 (.o(n247991),
	.a(n247969),
	.b(n247968),
	.c(n247967),
	.d(n247966));
   no04f03 U265058 (.o(n247990),
	.a(n247989),
	.b(n247988),
	.c(FE_OFN230_n247987),
	.d(n247986));
   na04f02 U265059 (.o(n247968),
	.a(n247957),
	.b(n247956),
	.c(n247955),
	.d(n247954));
   no04f03 U265060 (.o(n247697),
	.a(n247649),
	.b(n247648),
	.c(n247647),
	.d(n247646));
   na04f01 U265061 (.o(n247647),
	.a(n247635),
	.b(n247634),
	.c(n247633),
	.d(n247632));
   no04f02 U265062 (.o(n247739),
	.a(n247717),
	.b(n247716),
	.c(n247715),
	.d(n247714));
   no04f02 U265063 (.o(n247738),
	.a(FE_OFN372_n247737),
	.b(n247736),
	.c(n247735),
	.d(n247734));
   na04f03 U265064 (.o(n247716),
	.a(n247705),
	.b(n247704),
	.c(n247703),
	.d(n247702));
   no04f03 U265065 (.o(n247781),
	.a(n247759),
	.b(n247758),
	.c(n247757),
	.d(n247756));
   na04f04 U265066 (.o(n247756),
	.a(n247755),
	.b(n247754),
	.c(n247753),
	.d(n247752));
   no04f03 U265067 (.o(n247823),
	.a(n247801),
	.b(n247800),
	.c(n247799),
	.d(n247798));
   no04f03 U265068 (.o(n247906),
	.a(n247905),
	.b(n247904),
	.c(FE_OFN228_n247903),
	.d(n247902));
   na04f06 U265069 (.o(n247905),
	.a(n247889),
	.b(n247888),
	.c(n247887),
	.d(n247886));
   no04s02 U265070 (.o(n247949),
	.a(n247927),
	.b(n247926),
	.c(n247925),
	.d(n247924));
   no04f06 U265071 (.o(n247948),
	.a(n247947),
	.b(n247946),
	.c(n247945),
	.d(n247944));
   na04f02 U265072 (.o(n247926),
	.a(n247915),
	.b(n247914),
	.c(n247913),
	.d(n247912));
   no04f04 U265073 (.o(n248466),
	.a(FE_OFN246_n248465),
	.b(n248464),
	.c(FE_OFN244_n248463),
	.d(n248462));
   no04f04 U265074 (.o(n248467),
	.a(n248445),
	.b(n248444),
	.c(n248443),
	.d(FE_OFN581_n248442));
   na04f03 U265075 (.o(n248464),
	.a(n248453),
	.b(n248452),
	.c(n248451),
	.d(n248450));
   no04f01 U265076 (.o(n248075),
	.a(n248053),
	.b(n248052),
	.c(n248051),
	.d(n248050));
   no04f02 U265077 (.o(n248074),
	.a(n248073),
	.b(n248072),
	.c(n248071),
	.d(n248070));
   na04f03 U265078 (.o(n248052),
	.a(n248041),
	.b(n248040),
	.c(n248039),
	.d(n248038));
   no04f06 U265079 (.o(n248116),
	.a(FE_OFN234_n248115),
	.b(n248114),
	.c(n248113),
	.d(n248112));
   no04f01 U265080 (.o(n248117),
	.a(n248095),
	.b(n248094),
	.c(n248093),
	.d(n248092));
   na04f06 U265081 (.o(n248113),
	.a(n248107),
	.b(n248106),
	.c(n248105),
	.d(n248104));
   no04f02 U265082 (.o(n248719),
	.a(n248697),
	.b(n248696),
	.c(n248695),
	.d(n248694));
   no04f08 U265083 (.o(n248718),
	.a(n248717),
	.b(n248716),
	.c(n248715),
	.d(n248714));
   na04f04 U265084 (.o(n248696),
	.a(n248685),
	.b(n248684),
	.c(n248683),
	.d(n248682));
   no04f02 U265085 (.o(n248760),
	.a(n248759),
	.b(n248758),
	.c(n248757),
	.d(n248756));
   no04f01 U265086 (.o(n248761),
	.a(n248739),
	.b(n248738),
	.c(n248737),
	.d(n248736));
   na04f02 U265087 (.o(n248756),
	.a(n248755),
	.b(n248754),
	.c(n248753),
	.d(n248752));
   no04f01 U265088 (.o(n248354),
	.a(n248332),
	.b(n248331),
	.c(n248330),
	.d(n248329));
   no04f06 U265089 (.o(n248353),
	.a(FE_OFN376_n248352),
	.b(n248351),
	.c(n248350),
	.d(n248349));
   na04f03 U265090 (.o(n248332),
	.a(n248316),
	.b(n248315),
	.c(n248314),
	.d(n248313));
   no04f01 U265091 (.o(n248803),
	.a(n248781),
	.b(n248780),
	.c(n248779),
	.d(n248778));
   na04s02 U265092 (.o(n248780),
	.a(n248769),
	.b(n248768),
	.c(n248767),
	.d(n248766));
   na02s01 U265093 (.o(regtop_w1_hdi00_q[5]),
	.a(FE_OFN384_n248677),
	.b(n248676));
   no04f03 U265094 (.o(n248677),
	.a(n248655),
	.b(n248654),
	.c(n248653),
	.d(n248652));
   na04f04 U265095 (.o(n248654),
	.a(n248643),
	.b(n248642),
	.c(n248641),
	.d(n248640));
   no04f03 U265096 (.o(n248593),
	.a(n248571),
	.b(n248570),
	.c(n248569),
	.d(n248568));
   na04f03 U265097 (.o(n248570),
	.a(n248559),
	.b(n248558),
	.c(n248557),
	.d(n248556));
   no04f02 U265098 (.o(n248551),
	.a(n248529),
	.b(n248528),
	.c(FE_OFN248_n248527),
	.d(n248526));
   na04f02 U265099 (.o(n248527),
	.a(n248521),
	.b(n248520),
	.c(n248519),
	.d(n248518));
   no04f04 U265100 (.o(n248033),
	.a(n248011),
	.b(n248010),
	.c(n248009),
	.d(n248008));
   na04f02 U265101 (.o(n248010),
	.a(n247999),
	.b(n247998),
	.c(n247997),
	.d(n247996));
   no04f04 U265102 (.o(n248635),
	.a(n248613),
	.b(n248612),
	.c(n248611),
	.d(n248610));
   na04f06 U265103 (.o(n248610),
	.a(n248609),
	.b(n248608),
	.c(n248607),
	.d(n248606));
   no04f04 U265104 (.o(n248228),
	.a(n248206),
	.b(n248205),
	.c(n248204),
	.d(n248203));
   na02f01 U265105 (.o(busrtop_b_rreq_N104),
	.a(n245611),
	.b(n245610));
   no02f01 U265106 (.o(busrtop_b_rreq_N103),
	.a(n245618),
	.b(n245617));
   no02f01 U265107 (.o(n245617),
	.a(n245616),
	.b(n245615));
   na02f01 U265108 (.o(busrtop_b_rreq_N102),
	.a(n245626),
	.b(n245625));
   na02f01 U265109 (.o(n245625),
	.a(n245624),
	.b(n245623));
   no02f01 U265110 (.o(busrtop_b_rreq_N101),
	.a(n245633),
	.b(n245632));
   no02f01 U265111 (.o(n245632),
	.a(n245631),
	.b(n245630));
   no02s01 U265112 (.o(n245647),
	.a(n245646),
	.b(n245645));
   no02s01 U265113 (.o(n245674),
	.a(n245670),
	.b(n245671));
   no02f08 U265114 (.o(n249639),
	.a(n246372),
	.b(n245470));
   no02f06 U265115 (.o(n249787),
	.a(n246372),
	.b(n245461));
   in01s01 U265117 (.o(n246805),
	.a(n246365));
   in01f01 U265118 (.o(n246128),
	.a(regtop_g_udb2_r[6]));
   na02f04 U265119 (.o(n246068),
	.a(regtop_g_udb2_r[2]),
	.b(n246076));
   na02f03 U265120 (.o(n246077),
	.a(n246070),
	.b(regtop_g_udb0_r[2]));
   in01s01 U265121 (.o(n245875),
	.a(n245895));
   na02s01 U265122 (.o(n245582),
	.a(n252517),
	.b(regtop_g_paramadr_r[2]));
   ao22f01 U265123 (.o(n245971),
	.a(vldtop_vld_syndec_UREG[23]),
	.b(vldtop_vld_syndec_ADP[1]),
	.c(vldtop_vld_syndec_UREG[25]),
	.d(n246419));
   in01s01 U265124 (.o(n246038),
	.a(vldtop_vld_syndec_UREG[14]));
   ao22s01 U265125 (.o(n246273),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(vldtop_vld_syndec_vld_vlfeed_lower[13]),
	.c(n246419),
	.d(vldtop_vld_syndec_vld_vlfeed_lower[15]));
   na02s01 U265126 (.o(n245876),
	.a(n245875),
	.b(vh_1_ph_add[8]));
   no02s01 U265127 (.o(n252247),
	.a(regtop_g_paramadr_r[1]),
	.b(n252255));
   in01s01 U265128 (.o(n246657),
	.a(n246656));
   na02s01 U265129 (.o(n246049),
	.a(n246419),
	.b(n246048));
   na02s01 U265130 (.o(n246499),
	.a(n246568),
	.b(n246571));
   ao22s01 U265131 (.o(n246381),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n247368),
	.c(n246419),
	.d(FE_OFN543_vldtop_vld_syndec_vld_vlfeed_lower_26_));
   in01s01 U265132 (.o(n246694),
	.a(n246271));
   in01s01 U265133 (.o(n245987),
	.a(n249319));
   in01s01 U265134 (.o(n245832),
	.a(n245830));
   ao22s01 U265135 (.o(n249719),
	.a(n249718),
	.b(regtop_g_hclr_r_s),
	.c(n252867),
	.d(regtop_g_dcnt_r));
   na02f04 U265136 (.o(n249040),
	.a(n249038),
	.b(n249051));
   in01s01 U265137 (.o(n246544),
	.a(n246543));
   in01s01 U265138 (.o(n246037),
	.a(vldtop_vld_syndec_UREG[22]));
   ao22f01 U265139 (.o(n245974),
	.a(n246653),
	.b(n246337),
	.c(n246658),
	.d(n246285));
   in01s01 U265140 (.o(n246718),
	.a(n246713));
   in01s01 U265141 (.o(n246463),
	.a(n246315));
   in01s01 U265142 (.o(n246394),
	.a(n246663));
   in01s01 U265143 (.o(n246424),
	.a(n246423));
   no02s01 U265147 (.o(n245316),
	.a(g_field_start_add_r[31]),
	.b(n245314));
   no04s01 U265148 (.o(n245993),
	.a(y1_bs_data_r[8]),
	.b(y1_bs_data_r[9]),
	.c(y1_bs_data_r[10]),
	.d(y1_bs_data_r[11]));
   na02s01 U265149 (.o(n245814),
	.a(n245829),
	.b(n245815));
   in01s01 U265150 (.o(n245575),
	.a(n246840));
   no02f08 U265151 (.o(n249637),
	.a(n246372),
	.b(n249697));
   in01s01 U265152 (.o(n247594),
	.a(regtop_g_hclr_r_s));
   no02m02 U265153 (.o(n246105),
	.a(n246101),
	.b(n246102));
   ao22f01 U265154 (.o(n246461),
	.a(n246700),
	.b(n246312),
	.c(n246568),
	.d(n246340));
   in01s01 U265155 (.o(n246664),
	.a(n246711));
   na02s01 U265156 (.o(n246414),
	.a(n246568),
	.b(n246536));
   in01s01 U265159 (.o(n245411),
	.a(n245406));
   in01s01 U265160 (.o(n245374),
	.a(n245364));
   in01f01 U265161 (.o(n245350),
	.a(n245341));
   in01s01 U265162 (.o(n249873),
	.a(busrtop_b_rreq_vrh_add1_r[6]));
   in01s01 U265163 (.o(n249912),
	.a(busrtop_b_rreq_vrh_add1_r[1]));
   na02s01 U265164 (.o(n249689),
	.a(n249733),
	.b(regtop_g_vbsv_r[1]));
   ao22f01 U265165 (.o(n249736),
	.a(n249731),
	.b(g_field_offset_r[0]),
	.c(n249730),
	.d(regtop_g_icsh_r));
   ao22f01 U265166 (.o(n249473),
	.a(FE_OFN392_n249635),
	.b(regtop_g_dvs_r[13]),
	.c(n249634),
	.d(regtop_g_tmc_r[13]));
   ao22f01 U265167 (.o(n249560),
	.a(regtop_g_vd_r[8]),
	.b(FE_OFN264_n249636),
	.c(regtop_g_fcvo2_r[8]),
	.d(n249639));
   ao22f02 U265168 (.o(n249428),
	.a(n249663),
	.b(regtop_g_isfp_r),
	.c(regtop_g_icfp_r),
	.d(n249547));
   ao22s01 U265169 (.o(n249442),
	.a(n249629),
	.b(regtop_g_brv_r[17]),
	.c(n249638),
	.d(regtop_g_cp_r[1]));
   in01s01 U265171 (.o(n249165),
	.a(regtop_g_paramdata_r[9]));
   ao12f01 U265172 (.o(n249130),
	.a(n249126),
	.b(n249127),
	.c(regtop_g_atscd_r[18]));
   in01s01 U265173 (.o(n247036),
	.a(n247039));
   na02s01 U265174 (.o(n245538),
	.a(n245762),
	.b(n245537));
   in01s01 U265175 (.o(n245966),
	.a(regtop_g_atscd_r[9]));
   in01s01 U265176 (.o(n245960),
	.a(regtop_g_atscd_r[8]));
   in01s01 U265177 (.o(n246621),
	.a(regtop_g_usrd_r[17]));
   in01s01 U265178 (.o(n246757),
	.a(regtop_g_usrd_r[29]));
   in01f01 U265179 (.o(n245585),
	.a(n245568));
   in01s01 U265180 (.o(n246977),
	.a(n246976));
   in01s01 U265181 (.o(n247139),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[6]));
   in01s01 U265182 (.o(n247446),
	.a(y1_bs_data[25]));
   in01s01 U265183 (.o(n247442),
	.a(y1_bs_data[11]));
   in01s01 U265184 (.o(n247378),
	.a(y1_bs_data[1]));
   ao22s01 U265185 (.o(n247578),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1052]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[28]));
   ao22s01 U265186 (.o(n247557),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1596]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[572]));
   ao22s01 U265187 (.o(n247534),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1307]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[283]));
   ao22s01 U265188 (.o(n247511),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1851]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[827]));
   ao22s01 U265189 (.o(n247500),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1147]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[123]));
   ao22s01 U265190 (.o(n247097),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1626]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[602]));
   ao22s01 U265191 (.o(n247418),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1881]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[857]));
   ao22s01 U265192 (.o(n248402),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1688]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[664]));
   ao22s01 U265193 (.o(n248459),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1292]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[268]));
   ao22s01 U265194 (.o(n248096),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1866]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[842]));
   ao22s01 U265195 (.o(n248744),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1928]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[904]));
   ao22s01 U265196 (.o(n248343),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1735]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[711]));
   ao22s01 U265197 (.o(n248670),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1541]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[517]));
   ao22s01 U265198 (.o(n248510),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1891]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[867]));
   ao22s01 U265199 (.o(n248598),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1953]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[929]));
   ao22s01 U265200 (.o(n248197),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1760]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[736]));
   in01s01 U265201 (.o(n245400),
	.a(n245642));
   in01s01 U265202 (.o(n245680),
	.a(n245678));
   ao12s01 U265203 (.o(n249887),
	.a(n249885),
	.b(n249893),
	.c(n249886));
   in01s01 U265204 (.o(n246213),
	.a(n246212));
   na02f02 U265205 (.o(n249057),
	.a(n249056),
	.b(n249055));
   ao12s01 U265206 (.o(n252271),
	.a(n252269),
	.b(n252270),
	.c(regtop_g_wd_r[2]));
   in01s01 U265207 (.o(n252570),
	.a(n252571));
   no02s01 U265208 (.o(n245543),
	.a(n245542),
	.b(n245545));
   in01f01 U265209 (.o(n247002),
	.a(n246025));
   oa12f02 U265210 (.o(n247017),
	.a(n246397),
	.b(n246399),
	.c(n246398));
   in01f01 U265211 (.o(n252822),
	.a(n252818));
   in01s01 U265212 (.o(n246690),
	.a(n246836));
   na02s01 U265213 (.o(n247170),
	.a(g_swrst_r_n),
	.b(n247169));
   na03f01 U265214 (.o(n247391),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247494),
	.c(n247390));
   na02s01 U265215 (.o(n249292),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[2]));
   na02f01 U265216 (.o(n249303),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[15]));
   in01s01 U265217 (.o(n245819),
	.a(n245818));
   na02s01 U265218 (.o(n249869),
	.a(n253125),
	.b(vh_1_ph_add[7]));
   na02s01 U265219 (.o(n249918),
	.a(n253125),
	.b(vh_1_ph_add[1]));
   no02s01 U265220 (.o(n249288),
	.a(busrtop_b_rreq_vrh_add1_r[0]),
	.b(n249287));
   ao22s01 U265221 (.o(n249683),
	.a(g_fcyc_r[2]),
	.b(n249841),
	.c(n249713),
	.d(regtop_g_nfst_r[2]));
   na02f03 U265222 (.o(n249478),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[13]));
   ao22s01 U265223 (.o(n249454),
	.a(FE_OFN546_n245460),
	.b(regtop_g_brv_r[15]),
	.c(FE_OFN552_n245462),
	.d(regtop_g_vd_r[15]));
   in01s01 U265224 (.o(n249797),
	.a(n249796));
   na02f02 U265225 (.o(n249446),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[17]));
   oa22s01 U265226 (.o(n250007),
	.a(n250018),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[457]),
	.d(FE_OFN402_n249999));
   oa22s01 U265227 (.o(n250041),
	.a(n250053),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[427]),
	.d(FE_OFN270_n250035));
   oa22s01 U265228 (.o(n250075),
	.a(n250089),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[397]),
	.d(n250071));
   oa22s01 U265229 (.o(n250093),
	.a(n250126),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[382]),
	.d(FE_OFN193_n250107));
   oa22s01 U265230 (.o(n250296),
	.a(n250307),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[202]),
	.d(FE_OFN408_n250289));
   oa22s01 U265231 (.o(n250329),
	.a(n250343),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[172]),
	.d(FE_OFN280_n250324));
   oa22s01 U265232 (.o(n250347),
	.a(n250378),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[157]),
	.d(FE_OFN410_n250360));
   oa22s01 U265233 (.o(n250380),
	.a(n250413),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[127]),
	.d(FE_OFN195_n250395));
   oa22s01 U265234 (.o(n250545),
	.a(n250556),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1001]),
	.d(FE_OFN288_n250540));
   oa22s01 U265235 (.o(n250579),
	.a(n250591),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[971]),
	.d(FE_OFN412_n250576));
   oa22s01 U265236 (.o(n250596),
	.a(n250626),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[956]),
	.d(FE_OFN290_n250611));
   oa22s01 U265237 (.o(n250629),
	.a(n250662),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[926]),
	.d(FE_OFN414_n250646));
   oa22s01 U265238 (.o(n250828),
	.a(n250839),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[746]),
	.d(n250824));
   oa22s01 U265239 (.o(n250861),
	.a(n250875),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[716]),
	.d(FE_OFN416_n250859));
   oa22s01 U265240 (.o(n250879),
	.a(n250910),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[701]),
	.d(FE_OFN300_n250895));
   oa22s01 U265241 (.o(n250912),
	.a(n250945),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[671]),
	.d(FE_OFN418_n250930));
   oa22s01 U265242 (.o(n251077),
	.a(n251088),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[521]),
	.d(FE_OFN306_n251072));
   oa22s01 U265243 (.o(n251111),
	.a(n251123),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1515]),
	.d(FE_OFN309_n251105));
   oa22s01 U265244 (.o(n251144),
	.a(n251158),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1485]),
	.d(FE_OFN420_n251140));
   oa22s01 U265245 (.o(n251161),
	.a(n251194),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1470]),
	.d(FE_OFN311_n251175));
   oa22s01 U265246 (.o(n251360),
	.a(n251371),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1290]),
	.d(FE_OFN318_n251353));
   oa22s01 U265247 (.o(n251393),
	.a(n251407),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1260]),
	.d(FE_OFN320_n251388));
   oa22s01 U265248 (.o(n251411),
	.a(n251442),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1245]),
	.d(FE_OFN426_n251424));
   oa22s01 U265249 (.o(n251444),
	.a(n251477),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1215]),
	.d(FE_OFN322_n251459));
   oa22s01 U265250 (.o(n251608),
	.a(n251619),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1065]),
	.d(FE_OFN327_n251600));
   oa22s01 U265251 (.o(n251643),
	.a(n251655),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1035]),
	.d(FE_OFN329_n251637));
   oa22s01 U265252 (.o(n251660),
	.a(n251690),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[2044]),
	.d(FE_OFN331_n251675));
   oa22s01 U265253 (.o(n251693),
	.a(n251726),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[2014]),
	.d(FE_OFN430_n251710));
   oa22s01 U265254 (.o(n251891),
	.a(n251902),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1834]),
	.d(FE_OFN337_n251887));
   oa22s01 U265255 (.o(n251925),
	.a(n251939),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1804]),
	.d(FE_OFN339_n251923));
   oa22s01 U265256 (.o(n251944),
	.a(n251975),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1789]),
	.d(FE_OFN341_n251960));
   oa22s01 U265257 (.o(n251978),
	.a(n252011),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1759]),
	.d(FE_OFN434_n251996));
   oa22s01 U265258 (.o(n252146),
	.a(n252157),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1609]),
	.d(FE_OFN345_n252141));
   oa22s01 U265259 (.o(n252181),
	.a(n252193),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1579]),
	.d(FE_OFN348_n252178));
   oa22s01 U265260 (.o(n252200),
	.a(n252230),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1564]),
	.d(FE_OFN350_n252215));
   na02s01 U265261 (.o(n249352),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[30]));
   na02s01 U265262 (.o(n249337),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[15]));
   na02s01 U265263 (.o(n249322),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[0]));
   ao12f01 U265264 (.o(n248988),
	.a(n248987),
	.b(n248991),
	.c(n249073));
   in01s01 U265265 (.o(n252297),
	.a(regtop_g_fbst_r[5]));
   in01s01 U265266 (.o(n246948),
	.a(regtop_g_udb0_r[0]));
   in01s01 U265268 (.o(n252558),
	.a(regtop_g_dhs_r[11]));
   in01s01 U265269 (.o(n252579),
	.a(regtop_g_adb_r[6]));
   in01s01 U265270 (.o(n252649),
	.a(regtop_g_dvs_r[4]));
   in01f04 U265271 (.o(n252664),
	.a(regtop_g_paramdata_r[21]));
   in01s01 U265272 (.o(n252789),
	.a(n252787));
   in01s01 U265274 (.o(n246748),
	.a(n246746));
   na02s01 U265275 (.o(n246584),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247009));
   na02s01 U265276 (.o(n246218),
	.a(n246964),
	.b(vldtop_vld_syndec_vld_seqhed_state_0_));
   na02s01 U265277 (.o(n246220),
	.a(vldtop_vld_syndec_vld_vscdet_v_detvald_r[1]),
	.b(n246779));
   in01s01 U265278 (.o(n252854),
	.a(g_vsdc_r[3]));
   oa12s01 U265279 (.o(n246208),
	.a(g_swrst_r_n),
	.b(vldtop_vld_syndec_vld_vlfeed_feed_on),
	.c(g_init_vld_r_s));
   in01s01 U265280 (.o(n252881),
	.a(g_mbc_r[9]));
   in01s01 U265281 (.o(n252895),
	.a(g_pcut_r[3]));
   in01s01 U265282 (.o(n252909),
	.a(regtop_g_wd_r[27]));
   in01s01 U265283 (.o(n252924),
	.a(regtop_g_wd_r[12]));
   in01s01 U265284 (.o(n252955),
	.a(g_vldmode_r[0]));
   oa22s01 U265285 (.o(n253004),
	.a(n253012),
	.b(regtop_g_wd_r[5]),
	.c(g_field_offset_r[5]),
	.d(n253011));
   in01s01 U265286 (.o(n253022),
	.a(g_cbcr_offset_r[7]));
   in01f02 U265287 (.o(n249313),
	.a(busiftop_vmem_ren_g));
   in01s01 U265288 (.o(n253122),
	.a(n249292));
   in01s01 U265289 (.o(n253109),
	.a(n249305));
   oa12s01 U265290 (.o(busiftop_N58),
	.a(n249293),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   oa12f01 U265291 (.o(busiftop_N41),
	.a(n246210),
	.b(busiftop_vmem_ch_r),
	.c(n245865));
   no02s01 U265292 (.o(busrtop_b_rreq_N428),
	.a(n249279),
	.b(n249278));
   oa12f02 U265293 (.o(n244981),
	.a(n249407),
	.b(n245444),
	.c(n249408));
   in01s01 U265294 (.o(n184635),
	.a(n249954));
   in01s01 U265295 (.o(n184650),
	.a(n249970));
   in01s01 U265296 (.o(n184665),
	.a(n249987));
   in01s01 U265297 (.o(n184680),
	.a(n250003));
   in01s01 U265298 (.o(n184695),
	.a(n250021));
   in01s01 U265299 (.o(n184710),
	.a(n250037));
   in01s01 U265300 (.o(n184725),
	.a(n250054));
   in01s01 U265301 (.o(n184740),
	.a(n250070));
   in01s01 U265302 (.o(n184755),
	.a(n250087));
   in01s01 U265303 (.o(n184770),
	.a(n250104));
   in01s01 U265304 (.o(n184785),
	.a(n250121));
   in01s01 U265305 (.o(n184800),
	.a(n250139));
   in01s01 U265306 (.o(n184815),
	.a(n250156));
   in01s01 U265307 (.o(n184830),
	.a(n250173));
   in01s01 U265308 (.o(n184845),
	.a(n250189));
   in01s01 U265309 (.o(n184860),
	.a(n250209));
   in01s01 U265310 (.o(n184875),
	.a(n250225));
   in01s01 U265311 (.o(n184890),
	.a(n250243));
   in01s01 U265312 (.o(n184905),
	.a(n250259));
   in01s01 U265313 (.o(n184920),
	.a(n250276));
   in01s01 U265314 (.o(n184935),
	.a(n250292));
   in01s01 U265315 (.o(n184950),
	.a(n250309));
   in01s01 U265316 (.o(n184965),
	.a(n250325));
   in01s01 U265317 (.o(n184980),
	.a(n250341));
   in01s01 U265318 (.o(n184995),
	.a(n250358));
   in01s01 U265319 (.o(n185010),
	.a(n250375));
   in01s01 U265320 (.o(n185025),
	.a(n250391));
   in01s01 U265321 (.o(n185040),
	.a(n250408));
   in01s01 U265322 (.o(n185055),
	.a(n250424));
   in01s01 U265323 (.o(n185070),
	.a(n250440));
   in01s01 U265324 (.o(n185085),
	.a(n250458));
   in01s01 U265325 (.o(n185100),
	.a(n250474));
   in01s01 U265326 (.o(n185115),
	.a(n250492));
   in01s01 U265327 (.o(n185130),
	.a(n250508));
   in01s01 U265328 (.o(n185145),
	.a(n250525));
   in01s01 U265329 (.o(n185160),
	.a(n250541));
   in01s01 U265330 (.o(n185175),
	.a(n250559));
   in01s01 U265331 (.o(n185190),
	.a(n250574));
   in01s01 U265332 (.o(n185205),
	.a(n250592));
   in01s01 U265333 (.o(n185220),
	.a(n250607));
   in01s01 U265334 (.o(n185235),
	.a(n250624));
   in01s01 U265335 (.o(n185250),
	.a(n250640));
   in01s01 U265336 (.o(n185265),
	.a(n250657));
   in01s01 U265337 (.o(n185280),
	.a(n250674));
   in01s01 U265338 (.o(n185295),
	.a(n250691));
   in01s01 U265339 (.o(n185310),
	.a(n250707));
   in01s01 U265340 (.o(n185325),
	.a(n250723));
   in01s01 U265341 (.o(n185340),
	.a(n250740));
   in01s01 U265342 (.o(n185355),
	.a(n250756));
   in01s01 U265343 (.o(n185370),
	.a(n250775));
   in01s01 U265344 (.o(n185385),
	.a(n250791));
   in01s01 U265345 (.o(n185400),
	.a(n250808));
   in01s01 U265346 (.o(n185415),
	.a(n250823));
   in01s01 U265347 (.o(n185430),
	.a(n250841));
   in01s01 U265348 (.o(n185445),
	.a(n250856));
   in01s01 U265349 (.o(n185460),
	.a(n250873));
   in01s01 U265350 (.o(n185475),
	.a(n250890));
   in01s01 U265351 (.o(n185490),
	.a(n250907));
   in01s01 U265352 (.o(n185505),
	.a(n250923));
   in01s01 U265353 (.o(n185520),
	.a(n250940));
   in01s01 U265354 (.o(n185535),
	.a(n250956));
   in01s01 U265355 (.o(n185550),
	.a(n250972));
   in01s01 U265356 (.o(n185565),
	.a(n250990));
   in01s01 U265357 (.o(n185580),
	.a(n251006));
   in01s01 U265358 (.o(n185595),
	.a(n251023));
   in01s01 U265359 (.o(n185610),
	.a(n251039));
   in01s01 U265360 (.o(n185625),
	.a(n251057));
   in01s01 U265361 (.o(n185640),
	.a(n251073));
   in01s01 U265362 (.o(n185655),
	.a(n251091));
   in01s01 U265363 (.o(n185670),
	.a(n251107));
   in01s01 U265364 (.o(n185685),
	.a(n251124));
   in01s01 U265365 (.o(n185700),
	.a(n251139));
   in01s01 U265366 (.o(n185715),
	.a(n251156));
   in01s01 U265367 (.o(n185730),
	.a(n251172));
   in01s01 U265368 (.o(n185745),
	.a(n251189));
   in01s01 U265369 (.o(n185760),
	.a(n251206));
   in01s01 U265370 (.o(n185775),
	.a(n251223));
   in01s01 U265371 (.o(n185790),
	.a(n251239));
   in01s01 U265372 (.o(n185805),
	.a(n251255));
   in01s01 U265373 (.o(n185820),
	.a(n251272));
   in01s01 U265374 (.o(n185835),
	.a(n251288));
   in01s01 U265375 (.o(n185850),
	.a(n251306));
   in01s01 U265376 (.o(n185865),
	.a(n251322));
   in01s01 U265377 (.o(n185880),
	.a(n251340));
   in01s01 U265378 (.o(n185895),
	.a(n251356));
   in01s01 U265379 (.o(n185910),
	.a(n251373));
   in01s01 U265380 (.o(n185925),
	.a(n251389));
   in01s01 U265381 (.o(n185940),
	.a(n251405));
   in01s01 U265382 (.o(n185955),
	.a(n251422));
   in01s01 U265383 (.o(n185970),
	.a(n251439));
   in01s01 U265384 (.o(n185985),
	.a(n251455));
   in01s01 U265385 (.o(n186000),
	.a(n251472));
   in01s01 U265386 (.o(n186015),
	.a(n251488));
   in01s01 U265387 (.o(n186030),
	.a(n251504));
   in01s01 U265388 (.o(n186045),
	.a(n251522));
   in01s01 U265389 (.o(n186060),
	.a(n251538));
   in01s01 U265390 (.o(n186075),
	.a(n251555));
   in01s01 U265391 (.o(n186090),
	.a(n251571));
   in01s01 U265392 (.o(n186105),
	.a(n251588));
   in01s01 U265393 (.o(n186120),
	.a(n251604));
   in01s01 U265394 (.o(n186135),
	.a(n251623));
   in01s01 U265395 (.o(n186150),
	.a(n251639));
   in01s01 U265396 (.o(n186165),
	.a(n251656));
   in01s01 U265397 (.o(n186180),
	.a(n251671));
   in01s01 U265398 (.o(n186195),
	.a(n251688));
   in01s01 U265399 (.o(n186210),
	.a(n251704));
   in01s01 U265400 (.o(n186225),
	.a(n251721));
   in01s01 U265401 (.o(n186240),
	.a(n251738));
   in01s01 U265402 (.o(n186255),
	.a(n251755));
   in01s01 U265403 (.o(n186270),
	.a(n251771));
   in01s01 U265404 (.o(n186285),
	.a(n251787));
   in01s01 U265405 (.o(n186300),
	.a(n251804));
   in01s01 U265406 (.o(n186315),
	.a(n251820));
   in01s01 U265407 (.o(n186330),
	.a(n251838));
   in01s01 U265408 (.o(n186345),
	.a(n251854));
   in01s01 U265409 (.o(n186360),
	.a(n251871));
   in01s01 U265410 (.o(n186375),
	.a(n251886));
   in01s01 U265411 (.o(n186390),
	.a(n251905));
   in01s01 U265412 (.o(n186405),
	.a(n251920));
   in01s01 U265413 (.o(n186420),
	.a(n251937));
   in01s01 U265414 (.o(n186435),
	.a(n251955));
   in01s01 U265415 (.o(n186450),
	.a(n251972));
   in01s01 U265416 (.o(n186465),
	.a(n251989));
   in01s01 U265417 (.o(n186480),
	.a(n252006));
   in01s01 U265418 (.o(n186495),
	.a(n252023));
   in01s01 U265419 (.o(n186510),
	.a(n252039));
   in01s01 U265420 (.o(n186525),
	.a(n252058));
   in01s01 U265421 (.o(n186540),
	.a(n252074));
   in01s01 U265422 (.o(n186555),
	.a(n252092));
   in01s01 U265423 (.o(n186570),
	.a(n252108));
   in01s01 U265424 (.o(n186585),
	.a(n252126));
   in01s01 U265425 (.o(n186600),
	.a(n252142));
   in01s01 U265426 (.o(n186615),
	.a(n252161));
   in01s01 U265427 (.o(n186630),
	.a(n252176));
   in01s01 U265428 (.o(n186645),
	.a(n252194));
   in01s01 U265429 (.o(n186660),
	.a(n252211));
   in01s01 U265430 (.o(n186675),
	.a(n252228));
   in01s01 U265431 (.o(regtop_N2012),
	.a(n249341));
   in01s01 U265432 (.o(regtop_N1997),
	.a(n249326));
   na02f01 U265433 (.o(n245012),
	.a(n249134),
	.b(n249133));
   in01s01 U265434 (.o(n186692),
	.a(n247596));
   in01s01 U265435 (.o(n186720),
	.a(n246866));
   in01s01 U265436 (.o(n211880),
	.a(n252318));
   in01s01 U265437 (.o(n211895),
	.a(n252333));
   in01s01 U265438 (.o(n211910),
	.a(n252354));
   in01s01 U265439 (.o(n211925),
	.a(n246602));
   in01s01 U265440 (.o(n211940),
	.a(n246587));
   oa12s01 U265441 (.o(n211962),
	.a(n252366),
	.b(n252818),
	.c(n252367));
   in01s01 U265442 (.o(n211977),
	.a(n252393));
   in01s01 U265443 (.o(n211992),
	.a(n252413));
   in01s01 U265444 (.o(n212007),
	.a(n252432));
   in01s01 U265445 (.o(n212022),
	.a(n252451));
   in01s01 U265446 (.o(n212037),
	.a(n252471));
   in01s01 U265447 (.o(n212067),
	.a(n252500));
   in01s01 U265448 (.o(n212082),
	.a(n252526));
   ao22s01 U265449 (.o(n212127),
	.a(n252563),
	.b(n252656),
	.c(n252553),
	.d(n252561));
   na02s01 U265450 (.o(n212142),
	.a(n246257),
	.b(n246256));
   in01s01 U265451 (.o(n212172),
	.a(n252627));
   ao22s01 U265452 (.o(n212187),
	.a(n252671),
	.b(n252650),
	.c(n252649),
	.d(FE_OFN43_n252668));
   in01s01 U265453 (.o(n212202),
	.a(n252688));
   in01s01 U265454 (.o(n212217),
	.a(n252712));
   in01s01 U265455 (.o(n212232),
	.a(n252729));
   in01s01 U265456 (.o(n212247),
	.a(n252746));
   oa12s01 U265457 (.o(n212262),
	.a(n252777),
	.b(n252778),
	.c(n252780));
   na02s01 U265458 (.o(n212277),
	.a(n246636),
	.b(n246635));
   in01s01 U265459 (.o(vldtop_vld_syndec_vld_outbuf_N484),
	.a(n246336));
   in01s01 U265460 (.o(vldtop_vld_syndec_vld_outbuf_N469),
	.a(n246475));
   oa12f01 U265461 (.o(n212423),
	.a(n247254),
	.b(n249028),
	.c(n247255));
   ao22s01 U265462 (.o(n212537),
	.a(FE_OFN454_n252863),
	.b(n252983),
	.c(n252838),
	.d(n252834));
   na02f01 U265463 (.o(n212592),
	.a(n247373),
	.b(n247372));
   ao12f01 U265464 (.o(n253084),
	.a(n247274),
	.b(n247275),
	.c(FE_OCPN583_n247126));
   na02f01 U265465 (.o(n212622),
	.a(n247263),
	.b(n247262));
   ao12f01 U265466 (.o(n253099),
	.a(n247384),
	.b(n247385),
	.c(n247126));
   na02s01 U265467 (.o(n212681),
	.a(n252873),
	.b(n252872));
   ao22s01 U265468 (.o(n212694),
	.a(n252875),
	.b(n252918),
	.c(n252891),
	.d(FE_OFN441_n252905));
   in01s01 U265469 (.o(n212739),
	.a(n252967));
   in01s01 U265470 (.o(n212754),
	.a(n252986));
   in01s01 U265471 (.o(n212769),
	.a(n253005));
   in01s01 U265472 (.o(n212784),
	.a(n253025));
   no02s01 U265473 (.o(busrtop_b_rreq_N97),
	.a(n245663),
	.b(n245662));
   na02f01 U265474 (.o(vmem_ren),
	.a(vmem_wen),
	.b(n249313));
   ao12f08 U265475 (.o(n249511),
	.a(n249548),
	.b(n252972),
	.c(g_field_start_add_r[10]));
   no02s01 U265491 (.o(n245430),
	.a(g_field_start_add_r[30]),
	.b(busrtop_b_rreq_vrh_rrq_fldstatadd_r[30]));
   in01s01 U265492 (.o(n245319),
	.a(n245430));
   no02s01 U265493 (.o(n245314),
	.a(g_field_start_add_r[31]),
	.b(busrtop_b_rreq_vrh_rrq_fldstatadd_r[31]));
   no02s01 U265494 (.o(n245315),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[31]),
	.b(n245314));
   no02s01 U265495 (.o(n245318),
	.a(n245316),
	.b(n245315));
   no02s01 U265496 (.o(n245317),
	.a(n245319),
	.b(n245318));
   in01s01 U265497 (.o(n245321),
	.a(n245317));
   na02s01 U265498 (.o(n245320),
	.a(n245319),
	.b(n245318));
   na02s01 U265499 (.o(n245438),
	.a(n245321),
	.b(n245320));
   in01f01 U265500 (.o(n245329),
	.a(n245324));
   in01s01 U265501 (.o(n245327),
	.a(g_field_start_add_r[11]));
   no02f01 U265502 (.o(n245751),
	.a(n245327),
	.b(busrtop_b_rreq_N296));
   no02f02 U265503 (.o(n245758),
	.a(busrtop_b_rreq_N295),
	.b(g_field_start_add_r[10]));
   na02f01 U265504 (.o(n245752),
	.a(n245327),
	.b(busrtop_b_rreq_N296));
   oa12f04 U265505 (.o(n245734),
	.a(n245752),
	.b(n245751),
	.c(n245758));
   oa12m02 U265506 (.o(n245331),
	.a(n245736),
	.b(n245735),
	.c(n245744));
   in01f01 U265507 (.o(n245347),
	.a(n245336));
   in01f01 U265508 (.o(n245346),
	.a(n245335));
   in01f01 U265509 (.o(n245351),
	.a(n245342));
   oa12f01 U265510 (.o(n245665),
	.a(n245713),
	.b(n245712),
	.c(n245727));
   no02f01 U265512 (.o(n245358),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[19]),
	.b(n245364));
   no02f01 U265513 (.o(n245357),
	.a(g_field_start_add_r[19]),
	.b(n245364));
   in01f01 U265514 (.o(n245369),
	.a(n245361));
   in01s01 U265515 (.o(n245368),
	.a(n245360));
   in01f01 U265516 (.o(n245721),
	.a(n245686));
   no02s01 U265517 (.o(n245366),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[20]),
	.b(n245379));
   no02s01 U265518 (.o(n245365),
	.a(g_field_start_add_r[20]),
	.b(n245379));
   no02f01 U265519 (.o(n245373),
	.a(n245366),
	.b(n245365));
   no02f01 U265520 (.o(n245678),
	.a(n245374),
	.b(n245373));
   na02f01 U265521 (.o(n245687),
	.a(n245370),
	.b(n245369));
   in01f01 U265522 (.o(n245371),
	.a(n245687));
   na02s01 U265523 (.o(n245679),
	.a(n245374),
	.b(n245373));
   no02s01 U265525 (.o(n245378),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[21]),
	.b(n245382));
   in01s01 U265526 (.o(n245380),
	.a(n245379));
   in01s01 U265528 (.o(n245387),
	.a(n245382));
   no02s01 U265529 (.o(n245384),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[22]),
	.b(n245391));
   no02s01 U265530 (.o(n245383),
	.a(g_field_start_add_r[22]),
	.b(n245391));
   in01s01 U265531 (.o(n245388),
	.a(n245657));
   no02s01 U265533 (.o(n245390),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[23]),
	.b(n245394));
   no02s01 U265534 (.o(n245389),
	.a(g_field_start_add_r[23]),
	.b(n245394));
   in01s01 U265535 (.o(n245392),
	.a(n245391));
   in01s01 U265537 (.o(n245399),
	.a(n245394));
   no02s01 U265538 (.o(n245396),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[24]),
	.b(n245403));
   no02s01 U265539 (.o(n245395),
	.a(g_field_start_add_r[24]),
	.b(n245403));
   in01s01 U265541 (.o(n245404),
	.a(n245403));
   no02s01 U265543 (.o(n245407),
	.a(g_field_start_add_r[26]),
	.b(n245413));
   in01f04 U265544 (.o(n245628),
	.a(n245409));
   in01s01 U265545 (.o(n245412),
	.a(n245627));
   in01s01 U265547 (.o(n245417),
	.a(n245413));
   no02s01 U265548 (.o(n245415),
	.a(g_field_start_add_r[27]),
	.b(n245420));
   no02s01 U265549 (.o(n245414),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[27]),
	.b(n245420));
   no02s01 U265551 (.o(n245419),
	.a(g_field_start_add_r[28]),
	.b(n245427));
   no02s01 U265552 (.o(n245418),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[28]),
	.b(n245427));
   in01f01 U265553 (.o(n245422),
	.a(n245420));
   in01s01 U265554 (.o(n245613),
	.a(n245421));
   in01s01 U265555 (.o(n245424),
	.a(n245612));
   no02s01 U265556 (.o(n245426),
	.a(g_field_start_add_r[29]),
	.b(n245433));
   no02s01 U265557 (.o(n245425),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[29]),
	.b(n245433));
   in01s01 U265558 (.o(n245428),
	.a(n245427));
   no02s01 U265559 (.o(n245432),
	.a(g_field_start_add_r[30]),
	.b(n245430));
   no02s01 U265560 (.o(n245431),
	.a(busrtop_b_rreq_vrh_rrq_fldstatadd_r[30]),
	.b(n245430));
   no02s01 U265561 (.o(n245436),
	.a(n245432),
	.b(n245431));
   in01s01 U265562 (.o(n245435),
	.a(n245433));
   no02s01 U265563 (.o(n245434),
	.a(n245436),
	.b(n245435));
   in01s01 U265564 (.o(n245598),
	.a(n245434));
   na02s01 U265565 (.o(n245597),
	.a(n245436),
	.b(n245435));
   in01s01 U265566 (.o(n245437),
	.a(n245597));
   ao12f04 U265567 (.o(n245439),
	.a(n245437),
	.b(n245599),
	.c(n245598));
   no02f01 U265568 (.o(n245442),
	.a(n245438),
	.b(n245439));
   na02f02 U265569 (.o(n245440),
	.a(n245439),
	.b(n245438));
   in01f02 U265570 (.o(n245441),
	.a(n245440));
   no02f01 U265571 (.o(busrtop_b_rreq_N106),
	.a(n245442),
	.b(n245441));
   ao12f01 U265572 (.o(n245486),
	.a(n249825),
	.b(FE_OFN489_n249763),
	.c(regtop_g_fcho0_r[0]));
   in01f02 U265573 (.o(n249547),
	.a(n252958));
   no02f02 U265574 (.o(n249721),
	.a(n245481),
	.b(n245452));
   ao22s01 U265575 (.o(n245476),
	.a(regtop_g_icnf_r),
	.b(n249547),
	.c(regtop_g_mpeg_r),
	.d(n249721));
   na02f03 U265577 (.o(n249375),
	.a(FE_OFN4_n245443),
	.b(n249637));
   in01f06 U265578 (.o(n249838),
	.a(n249375));
   ao22f01 U265579 (.o(n245475),
	.a(regtop_g_hsv_r[0]),
	.b(n249823),
	.c(regtop_g_fcho1_r[0]),
	.d(n249838));
   no02f03 U265580 (.o(n249768),
	.a(n246372),
	.b(n252286));
   ao22f01 U265581 (.o(n245456),
	.a(n249768),
	.b(regtop_g_tff_r),
	.c(n252972),
	.d(g_field_start_add_r[16]));
   ao22s01 U265582 (.o(n245455),
	.a(n249663),
	.b(regtop_g_isnf_r),
	.c(n252944),
	.d(g_pmod_r));
   in01s01 U265583 (.o(n245450),
	.a(n245480));
   ao22f01 U265584 (.o(n245454),
	.a(n249769),
	.b(regtop_g_cf_r[0]),
	.c(FE_OFN266_n249787),
	.d(regtop_g_sc_r));
   na02f06 U265585 (.o(n245453),
	.a(g_pcut_r[0]),
	.b(n249811));
   na04s02 U265586 (.o(n245469),
	.a(n245456),
	.b(n245455),
	.c(n245454),
	.d(n245453));
   no02f04 U265587 (.o(n249630),
	.a(n245491),
	.b(n249697));
   no03f10 U265588 (.o(n249584),
	.a(FE_OFN491_regtop_g_a_r_3_),
	.b(FE_OFN519_regtop_g_a_r_6_),
	.c(n245457));
   ao22f02 U265589 (.o(n245467),
	.a(n249630),
	.b(regtop_g_cpf_r),
	.c(n249584),
	.d(regtop_g_nfst_r[16]));
   ao12s01 U265590 (.o(n245466),
	.a(n249542),
	.b(g_fcyc_r[16]),
	.c(n252912));
   na02f01 U265591 (.o(n245462),
	.a(FE_OFN4_n245443),
	.b(FE_OFN264_n249636));
   in01f04 U265593 (.o(n249813),
	.a(n245463));
   na04f02 U265594 (.o(n245468),
	.a(n245467),
	.b(n245466),
	.c(n245465),
	.d(n245464));
   no02f01 U265595 (.o(n245474),
	.a(n245469),
	.b(n245468));
   na02f01 U265596 (.o(n245472),
	.a(FE_OFN4_n245443),
	.b(FE_OFN392_n249635));
   na02s01 U265597 (.o(n245473),
	.a(regtop_g_dhs_r[0]),
	.b(n249824));
   in01f01 U265599 (.o(n249718),
	.a(n252286));
   na02f02 U265600 (.o(n249396),
	.a(n245479),
	.b(n249718));
   ao12s01 U265602 (.o(n245484),
	.a(n249664),
	.b(n249812),
	.c(regtop_g_tmc_r[16]));
   na02f03 U265603 (.o(n245483),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[16]));
   ao22s01 U265604 (.o(n245513),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[4]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcvo0_r[4]));
   ao22s01 U265605 (.o(n245508),
	.a(n253014),
	.b(g_cbcr_offset_r[4]),
	.c(n249769),
	.d(regtop_g_pali_r[4]));
   na02f01 U265606 (.o(n245507),
	.a(n249630),
	.b(regtop_g_vbsv_r[4]));
   na02f01 U265607 (.o(n245498),
	.a(regtop_g_a_r[6]),
	.b(n245488));
   no02f04 U265608 (.o(n249652),
	.a(FE_OFN491_regtop_g_a_r_3_),
	.b(n245498));
   ao22f01 U265609 (.o(n245506),
	.a(n249652),
	.b(regtop_g_embv_adr_r[4]),
	.c(FE_OFN545_n245460),
	.d(regtop_g_brv_r[4]));
   ao22f01 U265610 (.o(n245496),
	.a(n252998),
	.b(g_field_offset_r[4]),
	.c(n249645),
	.d(regtop_g_adb_cpu_r[4]));
   ao22s01 U265611 (.o(n245495),
	.a(n249787),
	.b(regtop_g_scp_r[4]),
	.c(n249648),
	.d(regtop_g_udb_cpu_r[4]));
   ao22f01 U265612 (.o(n245494),
	.a(n252912),
	.b(g_fcyc_r[4]),
	.c(n249584),
	.d(regtop_g_nfst_r[4]));
   na02s01 U265613 (.o(n245493),
	.a(n249811),
	.b(g_mbc_r[4]));
   ao22f02 U265614 (.o(n245502),
	.a(FE_OFN552_n245462),
	.b(regtop_g_vd_r[4]),
	.c(n249838),
	.d(regtop_g_fcvo1_r[4]));
   ao22f02 U265615 (.o(n245501),
	.a(FE_OFN527_n249828),
	.b(regtop_g_fcvo2_r[4]),
	.c(n249823),
	.d(regtop_g_vsv_r[4]));
   no02f02 U265616 (.o(n249647),
	.a(FE_OFN520_regtop_g_a_r_6_),
	.b(n245497));
   no02f02 U265617 (.o(n249582),
	.a(regtop_g_a_r[3]),
	.b(n245498));
   ao22f03 U265618 (.o(n245500),
	.a(n249647),
	.b(regtop_g_fpst_r[4]),
	.c(n249582),
	.d(regtop_g_fbst_r[4]));
   ao22f01 U265619 (.o(n245499),
	.a(n249813),
	.b(regtop_g_mc_r[4]),
	.c(n249824),
	.d(regtop_g_dvs_r[4]));
   ao22f02 U265620 (.o(n245512),
	.a(g_vs60p_r[4]),
	.b(n249786),
	.c(FE_OFN4_n245443),
	.d(n245509));
   ao12s01 U265621 (.o(n245511),
	.a(n249664),
	.b(n249812),
	.c(regtop_g_tmc_r[4]));
   na02s01 U265622 (.o(n245510),
	.a(n249825),
	.b(regtop_g_vldstatus_r[0]));
   in01f01 U265623 (.o(n245537),
	.a(regtop_g_paramadr_r[7]));
   no02f02 U265624 (.o(n246608),
	.a(regtop_g_paramadr_r[2]),
	.b(regtop_g_paramadr_r[3]));
   in01s01 U265625 (.o(n245516),
	.a(n245515));
   in01s01 U265626 (.o(n245551),
	.a(n245560));
   no02s01 U265627 (.o(n245540),
	.a(n246865),
	.b(n245530));
   in01s01 U265628 (.o(n245522),
	.a(n245540));
   in01s01 U265629 (.o(n245519),
	.a(n245762));
   na02f01 U265630 (.o(n245518),
	.a(regtop_g_paramadr_r[3]),
	.b(n246609));
   no02s01 U265631 (.o(n245520),
	.a(n245519),
	.b(n245848));
   na02s01 U265632 (.o(n245521),
	.a(n245520),
	.b(n252341));
   no02f01 U265633 (.o(n252376),
	.a(n245522),
	.b(n245521));
   no02f02 U265634 (.o(n252380),
	.a(regtop_g_paramadr_r[7]),
	.b(n246609));
   in01f02 U265635 (.o(n252404),
	.a(regtop_g_paramadr_r[2]));
   no02m02 U265636 (.o(n245523),
	.a(regtop_g_paramadr_r[3]),
	.b(n252404));
   na02f03 U265637 (.o(n252517),
	.a(n245527),
	.b(n245523));
   na02s01 U265638 (.o(n245524),
	.a(n252515),
	.b(n245544));
   in01s01 U265639 (.o(n245525),
	.a(n245524));
   no02s01 U265640 (.o(n252374),
	.a(n252676),
	.b(n245530));
   no02s01 U265641 (.o(n252372),
	.a(n245530),
	.b(n252752));
   na02s01 U265642 (.o(n245526),
	.a(regtop_g_paramadr_r[6]),
	.b(regtop_g_nferror_r));
   in01s01 U265643 (.o(n245554),
	.a(n245526));
   na02f01 U265644 (.o(n252826),
	.a(n245554),
	.b(n245939));
   in01s01 U265645 (.o(n245570),
	.a(n245530));
   na02s01 U265646 (.o(n252371),
	.a(n245570),
	.b(n245579));
   in01s01 U265647 (.o(n245535),
	.a(n246865));
   na02s01 U265648 (.o(n245532),
	.a(n245551),
	.b(n252613));
   in01s01 U265649 (.o(n245569),
	.a(n245532));
   in01s01 U265650 (.o(n245534),
	.a(n245533));
   na02f01 U265651 (.o(n252604),
	.a(n245535),
	.b(n245534));
   no02s01 U265652 (.o(n245539),
	.a(n245761),
	.b(n245538));
   na02f01 U265653 (.o(n246840),
	.a(n245540),
	.b(n245539));
   in01s01 U265654 (.o(n252253),
	.a(n252731));
   no02f01 U265655 (.o(n246001),
	.a(n245560),
	.b(n252253));
   na02s01 U265656 (.o(n245541),
	.a(n246001),
	.b(n245544));
   in01s01 U265657 (.o(n245553),
	.a(n245541));
   in01s01 U265658 (.o(n245768),
	.a(regtop_g_paramadr_r[1]));
   ao12s01 U265659 (.o(n245542),
	.a(n252404),
	.b(n252517),
	.c(n245768));
   na02s01 U265660 (.o(n252673),
	.a(n245551),
	.b(n245543));
   no02f01 U265661 (.o(n245558),
	.a(n245560),
	.b(n252575));
   in01s01 U265662 (.o(n245546),
	.a(n245544));
   na02f01 U265663 (.o(n252487),
	.a(n245558),
	.b(n252680));
   in01s01 U265664 (.o(n245548),
	.a(regtop_g_paramadr_r[3]));
   na02m01 U265665 (.o(n245767),
	.a(n252380),
	.b(n245548));
   no02m02 U265666 (.o(n245583),
	.a(n245762),
	.b(n245767));
   no02f01 U265667 (.o(n245549),
	.a(n245583),
	.b(n245763));
   na02f01 U265668 (.o(n245550),
	.a(n245766),
	.b(n245549));
   no02f01 U265669 (.o(n252238),
	.a(regtop_g_paramadr_r[0]),
	.b(n245585));
   na02f01 U265670 (.o(n252489),
	.a(n252567),
	.b(n245558));
   in01s01 U265671 (.o(n245557),
	.a(n252676));
   na02s01 U265672 (.o(n245576),
	.a(n252575),
	.b(n252253));
   na02s01 U265673 (.o(n245555),
	.a(n245554),
	.b(n245576));
   in01s01 U265674 (.o(n245556),
	.a(n245555));
   na02f01 U265675 (.o(n252547),
	.a(n245557),
	.b(n245556));
   na02f01 U265676 (.o(n252491),
	.a(n245558),
	.b(n245939));
   no02s01 U265677 (.o(n245561),
	.a(regtop_g_paramadr_r[1]),
	.b(n245560));
   ao22f01 U265678 (.o(n252606),
	.a(n245561),
	.b(n245583),
	.c(n245579),
	.d(n245569));
   no02s01 U265679 (.o(n245562),
	.a(regtop_g_paramadr_r[2]),
	.b(n246902));
   in01s01 U265680 (.o(n245563),
	.a(n245562));
   no02s01 U265681 (.o(n245564),
	.a(n245763),
	.b(n245563));
   na02s01 U265682 (.o(n245567),
	.a(n245564),
	.b(n252234));
   in01s01 U265683 (.o(n245565),
	.a(n245579));
   na02s01 U265684 (.o(n245566),
	.a(n245565),
	.b(n252752));
   no02f02 U265685 (.o(n252239),
	.a(n245567),
	.b(n245566));
   ao22f01 U265686 (.o(n252608),
	.a(n246001),
	.b(n245568),
	.c(n252239),
	.d(n245569));
   na02s01 U265687 (.o(n245573),
	.a(n252606),
	.b(n252608));
   na02s01 U265688 (.o(n245572),
	.a(n252567),
	.b(n245569));
   na02s01 U265689 (.o(n245571),
	.a(n245570),
	.b(n252680));
   na02s01 U265690 (.o(n252368),
	.a(n245572),
	.b(n245571));
   in01s01 U265691 (.o(n245588),
	.a(n245576));
   na02s01 U265692 (.o(n245577),
	.a(n245763),
	.b(n252404));
   in01s01 U265693 (.o(n245578),
	.a(n245577));
   in01s01 U265694 (.o(n245581),
	.a(n245580));
   in01s01 U265695 (.o(n245584),
	.a(n245582));
   ao12s01 U265696 (.o(n245586),
	.a(n245583),
	.b(n245763),
	.c(n245584));
   na02s01 U265697 (.o(n245587),
	.a(n245586),
	.b(n245585));
   na02f01 U265698 (.o(n252251),
	.a(regtop_g_paramadr_r[6]),
	.b(n245587));
   na02f02 U265699 (.o(n245589),
	.a(n252307),
	.b(regtop_g_nferror_r));
   no02f80 U265700 (.o(n253015),
	.a(regtop_g_write_r_n),
	.b(regtop_g_ms_r_n));
   na03s01 U265701 (.o(n245595),
	.a(n249924),
	.b(regtop_g_isnf_r),
	.c(n252273));
   in01s01 U265702 (.o(vmem_we[2]),
	.a(vmem_we_n[2]));
   in01s01 U265703 (.o(vmem_we[3]),
	.a(vmem_we_n[3]));
   in01s01 U265704 (.o(vmem_we[0]),
	.a(vmem_we_n[0]));
   no02f02 U265705 (.o(n245600),
	.a(n245599),
	.b(n245601));
   no02f01 U265706 (.o(n245603),
	.a(n245599),
	.b(n245600));
   no02f01 U265707 (.o(n245602),
	.a(n245601),
	.b(n245600));
   no02f01 U265708 (.o(busrtop_b_rreq_N105),
	.a(n245603),
	.b(n245602));
   in01s01 U265709 (.o(n245606),
	.a(n245604));
   na02s01 U265710 (.o(n245609),
	.a(n245606),
	.b(n245605));
   na02f01 U265711 (.o(n245608),
	.a(n245607),
	.b(n245609));
   na02f01 U265712 (.o(n245611),
	.a(n245607),
	.b(n245608));
   na02s01 U265713 (.o(n245616),
	.a(n245613),
	.b(n245612));
   no02m01 U265714 (.o(n245615),
	.a(n245614),
	.b(n245616));
   no02m01 U265715 (.o(n245618),
	.a(n245614),
	.b(n245615));
   in01s01 U265716 (.o(n245621),
	.a(n245619));
   na02s01 U265717 (.o(n245624),
	.a(n245621),
	.b(n245620));
   na02m01 U265718 (.o(n245623),
	.a(n245622),
	.b(n245624));
   na02s01 U265719 (.o(n245631),
	.a(n245628),
	.b(n245627));
   in01s01 U265720 (.o(n245636),
	.a(n245634));
   na02s01 U265721 (.o(n245638),
	.a(n245637),
	.b(n245639));
   na02s01 U265722 (.o(n245641),
	.a(n245637),
	.b(n245638));
   na02s01 U265723 (.o(n245640),
	.a(n245639),
	.b(n245638));
   na02s01 U265724 (.o(busrtop_b_rreq_N100),
	.a(n245641),
	.b(n245640));
   na02s01 U265725 (.o(n245646),
	.a(n245643),
	.b(n245642));
   no02s01 U265726 (.o(n245645),
	.a(n245644),
	.b(n245646));
   no02s01 U265727 (.o(n245648),
	.a(n245644),
	.b(n245645));
   no02s01 U265728 (.o(busrtop_b_rreq_N99),
	.a(n245648),
	.b(n245647));
   in01s01 U265729 (.o(n245651),
	.a(n245649));
   na02s01 U265730 (.o(n245654),
	.a(n245651),
	.b(n245650));
   na02s01 U265731 (.o(n245653),
	.a(n245652),
	.b(n245654));
   na02s01 U265732 (.o(n245656),
	.a(n245652),
	.b(n245653));
   na02s01 U265733 (.o(n245655),
	.a(n245654),
	.b(n245653));
   na02s01 U265734 (.o(busrtop_b_rreq_N98),
	.a(n245656),
	.b(n245655));
   na02s01 U265735 (.o(n245661),
	.a(n245658),
	.b(n245657));
   no02s01 U265736 (.o(n245660),
	.a(n245659),
	.b(n245661));
   no02s01 U265737 (.o(n245663),
	.a(n245659),
	.b(n245660));
   no02s01 U265738 (.o(n245662),
	.a(n245661),
	.b(n245660));
   in01s01 U265739 (.o(n245729),
	.a(n245664));
   in01s01 U265740 (.o(n245669),
	.a(n245667));
   na02s01 U265741 (.o(n245672),
	.a(n245669),
	.b(n245668));
   no02s01 U265742 (.o(n245673),
	.a(n245672),
	.b(n245671));
   no02s01 U265743 (.o(busrtop_b_rreq_N92),
	.a(n245674),
	.b(n245673));
   in01s01 U265744 (.o(n245722),
	.a(n245675));
   oa12s01 U265745 (.o(n245681),
	.a(n245676),
	.b(n245722),
	.c(n245677));
   no02s01 U265746 (.o(n245682),
	.a(n245681),
	.b(n245683));
   no02s01 U265747 (.o(n245685),
	.a(n245681),
	.b(n245682));
   no02s01 U265748 (.o(n245684),
	.a(n245683),
	.b(n245682));
   no02s01 U265749 (.o(busrtop_b_rreq_N95),
	.a(n245685),
	.b(n245684));
   na02s01 U265750 (.o(n245691),
	.a(n245688),
	.b(n245687));
   no02s01 U265751 (.o(n245690),
	.a(n245689),
	.b(n245691));
   no02s01 U265752 (.o(n245693),
	.a(n245689),
	.b(n245690));
   no02s01 U265753 (.o(n245692),
	.a(n245691),
	.b(n245690));
   no02s01 U265754 (.o(busrtop_b_rreq_N94),
	.a(n245693),
	.b(n245692));
   in01s01 U265755 (.o(n245696),
	.a(n245694));
   na02s01 U265756 (.o(n245699),
	.a(n245696),
	.b(n245695));
   na02s01 U265757 (.o(n245698),
	.a(n245697),
	.b(n245699));
   na02s01 U265758 (.o(n245701),
	.a(n245697),
	.b(n245698));
   na02s01 U265759 (.o(n245700),
	.a(n245699),
	.b(n245698));
   na02s01 U265760 (.o(busrtop_b_rreq_N96),
	.a(n245701),
	.b(n245700));
   in01s01 U265761 (.o(n245704),
	.a(n245702));
   na02s01 U265762 (.o(n245707),
	.a(n245704),
	.b(n245703));
   na02s01 U265763 (.o(n245706),
	.a(n245705),
	.b(n245707));
   na02s01 U265764 (.o(n245709),
	.a(n245705),
	.b(n245706));
   na02s01 U265765 (.o(n245708),
	.a(n245707),
	.b(n245706));
   na02s01 U265766 (.o(busrtop_b_rreq_N91),
	.a(n245709),
	.b(n245708));
   in01s01 U265767 (.o(n245728),
	.a(n245710));
   in01s01 U265768 (.o(n245711),
	.a(n245727));
   ao12s01 U265769 (.o(n245715),
	.a(n245711),
	.b(n245729),
	.c(n245728));
   in01s01 U265770 (.o(n245714),
	.a(n245712));
   na02s01 U265771 (.o(n245716),
	.a(n245715),
	.b(n245717));
   na02s01 U265772 (.o(n245719),
	.a(n245715),
	.b(n245716));
   na02s01 U265773 (.o(n245718),
	.a(n245717),
	.b(n245716));
   na02s01 U265774 (.o(busrtop_b_rreq_N90),
	.a(n245719),
	.b(n245718));
   na02s01 U265775 (.o(n245724),
	.a(n245721),
	.b(n245720));
   na02s01 U265776 (.o(n245723),
	.a(n245724),
	.b(n245722));
   na02s01 U265777 (.o(n245726),
	.a(n245722),
	.b(n245723));
   na02s01 U265778 (.o(n245725),
	.a(n245724),
	.b(n245723));
   na02s01 U265779 (.o(busrtop_b_rreq_N93),
	.a(n245726),
	.b(n245725));
   na02s01 U265780 (.o(n245731),
	.a(n245728),
	.b(n245727));
   no02s01 U265781 (.o(n245730),
	.a(n245731),
	.b(n245729));
   no02s01 U265782 (.o(n245733),
	.a(n245730),
	.b(n245729));
   no02s01 U265783 (.o(n245732),
	.a(n245731),
	.b(n245730));
   no02s01 U265784 (.o(busrtop_b_rreq_N89),
	.a(n245733),
	.b(n245732));
   in01s01 U265785 (.o(n245746),
	.a(n245734));
   oa12s01 U265786 (.o(n245738),
	.a(n245744),
	.b(n245746),
	.c(n245743));
   in01s01 U265787 (.o(n245737),
	.a(n245735));
   na02s01 U265788 (.o(n245740),
	.a(n245737),
	.b(n245736));
   no02s01 U265789 (.o(n245739),
	.a(n245738),
	.b(n245740));
   no02s01 U265790 (.o(n245742),
	.a(n245738),
	.b(n245739));
   no02s01 U265791 (.o(n245741),
	.a(n245740),
	.b(n245739));
   no02s01 U265792 (.o(busrtop_b_rreq_N88),
	.a(n245742),
	.b(n245741));
   in01s01 U265793 (.o(n245745),
	.a(n245743));
   na02s01 U265794 (.o(n245748),
	.a(n245745),
	.b(n245744));
   na02s01 U265795 (.o(n245747),
	.a(n245748),
	.b(n245746));
   na02s01 U265796 (.o(n245750),
	.a(n245746),
	.b(n245747));
   na02s01 U265797 (.o(n245749),
	.a(n245748),
	.b(n245747));
   na02s01 U265798 (.o(busrtop_b_rreq_N87),
	.a(n245750),
	.b(n245749));
   in01s01 U265799 (.o(n245753),
	.a(n245751));
   na02s01 U265800 (.o(n245754),
	.a(n245753),
	.b(n245752));
   na02s01 U265801 (.o(n245755),
	.a(n245754),
	.b(n245758));
   na02s01 U265802 (.o(n245757),
	.a(n245754),
	.b(n245755));
   na02s01 U265803 (.o(n245756),
	.a(n245758),
	.b(n245755));
   na02s01 U265804 (.o(busrtop_b_rreq_N86),
	.a(n245757),
	.b(n245756));
   no02s01 U265805 (.o(n245760),
	.a(busrtop_b_rreq_N295),
	.b(n245758));
   no02s01 U265806 (.o(n245759),
	.a(n245758),
	.b(g_field_start_add_r[10]));
   no02s01 U265807 (.o(busrtop_b_rreq_N85),
	.a(n245760),
	.b(n245759));
   in01s01 U265808 (.o(n245772),
	.a(n252380));
   in01f01 U265809 (.o(n245771),
	.a(n245766));
   in01s01 U265810 (.o(n245769),
	.a(n245767));
   in01s01 U265811 (.o(n245778),
	.a(n245777));
   in01f02 U265812 (.o(n253125),
	.a(busiftop_status_b_current_0_));
   in01s01 U265813 (.o(n252904),
	.a(g_pcut_r[9]));
   in01s01 U265814 (.o(n252893),
	.a(g_pcut_r[2]));
   in01s01 U265815 (.o(n252898),
	.a(g_pcut_r[5]));
   na02s01 U265816 (.o(n245779),
	.a(n252893),
	.b(n252898));
   in01s01 U265817 (.o(n245780),
	.a(n245779));
   na02s01 U265818 (.o(n245781),
	.a(n252895),
	.b(n245780));
   in01s01 U265819 (.o(n245782),
	.a(n245781));
   na02s01 U265820 (.o(n245794),
	.a(n252904),
	.b(n245782));
   in01s01 U265821 (.o(n252900),
	.a(g_pcut_r[6]));
   in01f01 U265822 (.o(n252897),
	.a(g_pcut_r[4]));
   in01s01 U265823 (.o(n252906),
	.a(g_pcut_r[10]));
   in01s01 U265824 (.o(n252903),
	.a(g_pcut_r[8]));
   na02s01 U265825 (.o(n245783),
	.a(n252906),
	.b(n252903));
   in01s01 U265826 (.o(n245784),
	.a(n245783));
   na02s01 U265827 (.o(n245785),
	.a(n252897),
	.b(n245784));
   in01s01 U265828 (.o(n245786),
	.a(n245785));
   na02s01 U265829 (.o(n245793),
	.a(n252900),
	.b(n245786));
   in01s01 U265830 (.o(n252908),
	.a(g_pcut_r[11]));
   in01s01 U265831 (.o(n245789),
	.a(g_pcut_r[7]));
   in01s01 U265832 (.o(n252892),
	.a(g_pcut_r[1]));
   in01s01 U265833 (.o(n252911),
	.a(g_pcut_r[0]));
   na02s01 U265834 (.o(n245787),
	.a(n252892),
	.b(g_pcut_r[0]));
   in01s01 U265835 (.o(n245788),
	.a(n245787));
   na02s01 U265836 (.o(n245790),
	.a(n245789),
	.b(n245788));
   in01s01 U265837 (.o(n245791),
	.a(n245790));
   in01s01 U265839 (.o(n252947),
	.a(g_pmod_r));
   no02f01 U265840 (.o(cntrltop_ctmg_ctpedet_c_tmg_ferr_pre),
	.a(cntrltop_ctmg_ctpedet_c_bigpictdet_r),
	.b(n252288));
   in01s01 U265841 (.o(n245796),
	.a(regtop_v1_hdi00_bs));
   no02s01 U265842 (.o(regtop_N1991),
	.a(regtop_v1_hdi00_we),
	.b(n245796));
   na02s01 U265843 (.o(n249307),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[19]));
   oa12s01 U265844 (.o(busiftop_N36),
	.a(n249307),
	.b(busiftop_vmem_ch_r),
	.c(vh_1_ph_add[0]));
   in01s01 U265845 (.o(n246214),
	.a(busrtop_b_rreq_vrh_cnt_16byte_r[0]));
   na02s01 U265846 (.o(n245797),
	.a(busiftop_status_b_current_0_),
	.b(n246214));
   oa12s01 U265847 (.o(n170939),
	.a(n245797),
	.b(busiftop_status_b_current_0_),
	.c(n246214));
   no02f02 U265848 (.o(n247029),
	.a(vldtop_vld_syndec_vld_seqhed_state_0_),
	.b(n249027));
   na02s01 U265849 (.o(vldtop_vld_syndec_vld_outbuf_N46),
	.a(g_swrst_r_n),
	.b(n247029));
   no02s01 U265850 (.o(n245798),
	.a(v_seqstrt_r),
	.b(vldtop_vld_syndec_vld_seqhed_state_0_));
   in01s01 U265851 (.o(n245799),
	.a(n245798));
   na02s01 U265852 (.o(vldtop_vld_syndec_vld_outbuf_N52),
	.a(g_swrst_r_n),
	.b(n245799));
   no02s01 U265853 (.o(n245812),
	.a(vh_1_ph_add[1]),
	.b(vh_1_ph_add[27]));
   in01s01 U265854 (.o(n245800),
	.a(n245812));
   na02s01 U265855 (.o(n245810),
	.a(vh_1_ph_add[1]),
	.b(vh_1_ph_add[27]));
   na02s01 U265856 (.o(n245801),
	.a(n245800),
	.b(n245810));
   in01s01 U265857 (.o(n245811),
	.a(vh_1_ph_add[0]));
   na02s01 U265858 (.o(n245802),
	.a(n245801),
	.b(n245811));
   na02s01 U265859 (.o(n245804),
	.a(n245801),
	.b(n245802));
   na02s01 U265860 (.o(n245803),
	.a(n245811),
	.b(n245802));
   na02s01 U265861 (.o(n245805),
	.a(n245804),
	.b(n245803));
   in01s01 U265862 (.o(n245806),
	.a(n245805));
   na02s01 U265863 (.o(n249308),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[20]));
   oa12s01 U265864 (.o(busiftop_N37),
	.a(n249308),
	.b(busiftop_vmem_ch_r),
	.c(n245806));
   in01s01 U265865 (.o(n249021),
	.a(v_vldstatus_r[0]));
   na02s01 U265866 (.o(n249023),
	.a(n246731),
	.b(n246796));
   in01s01 U265867 (.o(n245809),
	.a(n249023));
   in01s01 U265868 (.o(n245807),
	.a(y1_bs_wait_n));
   na02s01 U265869 (.o(n245808),
	.a(n245807),
	.b(n249015));
   na02s01 U265870 (.o(n249022),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n245808));
   oa22s01 U265871 (.o(n243163),
	.a(n245809),
	.b(n249022),
	.c(n249028),
	.d(n246731));
   in01s01 U265872 (.o(n245829),
	.a(n245823));
   in01s01 U265873 (.o(n245813),
	.a(n245828));
   na02s01 U265874 (.o(n245815),
	.a(n245813),
	.b(n245827));
   na02s01 U265875 (.o(n245817),
	.a(n245829),
	.b(n245814));
   na02s01 U265876 (.o(n245816),
	.a(n245815),
	.b(n245814));
   na02s01 U265877 (.o(n245818),
	.a(n245817),
	.b(n245816));
   na02s01 U265878 (.o(n249309),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[21]));
   oa12s01 U265879 (.o(busiftop_N38),
	.a(n249309),
	.b(busiftop_vmem_ch_r),
	.c(n245819));
   na02s01 U265880 (.o(n245831),
	.a(vh_1_ph_add[3]),
	.b(vh_1_ph_add[29]));
   na02s01 U265881 (.o(n245857),
	.a(vh_1_ph_add[5]),
	.b(vh_1_ph_add[31]));
   na02s01 U265882 (.o(n249294),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[4]));
   oa12s01 U265883 (.o(busiftop_N59),
	.a(n249294),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   na02s01 U265884 (.o(n249296),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[6]));
   oa12s01 U265885 (.o(busiftop_N61),
	.a(n249296),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   oa12s01 U265886 (.o(n245833),
	.a(n245827),
	.b(n245829),
	.c(n245828));
   na02s01 U265887 (.o(n245835),
	.a(n245832),
	.b(n245831));
   no02s01 U265888 (.o(n245834),
	.a(n245833),
	.b(n245835));
   no02s01 U265889 (.o(n245837),
	.a(n245833),
	.b(n245834));
   no02s01 U265890 (.o(n245836),
	.a(n245835),
	.b(n245834));
   no02s01 U265891 (.o(n245838),
	.a(n245837),
	.b(n245836));
   in01s01 U265892 (.o(n245839),
	.a(n245838));
   na02s01 U265893 (.o(n249310),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[22]));
   oa12s01 U265894 (.o(busiftop_N39),
	.a(n249310),
	.b(busiftop_vmem_ch_r),
	.c(n245839));
   in01s01 U265895 (.o(n245855),
	.a(n245841));
   na02s01 U265896 (.o(n245843),
	.a(n245855),
	.b(n245853));
   no02s01 U265897 (.o(n245842),
	.a(n245899),
	.b(n245843));
   no02s01 U265898 (.o(n245845),
	.a(n245899),
	.b(n245842));
   no02s01 U265899 (.o(n245844),
	.a(n245843),
	.b(n245842));
   no02s01 U265900 (.o(n245846),
	.a(n245845),
	.b(n245844));
   in01s01 U265901 (.o(n245847),
	.a(n245846));
   na02s01 U265902 (.o(n249311),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[23]));
   oa12s01 U265903 (.o(busiftop_N40),
	.a(n249311),
	.b(busiftop_vmem_ch_r),
	.c(n245847));
   in01s01 U265904 (.o(n252600),
	.a(regtop_g_adb_r[0]));
   in01f06 U265905 (.o(n252755),
	.a(regtop_g_paramdata_r[24]));
   in01s01 U265906 (.o(n252599),
	.a(regtop_g_adb_r[1]));
   na02f01 U265907 (.o(n245851),
	.a(FE_OFN218_n246238),
	.b(n252599));
   na02s01 U265908 (.o(n245850),
	.a(regtop_g_atscd_r[23]),
	.b(n245851));
   oa12s01 U265909 (.o(n212112),
	.a(n245850),
	.b(n245924),
	.c(n252755));
   na02s01 U265910 (.o(n245852),
	.a(regtop_g_atscd_r[22]),
	.b(n245851));
   oa12s01 U265911 (.o(n212111),
	.a(n245852),
	.b(n245924),
	.c(n252778));
   in01s01 U265912 (.o(n245854),
	.a(n245853));
   in01s01 U265913 (.o(n245858),
	.a(n245856));
   na02s01 U265914 (.o(n245861),
	.a(n245858),
	.b(n245857));
   na02s01 U265915 (.o(n245860),
	.a(n245859),
	.b(n245861));
   na02s01 U265916 (.o(n245863),
	.a(n245859),
	.b(n245860));
   in01s01 U265917 (.o(n245865),
	.a(n245864));
   na02s01 U265918 (.o(n246210),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[24]));
   in01s01 U265919 (.o(n245894),
	.a(n245887));
   no02s01 U265920 (.o(n245867),
	.a(n245894),
	.b(n249871));
   in01s01 U265921 (.o(n245896),
	.a(n245886));
   no02s01 U265922 (.o(n245866),
	.a(n245896),
	.b(n249871));
   in01s01 U265923 (.o(n245870),
	.a(vh_1_ph_add[7]));
   na02s01 U265924 (.o(n245869),
	.a(n245868),
	.b(n245870));
   na02s01 U265925 (.o(n245872),
	.a(n245868),
	.b(n245869));
   na02s01 U265926 (.o(n245871),
	.a(n245870),
	.b(n245869));
   na02s01 U265927 (.o(n245873),
	.a(n245872),
	.b(n245871));
   in01s01 U265928 (.o(n245874),
	.a(n245873));
   na02f01 U265929 (.o(n246211),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[12]));
   oa12s01 U265930 (.o(busiftop_N43),
	.a(n246211),
	.b(busiftop_vmem_ch_r),
	.c(n245874));
   no02s01 U265931 (.o(n245878),
	.a(n245876),
	.b(n245894));
   no02s01 U265932 (.o(n245877),
	.a(n245876),
	.b(n245896));
   in01s01 U265933 (.o(n245881),
	.a(vh_1_ph_add[9]));
   na02s01 U265934 (.o(n245880),
	.a(n245879),
	.b(n245881));
   na02s01 U265935 (.o(n245883),
	.a(n245879),
	.b(n245880));
   na02s01 U265936 (.o(n245882),
	.a(n245881),
	.b(n245880));
   na02s01 U265937 (.o(n245884),
	.a(n245883),
	.b(n245882));
   in01s01 U265938 (.o(n245885),
	.a(n245884));
   na02s01 U265939 (.o(n249302),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[14]));
   oa12s01 U265940 (.o(busiftop_N45),
	.a(n249302),
	.b(busiftop_vmem_ch_r),
	.c(n245885));
   na02s01 U265941 (.o(n245889),
	.a(n245888),
	.b(n249871));
   na02s01 U265942 (.o(n245891),
	.a(n245888),
	.b(n245889));
   na02s01 U265943 (.o(n245890),
	.a(n249871),
	.b(n245889));
   na02s01 U265944 (.o(n245892),
	.a(n245891),
	.b(n245890));
   in01s01 U265945 (.o(n245893),
	.a(n245892));
   na02s01 U265946 (.o(n246209),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[25]));
   oa12s01 U265947 (.o(busiftop_N42),
	.a(n246209),
	.b(busiftop_vmem_ch_r),
	.c(n245893));
   no02s01 U265948 (.o(n245898),
	.a(n245894),
	.b(n245895));
   no02s01 U265949 (.o(n245897),
	.a(n245896),
	.b(n245895));
   in01s01 U265950 (.o(n249856),
	.a(vh_1_ph_add[8]));
   na02s01 U265951 (.o(n245901),
	.a(n245900),
	.b(n249856));
   na02s01 U265952 (.o(n245903),
	.a(n245900),
	.b(n245901));
   na02s01 U265953 (.o(n245902),
	.a(n249856),
	.b(n245901));
   na02s01 U265954 (.o(n245904),
	.a(n245903),
	.b(n245902));
   in01s01 U265955 (.o(n245905),
	.a(n245904));
   na02f80 U265956 (.o(n249301),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[13]));
   oa12s01 U265957 (.o(busiftop_N44),
	.a(n249301),
	.b(busiftop_vmem_ch_r),
	.c(n245905));
   in01s01 U265958 (.o(n245906),
	.a(regtop_g_atscd_r[19]));
   na02f03 U265959 (.o(n249078),
	.a(regtop_g_adb_r[1]),
	.b(FE_OFN218_n246238));
   oa12s01 U265962 (.o(n212108),
	.a(n245908),
	.b(n252662),
	.c(n245924));
   in01f04 U265963 (.o(n252656),
	.a(regtop_g_paramdata_r[17]));
   in01s01 U265964 (.o(n245909),
	.a(regtop_g_atscd_r[16]));
   oa12s01 U265966 (.o(n212105),
	.a(n245911),
	.b(n252656),
	.c(n245924));
   in01s01 U265967 (.o(n245912),
	.a(regtop_g_atscd_r[21]));
   oa12s01 U265970 (.o(n212110),
	.a(n245914),
	.b(n252666),
	.c(n245924));
   in01f04 U265971 (.o(n252658),
	.a(regtop_g_paramdata_r[18]));
   in01s01 U265972 (.o(n245915),
	.a(regtop_g_atscd_r[17]));
   oa12s01 U265975 (.o(n212106),
	.a(n245917),
	.b(n252658),
	.c(n245924));
   in01s01 U265976 (.o(n245918),
	.a(regtop_g_atscd_r[20]));
   oa12s01 U265979 (.o(n212109),
	.a(n245920),
	.b(n252664),
	.c(n245924));
   in01s01 U265980 (.o(n245921),
	.a(regtop_g_atscd_r[18]));
   oa22s01 U265981 (.o(n245922),
	.a(FE_OFN218_n246238),
	.b(n245921),
	.c(n245921),
	.d(n249078));
   in01s01 U265982 (.o(n245923),
	.a(n245922));
   oa12s01 U265983 (.o(n212107),
	.a(n245923),
	.b(n252660),
	.c(n245924));
   in01s01 U265984 (.o(n249354),
	.a(regtop_g_init_cnt_r[2]));
   no02s01 U265985 (.o(n249355),
	.a(regtop_g_init_cnt_r[1]),
	.b(regtop_g_init_cnt_r[0]));
   na02f02 U265986 (.o(n252873),
	.a(n249354),
	.b(n249355));
   in01f08 U265987 (.o(n247591),
	.a(g_swrst_r_n));
   ao12s01 U265988 (.o(n212680),
	.a(FE_OFN492_n252377),
	.b(n252873),
	.c(n247591));
   in01s01 U265989 (.o(n246034),
	.a(vldtop_vld_syndec_UREG[0]));
   in01s01 U265990 (.o(n245925),
	.a(vldtop_vld_syndec_UREG[2]));
   ao22f01 U265991 (.o(n246498),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n246034),
	.c(n246419),
	.d(n245925));
   no02s01 U265992 (.o(n246402),
	.a(n246498),
	.b(n246697));
   in01s01 U265993 (.o(n247332),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[28]));
   na02s01 U265994 (.o(n245927),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n247332));
   in01s01 U265995 (.o(n247163),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[30]));
   na02s01 U265996 (.o(n245926),
	.a(n246419),
	.b(n247163));
   na02f02 U265997 (.o(n246564),
	.a(n245927),
	.b(n245926));
   in01s01 U265998 (.o(n245928),
	.a(n246564));
   na02f03 U265999 (.o(n246693),
	.a(vldtop_vld_syndec_ADP[2]),
	.b(vldtop_vld_syndec_ADP[3]));
   no02s01 U266000 (.o(n246403),
	.a(n245928),
	.b(n246693));
   na02s01 U266001 (.o(n245930),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n246359));
   in01s01 U266002 (.o(n246043),
	.a(vldtop_vld_syndec_UREG[10]));
   na02s01 U266003 (.o(n245929),
	.a(n246419),
	.b(n246043));
   na02f01 U266004 (.o(n246577),
	.a(n245930),
	.b(n245929));
   in01s01 U266005 (.o(n246379),
	.a(n246577));
   no02f06 U266006 (.o(n246568),
	.a(vldtop_vld_syndec_ADP[3]),
	.b(vldtop_vld_syndec_ADP[2]));
   in01f01 U266007 (.o(n246695),
	.a(n246568));
   in01s01 U266008 (.o(n245931),
	.a(vldtop_vld_syndec_UREG[4]));
   na02s01 U266009 (.o(n245933),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n245931));
   in01s01 U266010 (.o(n249001),
	.a(vldtop_vld_syndec_UREG[6]));
   na02s01 U266011 (.o(n245932),
	.a(n246419),
	.b(n249001));
   na02f02 U266012 (.o(n246567),
	.a(n245933),
	.b(n245932));
   in01s01 U266013 (.o(n246380),
	.a(n246567));
   na02f03 U266014 (.o(n246527),
	.a(vldtop_vld_syndec_ADP[2]),
	.b(n246743));
   na02f03 U266015 (.o(n246708),
	.a(n246568),
	.b(n246670));
   in01s01 U266016 (.o(n246658),
	.a(n246708));
   in01f01 U266017 (.o(n246783),
	.a(vldtop_vld_syndec_UREG[24]));
   in01s01 U266018 (.o(n246325),
	.a(vldtop_vld_syndec_UREG[26]));
   oa22f01 U266019 (.o(n246543),
	.a(n246419),
	.b(n246783),
	.c(vldtop_vld_syndec_ADP[1]),
	.d(n246325));
   in01f04 U266020 (.o(n246670),
	.a(vldtop_vld_syndec_ADP[4]));
   in01s01 U266021 (.o(n246039),
	.a(vldtop_vld_syndec_UREG[16]));
   in01s01 U266022 (.o(n246047),
	.a(vldtop_vld_syndec_UREG[18]));
   ao22s01 U266023 (.o(n246492),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n246039),
	.c(n246419),
	.d(n246047));
   na02f03 U266024 (.o(n246578),
	.a(n246570),
	.b(n246670));
   na02s01 U266025 (.o(n246555),
	.a(n246419),
	.b(n246038));
   in01s01 U266026 (.o(n246044),
	.a(vldtop_vld_syndec_UREG[12]));
   na02s01 U266027 (.o(n246554),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n246044));
   na02f01 U266028 (.o(n246576),
	.a(n246555),
	.b(n246554));
   in01s01 U266029 (.o(n246377),
	.a(n246576));
   na02f04 U266030 (.o(n246714),
	.a(n246700),
	.b(n246670));
   in01s01 U266031 (.o(n246048),
	.a(vldtop_vld_syndec_UREG[20]));
   oa22s01 U266032 (.o(n246546),
	.a(n246419),
	.b(n246048),
	.c(vldtop_vld_syndec_ADP[1]),
	.d(n246037));
   no02s01 U266033 (.o(vldtop_vld_syndec_vld_outbuf_N482),
	.a(n246890),
	.b(n247591));
   in01s01 U266034 (.o(n245941),
	.a(regtop_g_vsv_r[9]));
   in01s01 U266035 (.o(n252670),
	.a(regtop_g_paramdata_r[10]));
   oa22s01 U266036 (.o(n211937),
	.a(FE_OFN488_n245940),
	.b(n245941),
	.c(n252670),
	.d(n246585));
   oa12s01 U266037 (.o(busiftop_N46),
	.a(n249303),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   na02s01 U266038 (.o(n249295),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[5]));
   oa12s01 U266039 (.o(busiftop_N60),
	.a(n249295),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   oa12s01 U266040 (.o(busiftop_N54),
	.a(n246211),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   na02s01 U266041 (.o(n249293),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[3]));
   oa12s01 U266042 (.o(busiftop_N57),
	.a(n249292),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   na02f03 U266043 (.o(n249291),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[1]));
   oa12s01 U266044 (.o(busiftop_N56),
	.a(n249291),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   na02s01 U266045 (.o(n249306),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[18]));
   oa12s01 U266046 (.o(busiftop_N49),
	.a(n249306),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   na02s01 U266047 (.o(n249305),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[17]));
   oa12s01 U266048 (.o(busiftop_N48),
	.a(n249305),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   na02f03 U266049 (.o(n249298),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[9]));
   oa12s01 U266050 (.o(busiftop_N51),
	.a(n249298),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   na02f03 U266051 (.o(n249290),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[0]));
   oa12s01 U266052 (.o(busiftop_N55),
	.a(n249290),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   in01s01 U266053 (.o(n245945),
	.a(regtop_g_atscd_r[12]));
   oa22s01 U266054 (.o(n245946),
	.a(FE_OFN218_n246238),
	.b(n245945),
	.c(n245945),
	.d(n249140));
   in01s01 U266055 (.o(n245947),
	.a(n245946));
   oa12s01 U266056 (.o(n212101),
	.a(n245947),
	.b(n252664),
	.c(n249247));
   in01s01 U266057 (.o(n245948),
	.a(regtop_g_atscd_r[13]));
   oa22s01 U266058 (.o(n245949),
	.a(FE_OFN218_n246238),
	.b(n245948),
	.c(n245948),
	.d(n249140));
   in01s01 U266059 (.o(n245950),
	.a(n245949));
   oa12s01 U266060 (.o(n212102),
	.a(n245950),
	.b(n252666),
	.c(n249247));
   in01s01 U266061 (.o(n245951),
	.a(regtop_g_atscd_r[15]));
   oa22s01 U266062 (.o(n245952),
	.a(FE_OFN218_n246238),
	.b(n245951),
	.c(n245951),
	.d(n249140));
   in01s01 U266063 (.o(n245953),
	.a(n245952));
   oa12s01 U266064 (.o(n212104),
	.a(n245953),
	.b(n252755),
	.c(n249247));
   in01s01 U266065 (.o(n245954),
	.a(regtop_g_atscd_r[11]));
   oa22s01 U266066 (.o(n245955),
	.a(FE_OFN218_n246238),
	.b(n245954),
	.c(n245954),
	.d(n249140));
   in01s01 U266067 (.o(n245956),
	.a(n245955));
   oa12s01 U266068 (.o(n212100),
	.a(n245956),
	.b(n252662),
	.c(n249247));
   in01s01 U266069 (.o(n245957),
	.a(regtop_g_atscd_r[14]));
   oa22s01 U266070 (.o(n245958),
	.a(FE_OFN218_n246238),
	.b(n245957),
	.c(n245957),
	.d(n249140));
   in01s01 U266071 (.o(n245959),
	.a(n245958));
   oa12s01 U266072 (.o(n212103),
	.a(n245959),
	.b(n252778),
	.c(n249247));
   oa22s01 U266073 (.o(n245961),
	.a(FE_OFN218_n246238),
	.b(n245960),
	.c(n245960),
	.d(n249140));
   in01s01 U266074 (.o(n245962),
	.a(n245961));
   oa12s01 U266075 (.o(n212121),
	.a(n245962),
	.b(n252656),
	.c(n249247));
   in01s01 U266076 (.o(n245963),
	.a(regtop_g_atscd_r[10]));
   oa22s01 U266077 (.o(n245964),
	.a(FE_OFN218_n246238),
	.b(n245963),
	.c(n245963),
	.d(n249140));
   in01s01 U266078 (.o(n245965),
	.a(n245964));
   oa12s01 U266079 (.o(n212099),
	.a(n245965),
	.b(n252660),
	.c(n249247));
   oa22s01 U266080 (.o(n245967),
	.a(FE_OFN218_n246238),
	.b(n245966),
	.c(n245966),
	.d(n249140));
   in01s01 U266081 (.o(n245968),
	.a(n245967));
   oa12s01 U266082 (.o(n212098),
	.a(n245968),
	.b(n252658),
	.c(n249247));
   na02s01 U266083 (.o(n249299),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[10]));
   oa12s01 U266084 (.o(busiftop_N52),
	.a(n249299),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   na02s01 U266085 (.o(n249297),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[8]));
   oa12s01 U266086 (.o(busiftop_N50),
	.a(n249297),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   na02s01 U266087 (.o(n249300),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[11]));
   oa12s01 U266088 (.o(busiftop_N53),
	.a(n249300),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   na02s01 U266089 (.o(n249304),
	.a(busiftop_vmem_ch_r),
	.b(y1_bs_data_r[16]));
   oa12s01 U266090 (.o(busiftop_N47),
	.a(n249304),
	.b(busiftop_vmem_ch_r),
	.c(n245942));
   no02f01 U266091 (.o(n246289),
	.a(vldtop_vld_syndec_UREG[15]),
	.b(n246419));
   no02s01 U266092 (.o(n246293),
	.a(vldtop_vld_syndec_UREG[17]),
	.b(vldtop_vld_syndec_ADP[1]));
   no02s01 U266093 (.o(n245970),
	.a(n246289),
	.b(n246293));
   in01s01 U266094 (.o(n246341),
	.a(n245970));
   no02s01 U266095 (.o(n245976),
	.a(n246711),
	.b(n246341));
   in01s01 U266096 (.o(n246019),
	.a(vldtop_vld_syndec_UREG[21]));
   in01s01 U266097 (.o(n246016),
	.a(vldtop_vld_syndec_UREG[19]));
   oa22f01 U266098 (.o(n246337),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n246019),
	.c(n246016),
	.d(n246419));
   in01s01 U266099 (.o(n246285),
	.a(n245971));
   oa22f02 U266100 (.o(n246340),
	.a(vldtop_vld_syndec_UREG[11]),
	.b(n246419),
	.c(vldtop_vld_syndec_UREG[13]),
	.d(vldtop_vld_syndec_ADP[1]));
   in01s01 U266101 (.o(n245972),
	.a(n246340));
   in01s01 U266102 (.o(n245978),
	.a(vldtop_vld_syndec_UREG[3]));
   in01s01 U266103 (.o(n245977),
	.a(vldtop_vld_syndec_UREG[5]));
   ao22f01 U266104 (.o(n246297),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n245978),
	.c(n246419),
	.d(n245977));
   in01s01 U266105 (.o(n246344),
	.a(n246297));
   in01s01 U266106 (.o(n247210),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[27]));
   in01s01 U266107 (.o(n247289),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[29]));
   ao22f01 U266108 (.o(n245979),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n247210),
	.c(n246419),
	.d(n247289));
   in01s01 U266109 (.o(n246465),
	.a(n245979));
   oa22f01 U266110 (.o(n246312),
	.a(vldtop_vld_syndec_UREG[9]),
	.b(vldtop_vld_syndec_ADP[1]),
	.c(vldtop_vld_syndec_UREG[7]),
	.d(n246419));
   in01s01 U266111 (.o(n246338),
	.a(n246312));
   in01s01 U266112 (.o(n247159),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[31]));
   in01s01 U266113 (.o(n245980),
	.a(vldtop_vld_syndec_UREG[1]));
   ao22f01 U266114 (.o(n245981),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n247159),
	.c(n246419),
	.d(n245980));
   in01f01 U266115 (.o(n246345),
	.a(n245981));
   na02s01 U266116 (.o(n245982),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246444));
   no02s01 U266117 (.o(n245983),
	.a(n246446),
	.b(n245982));
   na02s01 U266118 (.o(n245984),
	.a(n246448),
	.b(n245983));
   in01s01 U266119 (.o(n246056),
	.a(n245986));
   no02s01 U266120 (.o(vldtop_vld_syndec_vld_outbuf_N481),
	.a(n246056),
	.b(n247591));
   no04s01 U266121 (.o(n245991),
	.a(y1_bs_data_r[20]),
	.b(y1_bs_data_r[21]),
	.c(y1_bs_data_r[22]),
	.d(y1_bs_data_r[23]));
   no04s01 U266122 (.o(n245990),
	.a(y1_bs_data_r[16]),
	.b(y1_bs_data_r[17]),
	.c(y1_bs_data_r[18]),
	.d(y1_bs_data_r[19]));
   no03f01 U266123 (.o(n245989),
	.a(y1_bs_data_r[29]),
	.b(y1_bs_data_r[27]),
	.c(y1_bs_data_r[26]));
   no03s01 U266124 (.o(n245988),
	.a(y1_bs_data_r[24]),
	.b(y1_bs_data_r[25]),
	.c(n245987));
   in01s01 U266125 (.o(n245999),
	.a(n245992));
   no04s01 U266126 (.o(n245996),
	.a(y1_bs_data_r[2]),
	.b(y1_bs_data_r[4]),
	.c(y1_bs_data_r[6]),
	.d(y1_bs_data_r[7]));
   no03s01 U266127 (.o(n245995),
	.a(y1_bs_data_r[31]),
	.b(y1_bs_data_r[0]),
	.c(y1_bs_data_r[1]));
   no04s01 U266128 (.o(n245994),
	.a(y1_bs_data_r[12]),
	.b(y1_bs_data_r[13]),
	.c(y1_bs_data_r[14]),
	.d(y1_bs_data_r[15]));
   in01s01 U266129 (.o(n245998),
	.a(n245997));
   na02f04 U266130 (.o(busiftop_N28),
	.a(n246000),
	.b(vmem_ch));
   na02s01 U266131 (.o(n252682),
	.a(n246001),
	.b(n252377));
   na02s01 U266132 (.o(n246005),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n247289));
   na02s01 U266133 (.o(n246004),
	.a(n246419),
	.b(n247159));
   na02f02 U266134 (.o(n246699),
	.a(n246005),
	.b(n246004));
   in01s01 U266135 (.o(n246006),
	.a(vldtop_vld_syndec_UREG[9]));
   na02s01 U266136 (.o(n246009),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n246006));
   in01s01 U266137 (.o(n246007),
	.a(vldtop_vld_syndec_UREG[11]));
   na02s01 U266138 (.o(n246008),
	.a(n246419),
	.b(n246007));
   no02s01 U266139 (.o(n246011),
	.a(vldtop_vld_syndec_UREG[5]),
	.b(n246419));
   no02s01 U266140 (.o(n246010),
	.a(vldtop_vld_syndec_UREG[7]),
	.b(vldtop_vld_syndec_ADP[1]));
   no02s01 U266141 (.o(n246303),
	.a(n246707),
	.b(n246527));
   oa22s01 U266142 (.o(n246012),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(vldtop_vld_syndec_UREG[3]),
	.c(vldtop_vld_syndec_UREG[1]),
	.d(n246419));
   in01f01 U266143 (.o(n246696),
	.a(n246012));
   no02s01 U266144 (.o(n246302),
	.a(n246696),
	.b(n246697));
   ao22f01 U266145 (.o(n246651),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(vldtop_vld_syndec_UREG[25]),
	.c(n246419),
	.d(vldtop_vld_syndec_UREG[27]));
   in01s01 U266146 (.o(n246014),
	.a(vldtop_vld_syndec_UREG[13]));
   in01s01 U266147 (.o(n246013),
	.a(vldtop_vld_syndec_UREG[15]));
   ao22s01 U266148 (.o(n246015),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n246014),
	.c(n246419),
	.d(n246013));
   in01s01 U266149 (.o(n246715),
	.a(n246015));
   in01s01 U266150 (.o(n246017),
	.a(vldtop_vld_syndec_UREG[17]));
   oa22s01 U266151 (.o(n246650),
	.a(n246419),
	.b(n246017),
	.c(vldtop_vld_syndec_ADP[1]),
	.d(n246016));
   in01s01 U266152 (.o(n246709),
	.a(n246650));
   in01s01 U266153 (.o(n246018),
	.a(vldtop_vld_syndec_UREG[23]));
   oa22s01 U266154 (.o(n246663),
	.a(n246419),
	.b(n246019),
	.c(vldtop_vld_syndec_ADP[1]),
	.d(n246018));
   in01s01 U266155 (.o(n246023),
	.a(n246022));
   no02s01 U266156 (.o(n246027),
	.a(vldtop_vld_syndec_UREG[2]),
	.b(n246419));
   no02s01 U266157 (.o(n246026),
	.a(vldtop_vld_syndec_UREG[4]),
	.b(vldtop_vld_syndec_ADP[1]));
   no02f01 U266158 (.o(n246430),
	.a(n246027),
	.b(n246026));
   na02s01 U266160 (.o(n246028),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(FE_OFN543_vldtop_vld_syndec_vld_vlfeed_lower_26_));
   in01s01 U266161 (.o(n246031),
	.a(n246028));
   na02s01 U266162 (.o(n246029),
	.a(n246419),
	.b(n247332));
   in01s01 U266163 (.o(n246030),
	.a(n246029));
   na02s01 U266164 (.o(n246033),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n249001));
   na02s01 U266165 (.o(n246032),
	.a(n246419),
	.b(n246359));
   na02f02 U266166 (.o(n246536),
	.a(n246033),
	.b(n246032));
   na02f01 U266167 (.o(n246036),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n247163));
   na02s01 U266168 (.o(n246035),
	.a(n246419),
	.b(n246034));
   na02f02 U266169 (.o(n246524),
	.a(n246036),
	.b(n246035));
   na02s01 U266170 (.o(n246415),
	.a(n246565),
	.b(n246524));
   na03s01 U266171 (.o(n246054),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246414),
	.c(n246415));
   oa22s01 U266172 (.o(n246327),
	.a(n246419),
	.b(n246037),
	.c(vldtop_vld_syndec_ADP[1]),
	.d(n246783));
   in01s01 U266173 (.o(n246042),
	.a(n246327));
   na02s01 U266174 (.o(n246041),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n246038));
   na02s01 U266175 (.o(n246040),
	.a(n246419),
	.b(n246039));
   na02f06 U266176 (.o(n246533),
	.a(n246041),
	.b(n246040));
   na02s01 U266177 (.o(n246046),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n246043));
   na02s01 U266178 (.o(n246045),
	.a(n246419),
	.b(n246044));
   na02f02 U266179 (.o(n246535),
	.a(n246046),
	.b(n246045));
   na02s01 U266180 (.o(n246050),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n246047));
   na02f01 U266181 (.o(n246435),
	.a(n246050),
	.b(n246049));
   in01s01 U266182 (.o(n246301),
	.a(n246055));
   in01s01 U266183 (.o(n246057),
	.a(n247000));
   no02m01 U266184 (.o(vldtop_vld_syndec_vld_outbuf_N44),
	.a(n246059),
	.b(n247591));
   in01s01 U266185 (.o(n246061),
	.a(n246060));
   na02f01 U266186 (.o(n246167),
	.a(regtop_g_udb1_r[0]),
	.b(regtop_g_udb0_r[0]));
   na02f02 U266187 (.o(n246064),
	.a(regtop_g_udb0_r[1]),
	.b(n246073));
   na02f02 U266188 (.o(n246063),
	.a(regtop_g_udb1_r[1]),
	.b(n246073));
   na02f02 U266189 (.o(n246066),
	.a(n246064),
	.b(n246063));
   in01f01 U266190 (.o(n246160),
	.a(n246065));
   na02f01 U266191 (.o(n246159),
	.a(n246066),
	.b(regtop_g_udb2_r[1]));
   in01f01 U266192 (.o(n246067),
	.a(n246159));
   na02f10 U266193 (.o(n246076),
	.a(regtop_g_udb1_r[2]),
	.b(regtop_g_udb2_r[2]));
   na02f02 U266194 (.o(n246070),
	.a(n246069),
	.b(n246068));
   na02f03 U266195 (.o(n246075),
	.a(n246072),
	.b(n246071));
   no02f03 U266196 (.o(n246173),
	.a(n246075),
	.b(n246074));
   na02f03 U266197 (.o(n246174),
	.a(n246075),
	.b(n246074));
   in01f01 U266199 (.o(n246079),
	.a(n246076));
   na02f02 U266200 (.o(n246082),
	.a(regtop_g_udb1_r[3]),
	.b(n246088));
   na02f02 U266201 (.o(n246081),
	.a(regtop_g_udb2_r[3]),
	.b(n246088));
   na02f02 U266202 (.o(n246083),
	.a(n246082),
	.b(n246081));
   na02f03 U266203 (.o(n246089),
	.a(regtop_g_udb0_r[3]),
	.b(n246083));
   na02f01 U266204 (.o(n246085),
	.a(n246083),
	.b(n246089));
   na02f01 U266205 (.o(n246084),
	.a(regtop_g_udb0_r[3]),
	.b(n246089));
   na02f02 U266206 (.o(n246086),
	.a(n246085),
	.b(n246084));
   no02f03 U266207 (.o(n246151),
	.a(n246087),
	.b(n246086));
   oa12f01 U266208 (.o(n246101),
	.a(n246152),
	.b(n246156),
	.c(n246151));
   no02m02 U266209 (.o(n246092),
	.a(n246091),
	.b(n246090));
   na02f03 U266210 (.o(n246111),
	.a(regtop_g_udb0_r[4]),
	.b(regtop_g_udb1_r[4]));
   na02m02 U266211 (.o(n246094),
	.a(n246111),
	.b(regtop_g_udb1_r[4]));
   na02m02 U266212 (.o(n246093),
	.a(n246111),
	.b(regtop_g_udb0_r[4]));
   na02f02 U266213 (.o(n246095),
	.a(n246094),
	.b(n246093));
   no02f04 U266214 (.o(n246107),
	.a(n246099),
	.b(n246098));
   no02f04 U266215 (.o(n246110),
	.a(n246107),
	.b(n246151));
   in01s01 U266218 (.o(n246114),
	.a(n246111));
   na02f01 U266219 (.o(n246117),
	.a(regtop_g_udb0_r[5]),
	.b(n246123));
   na02f01 U266220 (.o(n246116),
	.a(regtop_g_udb1_r[5]),
	.b(n246123));
   na02f02 U266221 (.o(n246118),
	.a(n246117),
	.b(n246116));
   na02f02 U266222 (.o(n246124),
	.a(regtop_g_udb2_r[5]),
	.b(n246118));
   oa12f02 U266223 (.o(n246138),
	.a(n246144),
	.b(n246146),
	.c(n246143));
   in01s01 U266224 (.o(n246126),
	.a(n246123));
   in01f01 U266225 (.o(n246125),
	.a(n246124));
   in01f01 U266226 (.o(n246924),
	.a(regtop_g_udb0_r[6]));
   no02f02 U266227 (.o(n246139),
	.a(n246138),
	.b(n246140));
   no02f02 U266228 (.o(n246142),
	.a(n246138),
	.b(n246139));
   no02f02 U266229 (.o(n246141),
	.a(n246140),
	.b(n246139));
   no02f03 U266230 (.o(n249042),
	.a(n246142),
	.b(n246141));
   na02f02 U266231 (.o(n246147),
	.a(n246146),
	.b(n246148));
   na02f01 U266232 (.o(n246150),
	.a(n246146),
	.b(n246147));
   na02f01 U266233 (.o(n246149),
	.a(n246148),
	.b(n246147));
   na02f03 U266234 (.o(n249036),
	.a(n246150),
	.b(n246149));
   in01f02 U266235 (.o(n246183),
	.a(n249036));
   in01f01 U266236 (.o(n246153),
	.a(n246151));
   na02m02 U266237 (.o(n246154),
	.a(n246153),
	.b(n246152));
   na02m02 U266238 (.o(n246155),
	.a(n246154),
	.b(n246156));
   in01f01 U266239 (.o(n246182),
	.a(n248990));
   in01s01 U266240 (.o(n246168),
	.a(n246166));
   in01f01 U266241 (.o(n246175),
	.a(n246173));
   na02f01 U266242 (.o(n246177),
	.a(n246176),
	.b(n246178));
   na02f01 U266243 (.o(n246180),
	.a(n246176),
	.b(n246177));
   na02f01 U266244 (.o(n246179),
	.a(n246178),
	.b(n246177));
   na02f02 U266245 (.o(n248984),
	.a(n246180),
	.b(n246179));
   na02f04 U266246 (.o(n246181),
	.a(n248952),
	.b(n248984));
   no02f10 U266247 (.o(n249066),
	.a(n246904),
	.b(n246189));
   na02s01 U266248 (.o(n246190),
	.a(regtop_g_adb_r[5]),
	.b(regtop_g_adb_r[3]));
   in01s01 U266249 (.o(n246191),
	.a(n246190));
   in01s01 U266250 (.o(n246195),
	.a(n246194));
   na02s01 U266251 (.o(n246207),
	.a(y1_bs_data_r[7]),
	.b(busiftop_vmem_ch_r));
   in01s01 U266252 (.o(n244245),
	.a(n246207));
   in01s01 U266253 (.o(n212679),
	.a(n246208));
   in01s01 U266254 (.o(n244263),
	.a(n246209));
   in01s01 U266255 (.o(n244262),
	.a(n246210));
   in01s01 U266256 (.o(n244250),
	.a(n246211));
   no02s01 U266257 (.o(n212573),
	.a(n246726),
	.b(FE_OFN68_n247591));
   in01s01 U266258 (.o(n246215),
	.a(busrtop_b_rreq_vrh_cnt_16byte_r[1]));
   na02s01 U266259 (.o(n246212),
	.a(busrtop_b_rreq_vrh_cnt_16byte_r[1]),
	.b(busrtop_b_rreq_vrh_cnt_16byte_r[0]));
   oa22s01 U266260 (.o(n170938),
	.a(n246229),
	.b(n253125),
	.c(busiftop_status_b_current_0_),
	.d(n246215));
   in01f01 U266261 (.o(n246964),
	.a(n246370));
   na02s01 U266262 (.o(n246216),
	.a(n249064),
	.b(vldtop_vld_syndec_vld_seqhed_pre_SHIFT[1]));
   na02s01 U266263 (.o(n212415),
	.a(n246218),
	.b(n246216));
   na02s01 U266264 (.o(n246217),
	.a(n249064),
	.b(vldtop_vld_syndec_vld_seqhed_pre_SHIFT[4]));
   na02s01 U266265 (.o(n212416),
	.a(n246218),
	.b(n246217));
   na02s01 U266266 (.o(n246219),
	.a(FE_OFN2_g_swrst_r_n),
	.b(vldtop_vld_syndec_vld_vscdet_v_search_1st_r));
   in01s01 U266267 (.o(n246224),
	.a(n246219));
   na02s01 U266268 (.o(n212486),
	.a(n246224),
	.b(n246220));
   in01s01 U266269 (.o(n246221),
	.a(vldtop_vld_syndec_vld_vscdet_v_detvald_r[0]));
   na02s01 U266270 (.o(n246222),
	.a(n246779),
	.b(n246221));
   oa12s01 U266271 (.o(n246223),
	.a(n246222),
	.b(n246779),
	.c(n248999));
   na02s01 U266272 (.o(n212487),
	.a(n246224),
	.b(n246223));
   in01s01 U266273 (.o(n246227),
	.a(regtop_g_ari_r[3]));
   na02s01 U266274 (.o(n246226),
	.a(regtop_g_paramdata_r[24]),
	.b(FE_OFN220_n246261));
   oa12s01 U266275 (.o(n212140),
	.a(n246226),
	.b(FE_OFN220_n246261),
	.c(n246227));
   in01s01 U266276 (.o(n253038),
	.a(busrtop_b_rreq_vrh_add1_r[0]));
   na02s01 U266277 (.o(n246228),
	.a(n253125),
	.b(vh_1_ph_add[0]));
   in01s01 U266278 (.o(n246232),
	.a(n246228));
   no02s01 U266279 (.o(n246231),
	.a(n249913),
	.b(n253038));
   no02s01 U266280 (.o(n246236),
	.a(n246232),
	.b(n246231));
   na02s01 U266281 (.o(n246235),
	.a(n249916),
	.b(n245811));
   na02s01 U266282 (.o(n157840),
	.a(n246236),
	.b(n246235));
   no02s01 U266283 (.o(n212571),
	.a(n246786),
	.b(FE_OFN68_n247591));
   na02s01 U266284 (.o(n246239),
	.a(regtop_g_atscd_r[29]),
	.b(n246247));
   oa12s01 U266285 (.o(n212118),
	.a(n246239),
	.b(n246247),
	.c(n252666));
   na02s01 U266286 (.o(n246240),
	.a(regtop_g_atscd_r[25]),
	.b(n246247));
   oa12s01 U266287 (.o(n212114),
	.a(n246240),
	.b(n246247),
	.c(n252658));
   na02s01 U266288 (.o(n246241),
	.a(regtop_g_atscd_r[26]),
	.b(n246247));
   oa12s01 U266289 (.o(n212115),
	.a(n246241),
	.b(n246247),
	.c(n252660));
   na02s01 U266290 (.o(n246242),
	.a(regtop_g_atscd_r[31]),
	.b(n246247));
   oa12s01 U266291 (.o(n212120),
	.a(n246242),
	.b(n246247),
	.c(n252755));
   na02s01 U266292 (.o(n246243),
	.a(regtop_g_atscd_r[30]),
	.b(n246247));
   oa12s01 U266293 (.o(n212119),
	.a(n246243),
	.b(n246247),
	.c(n252778));
   na02s01 U266294 (.o(n246244),
	.a(regtop_g_atscd_r[27]),
	.b(n246247));
   oa12s01 U266295 (.o(n212116),
	.a(n246244),
	.b(n246247),
	.c(n252662));
   na02s01 U266296 (.o(n246245),
	.a(regtop_g_atscd_r[24]),
	.b(n246247));
   oa12s01 U266297 (.o(n212113),
	.a(n246245),
	.b(n246247),
	.c(n252656));
   na02s01 U266298 (.o(n246246),
	.a(regtop_g_atscd_r[28]),
	.b(n246247));
   oa12s01 U266299 (.o(n212117),
	.a(n246246),
	.b(n246247),
	.c(n252664));
   na02s01 U266300 (.o(n246249),
	.a(n246260),
	.b(regtop_g_ari_r[0]));
   na02s01 U266301 (.o(n246248),
	.a(regtop_g_paramdata_r[21]),
	.b(FE_OFN220_n246261));
   na02s01 U266302 (.o(n212139),
	.a(n246249),
	.b(n246248));
   na02s01 U266303 (.o(n246251),
	.a(n246260),
	.b(regtop_g_ari_r[2]));
   na02s01 U266304 (.o(n246250),
	.a(regtop_g_paramdata_r[23]),
	.b(FE_OFN220_n246261));
   na02s01 U266305 (.o(n212141),
	.a(n246251),
	.b(n246250));
   na02s01 U266306 (.o(n246253),
	.a(n246260),
	.b(regtop_g_frc_r[1]));
   na02s01 U266307 (.o(n246252),
	.a(regtop_g_paramdata_r[18]),
	.b(FE_OFN220_n246261));
   na02s01 U266308 (.o(n212143),
	.a(n246253),
	.b(n246252));
   na02s01 U266309 (.o(n246255),
	.a(n246260),
	.b(regtop_g_frc_r[0]));
   na02s01 U266310 (.o(n246254),
	.a(regtop_g_paramdata_r[17]),
	.b(FE_OFN220_n246261));
   na02s01 U266311 (.o(n212146),
	.a(n246255),
	.b(n246254));
   na02s01 U266312 (.o(n246257),
	.a(n246260),
	.b(regtop_g_ari_r[1]));
   na02s01 U266313 (.o(n246256),
	.a(regtop_g_paramdata_r[22]),
	.b(FE_OFN220_n246261));
   na02s01 U266314 (.o(n246259),
	.a(n246260),
	.b(regtop_g_frc_r[3]));
   na02s01 U266315 (.o(n246258),
	.a(regtop_g_paramdata_r[20]),
	.b(FE_OFN220_n246261));
   na02s01 U266316 (.o(n212145),
	.a(n246259),
	.b(n246258));
   na02s01 U266317 (.o(n246263),
	.a(n246260),
	.b(regtop_g_frc_r[2]));
   na02s01 U266318 (.o(n246262),
	.a(regtop_g_paramdata_r[19]),
	.b(FE_OFN220_n246261));
   na02s01 U266319 (.o(n212144),
	.a(n246263),
	.b(n246262));
   ao22s01 U266320 (.o(n246264),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[4]),
	.c(n245940),
	.d(regtop_g_vsv_r[3]));
   in01s01 U266321 (.o(n211931),
	.a(n246264));
   ao22s01 U266322 (.o(n246265),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[2]),
	.c(FE_OFN486_n245940),
	.d(regtop_g_vsv_r[1]));
   in01s01 U266323 (.o(n211929),
	.a(n246265));
   ao22s01 U266324 (.o(n246267),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[3]),
	.c(FE_OFN486_n245940),
	.d(regtop_g_vsv_r[2]));
   in01s01 U266325 (.o(n211930),
	.a(n246267));
   oa22s01 U266326 (.o(n246268),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[27]),
	.b(vldtop_vld_syndec_ADP[1]),
	.c(vldtop_vld_syndec_vld_vlfeed_lower[25]),
	.d(n246419));
   in01s01 U266327 (.o(n246698),
	.a(n246268));
   oa22s01 U266328 (.o(n246399),
	.a(n246707),
	.b(n246695),
	.c(n246698),
	.d(n246693));
   no02s01 U266329 (.o(n246391),
	.a(n246696),
	.b(n246527));
   no02s01 U266330 (.o(n246269),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246391));
   na02s01 U266331 (.o(n246392),
	.a(n246565),
	.b(n246699));
   na02s01 U266332 (.o(n246270),
	.a(n246269),
	.b(n246392));
   no02s01 U266333 (.o(n246279),
	.a(n246399),
	.b(n246270));
   in01f01 U266334 (.o(n246512),
	.a(n246466));
   oa22s01 U266335 (.o(n246271),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[23]),
	.b(vldtop_vld_syndec_ADP[1]),
	.c(vldtop_vld_syndec_vld_vlfeed_lower[21]),
	.d(n246419));
   in01f01 U266336 (.o(n246511),
	.a(n246464));
   oa22s01 U266337 (.o(n246272),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[19]),
	.b(vldtop_vld_syndec_ADP[1]),
	.c(vldtop_vld_syndec_vld_vlfeed_lower[17]),
	.d(n246419));
   in01s01 U266338 (.o(n246514),
	.a(n246272));
   ao22s01 U266339 (.o(n246277),
	.a(n246512),
	.b(n246694),
	.c(n246511),
	.d(n246514));
   na02f02 U266340 (.o(n246485),
	.a(n246565),
	.b(vldtop_vld_syndec_ADP[4]));
   in01s01 U266341 (.o(n246516),
	.a(n246485));
   in01s01 U266342 (.o(n246304),
	.a(n246273));
   ao22s01 U266343 (.o(n246274),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(vldtop_vld_syndec_vld_vlfeed_lower[9]),
	.c(n246419),
	.d(vldtop_vld_syndec_vld_vlfeed_lower[11]));
   in01s01 U266344 (.o(n246275),
	.a(n246274));
   na02s01 U266345 (.o(n246278),
	.a(n246277),
	.b(n246276));
   no02s01 U266346 (.o(n246280),
	.a(n246279),
	.b(n246278));
   in01s01 U266347 (.o(n246281),
	.a(n246280));
   na02s01 U266348 (.o(n246282),
	.a(g_swrst_r_n),
	.b(n246281));
   in01s01 U266349 (.o(vldtop_vld_syndec_vld_outbuf_N463),
	.a(n246282));
   in01s01 U266350 (.o(n246283),
	.a(vldtop_vld_syndec_UREG[27]));
   na02s01 U266351 (.o(n246284),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n246283));
   ao22f01 U266352 (.o(n246287),
	.a(vldtop_vld_syndec_ADP[2]),
	.b(n246285),
	.c(n246692),
	.d(n246284));
   oa12s01 U266353 (.o(n246286),
	.a(n246659),
	.b(vldtop_vld_syndec_UREG[29]),
	.c(n246684));
   no02s01 U266354 (.o(n246296),
	.a(n246287),
	.b(n246286));
   in01s01 U266355 (.o(n246294),
	.a(n246337));
   na02s01 U266356 (.o(n246288),
	.a(vldtop_vld_syndec_ADP[3]),
	.b(n246670));
   no02f01 U266357 (.o(n246291),
	.a(n246692),
	.b(n246288));
   in01s01 U266358 (.o(n246290),
	.a(n246289));
   na02s01 U266359 (.o(n246292),
	.a(n246291),
	.b(n246290));
   oa22f01 U266360 (.o(n246295),
	.a(n246294),
	.b(n246711),
	.c(n246293),
	.d(n246292));
   no02s01 U266361 (.o(n246459),
	.a(n246297),
	.b(n246697));
   na02s01 U266362 (.o(n246298),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246457));
   no02s01 U266363 (.o(n246299),
	.a(n246459),
	.b(n246298));
   na02s01 U266364 (.o(n246300),
	.a(g_swrst_r_n),
	.b(n246885));
   in01s01 U266365 (.o(vldtop_vld_syndec_vld_outbuf_N485),
	.a(n246300));
   no02s01 U266366 (.o(vldtop_vld_syndec_vld_outbuf_N480),
	.a(n246301),
	.b(FE_OFN68_n247591));
   in01s01 U266367 (.o(n246310),
	.a(n246988));
   na02s01 U266368 (.o(n246311),
	.a(g_swrst_r_n),
	.b(n246310));
   in01s01 U266369 (.o(vldtop_vld_syndec_vld_outbuf_N467),
	.a(n246311));
   in01s01 U266370 (.o(n247293),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[23]));
   in01s01 U266371 (.o(n247131),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[25]));
   ao22s01 U266372 (.o(n246315),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n247293),
	.c(n246419),
	.d(n247131));
   ao22s01 U266373 (.o(n246319),
	.a(n246700),
	.b(n246465),
	.c(n246565),
	.d(n246463));
   in01s01 U266374 (.o(n247364),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[19]));
   in01s01 U266375 (.o(n247127),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[21]));
   ao22s01 U266376 (.o(n246316),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n247364),
	.c(n246419),
	.d(n247127));
   in01s01 U266377 (.o(n246467),
	.a(n246316));
   na02s01 U266378 (.o(n246318),
	.a(n246570),
	.b(n246467));
   na02s01 U266379 (.o(n246317),
	.a(n246568),
	.b(n246345));
   na02s01 U266380 (.o(n246322),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n246982));
   in01s01 U266381 (.o(vldtop_vld_syndec_vld_outbuf_N473),
	.a(n246322));
   ao22f01 U266382 (.o(n246480),
	.a(n246700),
	.b(n246536),
	.c(n246570),
	.d(n246524));
   in01s01 U266383 (.o(n246323),
	.a(n246535));
   no02f01 U266384 (.o(n246477),
	.a(n246323),
	.b(n246695));
   no02f01 U266385 (.o(n246476),
	.a(n246430),
	.b(n246697));
   na02s01 U266386 (.o(n246335),
	.a(n246570),
	.b(n246533));
   na02s01 U266387 (.o(n246334),
	.a(n246565),
	.b(n246435));
   no02s01 U266388 (.o(n246326),
	.a(n246419),
	.b(n246325));
   no02s01 U266389 (.o(n246332),
	.a(vldtop_vld_syndec_ADP[2]),
	.b(n246326));
   no02s01 U266390 (.o(n246331),
	.a(n246692),
	.b(n246327));
   in01s01 U266391 (.o(n246328),
	.a(vldtop_vld_syndec_UREG[28]));
   no02s01 U266392 (.o(n246329),
	.a(n246684),
	.b(n246328));
   no02s01 U266393 (.o(n246330),
	.a(vldtop_vld_syndec_ADP[3]),
	.b(n246329));
   oa12f01 U266394 (.o(n246333),
	.a(n246330),
	.b(n246332),
	.c(n246331));
   na02s01 U266395 (.o(n246336),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n246884));
   ao22s01 U266396 (.o(n246348),
	.a(n246568),
	.b(n246344),
	.c(n246565),
	.d(n246465));
   na02s01 U266397 (.o(n246346),
	.a(n246700),
	.b(n246345));
   na02s01 U266398 (.o(n246351),
	.a(g_swrst_r_n),
	.b(n246997));
   in01s01 U266399 (.o(vldtop_vld_syndec_vld_outbuf_N477),
	.a(n246351));
   no02s01 U266400 (.o(n246352),
	.a(vldtop_vld_syndec_vld_vlfeed_feed_on),
	.b(FE_OFN68_n247591));
   no03f02 U266401 (.o(n246358),
	.a(vldtop_vld_syndec_UREG[21]),
	.b(vldtop_vld_syndec_UREG[18]),
	.c(vldtop_vld_syndec_UREG[19]));
   no04f02 U266402 (.o(n246357),
	.a(vldtop_vld_syndec_UREG[22]),
	.b(vldtop_vld_syndec_UREG[23]),
	.c(vldtop_vld_syndec_UREG[17]),
	.d(vldtop_vld_syndec_UREG[20]));
   no04f04 U266403 (.o(n246360),
	.a(vldtop_vld_syndec_UREG[24]),
	.b(n246359),
	.c(n246785),
	.d(n249005));
   in01s01 U266404 (.o(n246367),
	.a(n246366));
   no02s01 U266405 (.o(n246368),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n246367));
   in01s01 U266406 (.o(n246369),
	.a(n246368));
   na02s01 U266407 (.o(n246371),
	.a(n246805),
	.b(n246369));
   oa22s01 U266408 (.o(n212579),
	.a(n246838),
	.b(n246419),
	.c(n246371),
	.d(n246836));
   in01s01 U266409 (.o(n246376),
	.a(g_line_offset_r));
   no02s01 U266410 (.o(n249717),
	.a(n246372),
	.b(n249720));
   na02s01 U266411 (.o(n246373),
	.a(n253015),
	.b(n249717));
   in01s01 U266412 (.o(n246375),
	.a(n246373));
   na02s01 U266413 (.o(n246374),
	.a(regtop_g_wd_r[0]),
	.b(n246375));
   oa12s01 U266414 (.o(n212788),
	.a(n246374),
	.b(n246376),
	.c(n246375));
   no02s01 U266415 (.o(n246378),
	.a(n246377),
	.b(n246695));
   no02s01 U266416 (.o(n246389),
	.a(n246553),
	.b(n246378));
   no02s01 U266417 (.o(n246552),
	.a(n246379),
	.b(n246527));
   no02s01 U266418 (.o(n246551),
	.a(n246380),
	.b(n246697));
   in01f02 U266419 (.o(n247368),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[24]));
   in01s01 U266420 (.o(n246569),
	.a(n246381));
   oa22s01 U266421 (.o(n246385),
	.a(n246466),
	.b(n246564),
	.c(n246464),
	.d(n246569));
   in01f01 U266422 (.o(n247173),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[20]));
   in01f01 U266423 (.o(n247276),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[22]));
   ao22s01 U266424 (.o(n246382),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n247173),
	.c(n246419),
	.d(n247276));
   in01s01 U266425 (.o(n246497),
	.a(n246382));
   ao22s01 U266428 (.o(n246383),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(FE_OFN525_vldtop_vld_syndec_vld_vlfeed_lower_16_),
	.c(n246419),
	.d(FE_OFN537_vldtop_vld_syndec_vld_vlfeed_lower_18_));
   in01s01 U266429 (.o(n246407),
	.a(n246383));
   oa22s01 U266430 (.o(n246384),
	.a(n246485),
	.b(n246497),
	.c(n246484),
	.d(n246407));
   no02s01 U266431 (.o(n246386),
	.a(n246385),
	.b(n246384));
   in01s01 U266432 (.o(n246387),
	.a(n246386));
   in01s01 U266433 (.o(n246974),
	.a(n246985));
   na02s01 U266434 (.o(n246390),
	.a(g_swrst_r_n),
	.b(n246974));
   in01s01 U266435 (.o(vldtop_vld_syndec_vld_outbuf_N470),
	.a(n246390));
   no02s01 U266436 (.o(n246393),
	.a(n246391),
	.b(n246670));
   na02s01 U266437 (.o(n246398),
	.a(n246393),
	.b(n246392));
   oa22s01 U266438 (.o(n246395),
	.a(n246712),
	.b(n246578),
	.c(n246715),
	.d(n246711));
   na02s01 U266439 (.o(n246400),
	.a(g_swrst_r_n),
	.b(n247017));
   in01s01 U266440 (.o(vldtop_vld_syndec_vld_outbuf_N479),
	.a(n246400));
   no02s01 U266441 (.o(n246412),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246404));
   ao22s01 U266444 (.o(n246405),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(FE_OFN540_vldtop_vld_syndec_vld_vlfeed_lower_12_),
	.c(n246419),
	.d(FE_OFN530_vldtop_vld_syndec_vld_vlfeed_lower_14_));
   in01s01 U266445 (.o(n246406),
	.a(n246405));
   oa22s01 U266446 (.o(n246408),
	.a(vldtop_vld_syndec_ADP[2]),
	.b(n246407),
	.c(n246406),
	.d(n246692));
   ao12f01 U266447 (.o(n246411),
	.a(n246670),
	.b(vldtop_vld_syndec_ADP[3]),
	.c(n246408));
   oa22s01 U266448 (.o(n246409),
	.a(n246466),
	.b(n246569),
	.c(n246464),
	.d(n246497));
   in01s01 U266449 (.o(n246410),
	.a(n246409));
   na02s01 U266450 (.o(n246413),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n246987));
   in01s01 U266451 (.o(vldtop_vld_syndec_vld_outbuf_N466),
	.a(n246413));
   in01s01 U266452 (.o(n246418),
	.a(n246414));
   na02s01 U266453 (.o(n246416),
	.a(n246670),
	.b(n246415));
   ao22f02 U266454 (.o(n246526),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n247276),
	.c(n246419),
	.d(n247368));
   ao22s01 U266455 (.o(n246482),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(FE_OFN537_vldtop_vld_syndec_vld_vlfeed_lower_18_),
	.c(n246419),
	.d(n247173));
   ao22s01 U266456 (.o(n246420),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(FE_OFN530_vldtop_vld_syndec_vld_vlfeed_lower_14_),
	.c(n246419),
	.d(FE_OFN525_vldtop_vld_syndec_vld_vlfeed_lower_16_));
   in01s01 U266457 (.o(n246483),
	.a(n246420));
   in01f01 U266458 (.o(n247222),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[10]));
   ao22s01 U266459 (.o(n246421),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(n247222),
	.c(n246419),
	.d(FE_OFN540_vldtop_vld_syndec_vld_vlfeed_lower_12_));
   in01s01 U266460 (.o(n246422),
	.a(n246421));
   in01s01 U266461 (.o(n246428),
	.a(n247007));
   in01s01 U266462 (.o(vldtop_vld_syndec_vld_outbuf_N464),
	.a(n246429));
   in01s01 U266463 (.o(n246534),
	.a(n246430));
   no02s01 U266464 (.o(n246432),
	.a(n246695),
	.b(n246534));
   no02s01 U266465 (.o(n246431),
	.a(n246527),
	.b(n246524));
   oa12s01 U266466 (.o(n246442),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246432),
	.c(n246431));
   ao22s01 U266467 (.o(n246434),
	.a(n246526),
	.b(vldtop_vld_syndec_ADP[2]),
	.c(n246528),
	.d(n246692));
   na02s01 U266468 (.o(n246433),
	.a(vldtop_vld_syndec_ADP[3]),
	.b(vldtop_vld_syndec_ADP[4]));
   na02f01 U266469 (.o(n246443),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n246998));
   in01s01 U266470 (.o(vldtop_vld_syndec_vld_outbuf_N476),
	.a(n246443));
   ao22s01 U266471 (.o(n246468),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(vldtop_vld_syndec_vld_vlfeed_lower[15]),
	.c(n246419),
	.d(vldtop_vld_syndec_vld_vlfeed_lower[17]));
   ao22s01 U266472 (.o(n246450),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(vldtop_vld_syndec_vld_vlfeed_lower[11]),
	.c(n246419),
	.d(vldtop_vld_syndec_vld_vlfeed_lower[13]));
   na02s01 U266473 (.o(n246456),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n246981));
   in01s01 U266474 (.o(vldtop_vld_syndec_vld_outbuf_N465),
	.a(n246456));
   na02s01 U266475 (.o(n246458),
	.a(n246670),
	.b(n246457));
   in01s01 U266476 (.o(n246473),
	.a(n246462));
   no02s01 U266477 (.o(n246471),
	.a(n246470),
	.b(n246469));
   in01s01 U266478 (.o(n246472),
	.a(n246471));
   in01s01 U266479 (.o(n246474),
	.a(n246989));
   na02s01 U266480 (.o(n246475),
	.a(g_swrst_r_n),
	.b(n246474));
   no02s01 U266481 (.o(n246479),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246476));
   in01s01 U266482 (.o(n246478),
	.a(n246477));
   in01s01 U266483 (.o(n246490),
	.a(n246481));
   in01s01 U266484 (.o(n246525),
	.a(n246482));
   in01s01 U266485 (.o(n246487),
	.a(n246486));
   in01s01 U266486 (.o(n246971),
	.a(n246984));
   na02s01 U266487 (.o(n246491),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n246971));
   in01s01 U266488 (.o(vldtop_vld_syndec_vld_outbuf_N468),
	.a(n246491));
   in01s01 U266489 (.o(n246574),
	.a(n246492));
   oa22s01 U266490 (.o(n246494),
	.a(n246578),
	.b(n246567),
	.c(n246708),
	.d(n246574));
   no02s01 U266491 (.o(n246505),
	.a(n246494),
	.b(n246493));
   na02s01 U266492 (.o(n246496),
	.a(n246565),
	.b(n246569));
   na02s01 U266493 (.o(n246495),
	.a(n246700),
	.b(n246564));
   na02s01 U266494 (.o(n246502),
	.a(n246496),
	.b(n246495));
   na02s01 U266495 (.o(n246500),
	.a(n246570),
	.b(n246497));
   in01s01 U266496 (.o(n246571),
	.a(n246498));
   na02s01 U266497 (.o(n246501),
	.a(n246500),
	.b(n246499));
   no02s01 U266498 (.o(n246503),
	.a(n246502),
	.b(n246501));
   na02s01 U266499 (.o(n246506),
	.a(g_swrst_r_n),
	.b(n246991));
   in01s01 U266500 (.o(vldtop_vld_syndec_vld_outbuf_N474),
	.a(n246506));
   na02s01 U266501 (.o(n246674),
	.a(n246700),
	.b(n246712));
   in01s01 U266502 (.o(n246510),
	.a(n246674));
   no02s01 U266503 (.o(n246671),
	.a(n246696),
	.b(n246693));
   na02s01 U266504 (.o(n246673),
	.a(n246568),
	.b(n246715));
   in01s01 U266505 (.o(n246509),
	.a(n246673));
   in01s01 U266506 (.o(n246507),
	.a(n246707));
   na02s01 U266507 (.o(n246672),
	.a(n246565),
	.b(n246507));
   in01s01 U266508 (.o(n246508),
	.a(n246672));
   in01s01 U266509 (.o(n246513),
	.a(n246699));
   na02s01 U266510 (.o(n246519),
	.a(n246518),
	.b(n246517));
   in01s01 U266511 (.o(n246521),
	.a(n246994));
   na02s01 U266512 (.o(n246522),
	.a(g_swrst_r_n),
	.b(n246521));
   in01s01 U266513 (.o(vldtop_vld_syndec_vld_outbuf_N471),
	.a(n246522));
   na02s01 U266514 (.o(n246523),
	.a(g_swrst_r_n),
	.b(n247002));
   in01s01 U266515 (.o(vldtop_vld_syndec_vld_outbuf_N483),
	.a(n246523));
   ao22s01 U266516 (.o(n246532),
	.a(n246570),
	.b(n246525),
	.c(n246568),
	.d(n246524));
   no02s01 U266517 (.o(n246530),
	.a(n246526),
	.b(n246697));
   no02s01 U266518 (.o(n246529),
	.a(n246528),
	.b(n246527));
   na02s01 U266519 (.o(n246541),
	.a(g_swrst_r_n),
	.b(n246980));
   in01s01 U266520 (.o(vldtop_vld_syndec_vld_outbuf_N472),
	.a(n246541));
   na02s01 U266521 (.o(n246542),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(vldtop_vld_syndec_UREG[28]));
   no02s01 U266522 (.o(n246550),
	.a(n246542),
	.b(n246708));
   no02s01 U266523 (.o(n246549),
	.a(n246544),
	.b(n246714));
   na02s01 U266524 (.o(n246545),
	.a(vldtop_vld_syndec_UREG[30]),
	.b(n246659));
   no02s01 U266525 (.o(n246548),
	.a(n246684),
	.b(n246545));
   in01s01 U266526 (.o(n246575),
	.a(n246546));
   oa22s01 U266527 (.o(n246547),
	.a(n246575),
	.b(n246711),
	.c(n246578),
	.d(n246574));
   no04s02 U266528 (.o(n246562),
	.a(n246550),
	.b(n246549),
	.c(n246548),
	.d(n246547));
   no02s01 U266529 (.o(n246560),
	.a(n246552),
	.b(n246551));
   in01s01 U266530 (.o(n246559),
	.a(n246553));
   na02s01 U266531 (.o(n246557),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246554));
   in01s01 U266532 (.o(n246556),
	.a(n246555));
   oa22s01 U266533 (.o(n246558),
	.a(n246568),
	.b(n246670),
	.c(n246557),
	.d(n246556));
   na03s01 U266534 (.o(n246561),
	.a(n246560),
	.b(n246559),
	.c(n246558));
   na02s01 U266535 (.o(n246563),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247018));
   in01s01 U266536 (.o(vldtop_vld_syndec_vld_outbuf_N486),
	.a(n246563));
   na02s01 U266537 (.o(n246566),
	.a(n246565),
	.b(n246564));
   na02s01 U266538 (.o(n246583),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246566));
   na02s01 U266539 (.o(n246572),
	.a(n246700),
	.b(n246571));
   oa22s01 U266540 (.o(n246579),
	.a(n246578),
	.b(n246577),
	.c(n246711),
	.d(n246576));
   oa12f02 U266541 (.o(n247009),
	.a(n246581),
	.b(n246583),
	.c(n246582));
   in01s01 U266542 (.o(vldtop_vld_syndec_vld_outbuf_N478),
	.a(n246584));
   in01s01 U266543 (.o(n211934),
	.a(n246586));
   ao22s01 U266544 (.o(n246587),
	.a(FE_OFN366_n246266),
	.b(regtop_g_paramdata_r[1]),
	.c(FE_OFN486_n245940),
	.d(regtop_g_vsv_r[0]));
   in01s01 U266545 (.o(n211921),
	.a(n246588));
   in01s01 U266546 (.o(n211919),
	.a(n246589));
   in01s01 U266547 (.o(n211918),
	.a(n246590));
   in01s01 U266548 (.o(n211932),
	.a(n246591));
   in01s01 U266549 (.o(n211922),
	.a(n246592));
   in01s01 U266550 (.o(n211935),
	.a(n246593));
   in01s01 U266551 (.o(n211920),
	.a(n246594));
   in01s01 U266552 (.o(n211917),
	.a(n246595));
   in01s01 U266553 (.o(n211933),
	.a(n246596));
   in01s01 U266554 (.o(n211938),
	.a(n246597));
   in01s01 U266555 (.o(n211928),
	.a(n246598));
   in01s01 U266556 (.o(n211939),
	.a(n246599));
   in01s01 U266557 (.o(n211927),
	.a(n246600));
   in01s01 U266558 (.o(n211926),
	.a(n246601));
   ao22s01 U266559 (.o(n246602),
	.a(regtop_g_paramdata_r[17]),
	.b(FE_OFN366_n246266),
	.c(FE_OFN486_n245940),
	.d(regtop_g_hsv_r[4]));
   in01s01 U266560 (.o(n211924),
	.a(n246603));
   in01s01 U266561 (.o(n211936),
	.a(n246604));
   in01s01 U266562 (.o(n211923),
	.a(n246606));
   in01s01 U266563 (.o(n246615),
	.a(regtop_g_usrd_r[16]));
   in01s01 U266565 (.o(n246617),
	.a(n249137));
   na02s01 U266566 (.o(n246619),
	.a(regtop_g_paramdata_r[17]),
	.b(n246647));
   na02s01 U266567 (.o(n212271),
	.a(n246620),
	.b(n246619));
   na02s01 U266570 (.o(n246623),
	.a(regtop_g_paramdata_r[18]),
	.b(n246647));
   na02s01 U266571 (.o(n212272),
	.a(n246624),
	.b(n246623));
   in01s01 U266572 (.o(n246625),
	.a(regtop_g_usrd_r[23]));
   na02s01 U266575 (.o(n246627),
	.a(regtop_g_paramdata_r[24]),
	.b(n246647));
   na02s01 U266576 (.o(n212278),
	.a(n246628),
	.b(n246627));
   in01s01 U266577 (.o(n246629),
	.a(regtop_g_usrd_r[18]));
   na02s01 U266580 (.o(n246631),
	.a(regtop_g_paramdata_r[19]),
	.b(n246647));
   na02s01 U266581 (.o(n212273),
	.a(n246632),
	.b(n246631));
   in01s01 U266582 (.o(n246633),
	.a(regtop_g_usrd_r[22]));
   na02s01 U266585 (.o(n246635),
	.a(regtop_g_paramdata_r[23]),
	.b(n246647));
   in01s01 U266586 (.o(n246637),
	.a(regtop_g_usrd_r[19]));
   oa22s01 U266587 (.o(n246638),
	.a(FE_OFN6_n246618),
	.b(n246637),
	.c(n246637),
	.d(n249079));
   in01s01 U266588 (.o(n246640),
	.a(n246638));
   na02s01 U266589 (.o(n246639),
	.a(regtop_g_paramdata_r[20]),
	.b(n246647));
   na02s01 U266590 (.o(n212274),
	.a(n246640),
	.b(n246639));
   in01s01 U266591 (.o(n246641),
	.a(regtop_g_usrd_r[21]));
   oa22s01 U266592 (.o(n246642),
	.a(FE_OFN6_n246618),
	.b(n246641),
	.c(n246641),
	.d(n249079));
   in01s01 U266593 (.o(n246644),
	.a(n246642));
   na02s01 U266594 (.o(n246643),
	.a(regtop_g_paramdata_r[22]),
	.b(n246647));
   na02s01 U266595 (.o(n212276),
	.a(n246644),
	.b(n246643));
   in01s01 U266596 (.o(n246645),
	.a(regtop_g_usrd_r[20]));
   oa22s01 U266597 (.o(n246646),
	.a(FE_OFN6_n246618),
	.b(n246645),
	.c(n246645),
	.d(n249079));
   in01s01 U266598 (.o(n246649),
	.a(n246646));
   na02s01 U266599 (.o(n246648),
	.a(regtop_g_paramdata_r[21]),
	.b(n246647));
   na02s01 U266600 (.o(n212275),
	.a(n246649),
	.b(n246648));
   na02s01 U266601 (.o(n246655),
	.a(n246706),
	.b(n246650));
   in01s01 U266602 (.o(n246652),
	.a(n246651));
   na02s01 U266603 (.o(n246654),
	.a(n246653),
	.b(n246652));
   na02s01 U266604 (.o(n246669),
	.a(n246655),
	.b(n246654));
   na02s01 U266605 (.o(n246656),
	.a(vldtop_vld_syndec_ADP[1]),
	.b(vldtop_vld_syndec_UREG[29]));
   na02s01 U266606 (.o(n246667),
	.a(n246658),
	.b(n246657));
   na02s01 U266607 (.o(n246660),
	.a(n246659),
	.b(vldtop_vld_syndec_UREG[31]));
   in01s01 U266608 (.o(n246661),
	.a(n246660));
   na02f01 U266609 (.o(n246666),
	.a(n246662),
	.b(n246661));
   na02f01 U266610 (.o(n246665),
	.a(n246664),
	.b(n246663));
   no02s01 U266611 (.o(n246675),
	.a(n246671),
	.b(n246670));
   na02s01 U266612 (.o(n246678),
	.a(g_swrst_r_n),
	.b(n246889));
   in01s01 U266613 (.o(vldtop_vld_syndec_vld_outbuf_N487),
	.a(n246678));
   in01s01 U266614 (.o(n245083),
	.a(regtop_g_dsts_r));
   in01f01 U266615 (.o(n252949),
	.a(regtop_g_dmod_r));
   na02f02 U266616 (.o(n246680),
	.a(regtop_g_dack32_r_n),
	.b(regtop_g_dacksh_r_n));
   in01s01 U266617 (.o(n246682),
	.a(n246679));
   oa12s01 U266618 (.o(n246681),
	.a(n246682),
	.b(n246680),
	.c(n245083));
   oa12s01 U266619 (.o(n246683),
	.a(n246681),
	.b(regtop_g_wd_r[0]),
	.c(n246682));
   in01s01 U266620 (.o(n186714),
	.a(n246683));
   no02s01 U266621 (.o(n246686),
	.a(n246794),
	.b(n246806));
   in01s01 U266622 (.o(n246687),
	.a(n246686));
   na02s01 U266623 (.o(n246689),
	.a(n246805),
	.b(n246687));
   in01s01 U266624 (.o(n246688),
	.a(n246831));
   oa12s01 U266625 (.o(n212578),
	.a(n246691),
	.b(n246838),
	.c(n246692));
   no02s01 U266626 (.o(n246705),
	.a(n246694),
	.b(n246693));
   no02s01 U266627 (.o(n246704),
	.a(n246696),
	.b(n246695));
   no02s01 U266628 (.o(n246703),
	.a(n246698),
	.b(n246697));
   na02s01 U266629 (.o(n246701),
	.a(n246700),
	.b(n246699));
   in01s01 U266630 (.o(n246702),
	.a(n246701));
   na02s01 U266631 (.o(n246720),
	.a(n246707),
	.b(n246706));
   no02s01 U266632 (.o(n246710),
	.a(n246709),
	.b(n246708));
   in01s01 U266633 (.o(n246719),
	.a(n246710));
   no02s01 U266634 (.o(n246713),
	.a(n246712),
	.b(n246711));
   no02s01 U266635 (.o(n246716),
	.a(n246715),
	.b(n246714));
   in01s01 U266636 (.o(n246717),
	.a(n246716));
   ao12f02 U266637 (.o(n246723),
	.a(n246721),
	.b(vldtop_vld_syndec_ADP[4]),
	.c(n246722));
   in01s01 U266638 (.o(n246965),
	.a(n246723));
   na02s01 U266639 (.o(n246724),
	.a(g_swrst_r_n),
	.b(n246965));
   in01s01 U266640 (.o(vldtop_vld_syndec_vld_outbuf_N475),
	.a(n246724));
   in01s01 U266641 (.o(busiftop_N32),
	.a(busiftop_N28));
   no02s01 U266642 (.o(n246741),
	.a(n246831),
	.b(n246806));
   in01s01 U266643 (.o(n246898),
	.a(v_vldstatus_r[1]));
   na02s01 U266644 (.o(n246740),
	.a(n246830),
	.b(n246828));
   na02s01 U266645 (.o(n246739),
	.a(n246741),
	.b(n246740));
   oa12s01 U266646 (.o(n246742),
	.a(n246739),
	.b(n246741),
	.c(n246740));
   oa22s01 U266647 (.o(n212577),
	.a(n246838),
	.b(n246743),
	.c(n246742),
	.d(n246836));
   in01s01 U266648 (.o(n246745),
	.a(regtop_g_usrd_r[31]));
   na02s01 U266649 (.o(n246747),
	.a(regtop_g_usrd_r[31]),
	.b(n248978));
   in01s01 U266650 (.o(n246749),
	.a(regtop_g_usrd_r[25]));
   in01s01 U266651 (.o(n246752),
	.a(n246750));
   na02s01 U266652 (.o(n246751),
	.a(regtop_g_usrd_r[25]),
	.b(n248978));
   na02s01 U266653 (.o(n212280),
	.a(n246752),
	.b(n246751));
   in01s01 U266654 (.o(n246753),
	.a(regtop_g_usrd_r[24]));
   in01s01 U266655 (.o(n246756),
	.a(n246754));
   na02s01 U266656 (.o(n246755),
	.a(regtop_g_usrd_r[24]),
	.b(n248978));
   na02s01 U266657 (.o(n212279),
	.a(n246756),
	.b(n246755));
   in01s01 U266658 (.o(n246760),
	.a(n246758));
   na02s01 U266659 (.o(n246759),
	.a(regtop_g_usrd_r[29]),
	.b(n248978));
   na02s01 U266660 (.o(n212284),
	.a(n246760),
	.b(n246759));
   in01s01 U266661 (.o(n246761),
	.a(regtop_g_usrd_r[30]));
   in01s01 U266662 (.o(n246764),
	.a(n246762));
   na02s01 U266663 (.o(n246763),
	.a(regtop_g_usrd_r[30]),
	.b(n248978));
   na02s01 U266664 (.o(n212285),
	.a(n246764),
	.b(n246763));
   in01s01 U266665 (.o(n246765),
	.a(regtop_g_usrd_r[28]));
   in01s01 U266666 (.o(n246768),
	.a(n246766));
   na02s01 U266667 (.o(n246767),
	.a(regtop_g_usrd_r[28]),
	.b(n248978));
   na02s01 U266668 (.o(n212283),
	.a(n246768),
	.b(n246767));
   in01s01 U266669 (.o(n246769),
	.a(regtop_g_usrd_r[27]));
   in01s01 U266670 (.o(n246772),
	.a(n246770));
   na02s01 U266671 (.o(n246771),
	.a(regtop_g_usrd_r[27]),
	.b(n248978));
   na02s01 U266672 (.o(n212282),
	.a(n246772),
	.b(n246771));
   in01s01 U266673 (.o(n246774),
	.a(regtop_g_usrd_r[26]));
   in01s01 U266674 (.o(n246777),
	.a(n246775));
   na02s01 U266675 (.o(n246776),
	.a(regtop_g_usrd_r[26]),
	.b(n248978));
   na02s01 U266676 (.o(n212281),
	.a(n246777),
	.b(n246776));
   in01f02 U266677 (.o(n246788),
	.a(n246782));
   na03f01 U266678 (.o(n246784),
	.a(vldtop_vld_syndec_UREG[16]),
	.b(vldtop_vld_syndec_vld_vscdet_v_detvald_r[0]),
	.c(n246783));
   no03f02 U266679 (.o(n246790),
	.a(vldtop_vld_syndec_vld_seqhed_pre_SHIFT[4]),
	.b(n246789),
	.c(n249020));
   no02f04 U266680 (.o(n246792),
	.a(v_seqstrt_r),
	.b(n246791));
   no02f04 U266681 (.o(n246809),
	.a(vldtop_vld_syndec_ADP[4]),
	.b(n246808));
   in01s01 U266682 (.o(n246807),
	.a(n246806));
   in01s01 U266683 (.o(n249016),
	.a(g_init_vld_r_s));
   oa12s01 U266684 (.o(n246823),
	.a(v1_bs_req_n),
	.b(vldtop_vld_syndec_vld_vlfeed_feed_on),
	.c(n249016));
   no02s01 U266685 (.o(n246824),
	.a(n246838),
	.b(n246823));
   no02s01 U266686 (.o(n246825),
	.a(n246824),
	.b(FE_OFN68_n247591));
   in01s01 U266687 (.o(n247145),
	.a(vldtop_vld_syndec_vld_vlfeed_dselect_r));
   na02s01 U266688 (.o(n246832),
	.a(n246827),
	.b(n246826));
   in01s01 U266689 (.o(n246835),
	.a(n246832));
   na02s01 U266690 (.o(n246829),
	.a(n246828),
	.b(n246807));
   in01s01 U266691 (.o(n246833),
	.a(n246834));
   na02s01 U266692 (.o(n246839),
	.a(n252485),
	.b(regtop_g_nfst_r[11]));
   ao12s01 U266693 (.o(n246841),
	.a(n252269),
	.b(n252270),
	.c(regtop_g_wd_r[0]));
   in01s01 U266694 (.o(n184629),
	.a(n246842));
   in01s01 U266695 (.o(n246844),
	.a(vldtop_vld_syndec_vld_vscdet_v_prezerotmp_r[0]));
   in01s01 U266696 (.o(n246913),
	.a(n249003));
   no04f03 U266697 (.o(n246843),
	.a(vldtop_vld_syndec_UREG[0]),
	.b(vldtop_vld_syndec_UREG[3]),
	.c(vldtop_vld_syndec_UREG[6]),
	.d(vldtop_vld_syndec_UREG[7]));
   na02s01 U266698 (.o(n246917),
	.a(n246964),
	.b(n246843));
   oa22s01 U266699 (.o(n212572),
	.a(n246844),
	.b(n249028),
	.c(n246913),
	.d(n246917));
   in01s01 U266700 (.o(n246851),
	.a(regtop_g_udb2_r[1]));
   ao22s01 U266701 (.o(n246852),
	.a(regtop_g_udb2_r[0]),
	.b(n246851),
	.c(regtop_g_udb2_r[1]),
	.d(n246062));
   in01s01 U266702 (.o(n246854),
	.a(y1_bs_data[9]));
   no03m01 U266703 (.o(n246856),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[9]),
	.b(n247494),
	.c(FE_OFN68_n247591));
   na02s01 U266704 (.o(n246858),
	.a(regtop_g_udb2_r[0]),
	.b(regtop_g_udb2_r[1]));
   in01s01 U266705 (.o(n246876),
	.a(n246858));
   na02s01 U266706 (.o(n246859),
	.a(regtop_g_udb2_r[2]),
	.b(n246876));
   in01s01 U266707 (.o(n246871),
	.a(n246859));
   in01s01 U266708 (.o(n246860),
	.a(regtop_g_udb2_r[3]));
   in01s01 U266709 (.o(n252299),
	.a(regtop_g_ferror_r));
   no02s01 U266710 (.o(n252240),
	.a(n252757),
	.b(n252299));
   na02s01 U266711 (.o(n246864),
	.a(n246863),
	.b(n252240));
   ao22s01 U266712 (.o(n246866),
	.a(n252377),
	.b(n252245),
	.c(regtop_g_fbst_r[0]),
	.d(n252300));
   na02s01 U266713 (.o(n246867),
	.a(regtop_g_udb2_r[3]),
	.b(regtop_g_udb2_r[4]));
   in01s01 U266714 (.o(n246868),
	.a(n246867));
   in01s01 U266715 (.o(n246875),
	.a(n246874));
   in01s01 U266716 (.o(n211959),
	.a(n246878));
   no02s01 U266717 (.o(n246879),
	.a(regtop_g_udb2_r[5]),
	.b(n246935));
   in01s01 U266718 (.o(n211956),
	.a(n246881));
   in01s01 U266719 (.o(n246897),
	.a(n246882));
   in01s01 U266720 (.o(n246888),
	.a(n246883));
   in01s01 U266721 (.o(n246887),
	.a(n246884));
   in01s01 U266722 (.o(n246886),
	.a(n246885));
   in01s01 U266723 (.o(n247028),
	.a(n246889));
   na02s01 U266724 (.o(n246895),
	.a(v_vldstatus_r[4]),
	.b(v_vldstatus_r[1]));
   in01s01 U266725 (.o(n246907),
	.a(regtop_g_udb0_r[2]));
   no02f01 U266726 (.o(n246949),
	.a(n246952),
	.b(n246907));
   ao12s01 U266727 (.o(n246905),
	.a(n246949),
	.b(n246952),
	.c(n246907));
   in01s01 U266728 (.o(n246912),
	.a(regtop_g_udb1_r[2]));
   na02f01 U266729 (.o(n246959),
	.a(regtop_g_udb1_r[0]),
	.b(regtop_g_udb1_r[1]));
   ao12s01 U266730 (.o(n246910),
	.a(n246956),
	.b(n246959),
	.c(n246912));
   in01s01 U266731 (.o(n246918),
	.a(vldtop_vld_syndec_vld_vscdet_v_prezerotmp_r[1]));
   no03s01 U266732 (.o(n246915),
	.a(vldtop_vld_syndec_UREG[8]),
	.b(n246914),
	.c(n246913));
   in01s01 U266733 (.o(n246916),
	.a(n246915));
   oa22s01 U266734 (.o(n212574),
	.a(n246918),
	.b(n249028),
	.c(n246917),
	.d(n246916));
   na02s01 U266735 (.o(n246919),
	.a(regtop_g_udb0_r[4]),
	.b(regtop_g_udb0_r[3]));
   in01s01 U266736 (.o(n246920),
	.a(n246919));
   in01s01 U266737 (.o(n246921),
	.a(regtop_g_udb0_r[5]));
   na02s01 U266738 (.o(n246927),
	.a(regtop_g_udb1_r[4]),
	.b(regtop_g_udb1_r[3]));
   in01s01 U266739 (.o(n246928),
	.a(n246927));
   in01s01 U266740 (.o(n246929),
	.a(regtop_g_udb1_r[5]));
   in01s01 U266741 (.o(n246932),
	.a(regtop_g_udb1_r[6]));
   in01s01 U266742 (.o(n246938),
	.a(n246935));
   in01s01 U266743 (.o(n246936),
	.a(regtop_g_udb2_r[5]));
   no02s01 U266744 (.o(n246937),
	.a(regtop_g_udb2_r[6]),
	.b(n246936));
   ao22s01 U266745 (.o(n246942),
	.a(n246938),
	.b(n246937),
	.c(regtop_g_udb2_r[6]),
	.d(n246936));
   na02s01 U266746 (.o(n246944),
	.a(regtop_g_paramadr_r[4]),
	.b(n252642));
   no02f01 U266747 (.o(n246947),
	.a(n252517),
	.b(n246944));
   in01s01 U266748 (.o(n246946),
	.a(regtop_g_ld_r));
   na02s01 U266749 (.o(n246945),
	.a(regtop_g_paramdata_r[24]),
	.b(n246947));
   oa12s01 U266750 (.o(n212175),
	.a(n246945),
	.b(n246947),
	.c(n246946));
   in01s01 U266751 (.o(n246951),
	.a(regtop_g_udb0_r[3]));
   na02s01 U266752 (.o(n247035),
	.a(n246949),
	.b(regtop_g_udb0_r[3]));
   oa12s01 U266753 (.o(n246950),
	.a(n247035),
	.b(n246949),
	.c(regtop_g_udb0_r[3]));
   in01s01 U266754 (.o(n246955),
	.a(regtop_g_udb0_r[1]));
   oa12s01 U266755 (.o(n246953),
	.a(n246952),
	.b(regtop_g_udb0_r[0]),
	.c(regtop_g_udb0_r[1]));
   in01s01 U266756 (.o(n246958),
	.a(regtop_g_udb1_r[3]));
   na02s01 U266757 (.o(n247046),
	.a(n246956),
	.b(regtop_g_udb1_r[3]));
   oa12s01 U266758 (.o(n246957),
	.a(n247046),
	.b(n246956),
	.c(regtop_g_udb1_r[3]));
   in01s01 U266759 (.o(n246961),
	.a(regtop_g_udb1_r[1]));
   oa12s01 U266760 (.o(n246960),
	.a(n246959),
	.b(regtop_g_udb1_r[0]),
	.c(regtop_g_udb1_r[1]));
   in01s01 U266761 (.o(n246962),
	.a(regtop_g_udb1_r[0]));
   na02s01 U266762 (.o(n246966),
	.a(n246994),
	.b(n246723));
   in01s01 U266763 (.o(n246975),
	.a(n246991));
   in01s01 U266764 (.o(n246986),
	.a(n246980));
   in01s01 U266765 (.o(n246993),
	.a(n246987));
   no02s02 U266766 (.o(n247005),
	.a(n247001),
	.b(n247000));
   in01s01 U266767 (.o(n247025),
	.a(n247009));
   in01f01 U266768 (.o(n247016),
	.a(n247014));
   na02f02 U266769 (.o(n247022),
	.a(n247016),
	.b(n247015));
   in01s01 U266770 (.o(n247032),
	.a(vldtop_vld_syndec_vld_vscdet_v_seqerr_r));
   oa22m01 U266771 (.o(n212463),
	.a(n246370),
	.b(n249255),
	.c(n249028),
	.d(n247032));
   no02s01 U266772 (.o(n247037),
	.a(n247036),
	.b(n247035));
   no02s01 U266773 (.o(n247041),
	.a(regtop_g_udb0_r[5]),
	.b(n247039));
   in01s01 U266774 (.o(n247047),
	.a(n247050));
   no02s01 U266775 (.o(n247048),
	.a(n247047),
	.b(n247046));
   no02s01 U266776 (.o(n247052),
	.a(regtop_g_udb1_r[5]),
	.b(n247050));
   no02f01 U266777 (.o(n248118),
	.a(n247062),
	.b(n251621));
   no02f01 U266778 (.o(n248355),
	.a(n247062),
	.b(FE_OFN24_n250486));
   ao22s01 U266779 (.o(n247066),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1146]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[122]));
   no02f01 U266780 (.o(n248357),
	.a(n247062),
	.b(n252195));
   ao22s01 U266781 (.o(n247065),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1658]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[634]));
   no02f01 U266782 (.o(n248119),
	.a(n247062),
	.b(FE_OFN28_n251337));
   no02f01 U266783 (.o(n247057),
	.a(n247062),
	.b(FE_OFN22_n250202));
   ao22s01 U266786 (.o(n247064),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1402]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[378]));
   no02f01 U266787 (.o(n248121),
	.a(n247062),
	.b(FE_OFN32_n251904));
   no02f01 U266788 (.o(n248120),
	.a(n247062),
	.b(FE_OFN556_n250770));
   ao22s01 U266789 (.o(n247063),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1914]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[890]));
   ao22s01 U266790 (.o(n247073),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1210]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[186]));
   ao22s01 U266791 (.o(n247072),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1722]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[698]));
   no02f01 U266792 (.o(n247067),
	.a(n247069),
	.b(FE_OFN22_n250202));
   ao22s01 U266794 (.o(n247071),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1466]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[442]));
   ao22s01 U266795 (.o(n247070),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1978]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[954]));
   no02f01 U266796 (.o(n248370),
	.a(FE_OFN8_n247076),
	.b(n251621));
   no02f01 U266797 (.o(n248369),
	.a(FE_OFN8_n247076),
	.b(FE_OFN24_n250486));
   ao22s01 U266798 (.o(n247080),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1274]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[250]));
   no02f01 U266799 (.o(n248372),
	.a(FE_OFN8_n247076),
	.b(n252195));
   no02f01 U266800 (.o(n248371),
	.a(FE_OFN8_n247076),
	.b(n251053));
   ao22s01 U266801 (.o(n247079),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1786]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[762]));
   no02f01 U266802 (.o(n248373),
	.a(FE_OFN8_n247076),
	.b(FE_OFN28_n251337));
   no02f01 U266803 (.o(n247074),
	.a(FE_OFN8_n247076),
	.b(FE_OFN22_n250202));
   ao22s01 U266806 (.o(n247078),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1530]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[506]));
   no02f01 U266807 (.o(n248375),
	.a(FE_OFN8_n247076),
	.b(FE_OFN32_n251904));
   no02f01 U266808 (.o(n248374),
	.a(FE_OFN8_n247076),
	.b(FE_OFN556_n250770));
   ao22f01 U266809 (.o(n247077),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2042]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1018]));
   no02f01 U266810 (.o(n248138),
	.a(n247082),
	.b(n251621));
   no02f01 U266811 (.o(n248380),
	.a(n247082),
	.b(FE_OFN24_n250486));
   ao22s01 U266812 (.o(n247086),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1082]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[58]));
   no02f01 U266813 (.o(n248382),
	.a(n247082),
	.b(n252195));
   no02f01 U266814 (.o(n248381),
	.a(n247082),
	.b(n251053));
   ao22s01 U266815 (.o(n247085),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1594]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[570]));
   no02f02 U266816 (.o(n248139),
	.a(n247082),
	.b(FE_OFN28_n251337));
   no02f01 U266817 (.o(n247509),
	.a(n247082),
	.b(FE_OFN22_n250202));
   ao22s01 U266818 (.o(n247084),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1338]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[314]));
   no02f01 U266819 (.o(n248141),
	.a(n247082),
	.b(FE_OFN32_n251904));
   ao22s01 U266820 (.o(n247083),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1850]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[826]));
   na04f03 U266821 (.o(n247087),
	.a(n247086),
	.b(n247085),
	.c(n247084),
	.d(n247083));
   no02f01 U266822 (.o(n248150),
	.a(n247094),
	.b(n251621));
   no02f01 U266823 (.o(n248391),
	.a(n247094),
	.b(FE_OFN24_n250486));
   ao22s01 U266824 (.o(n247098),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1114]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[90]));
   no02f01 U266825 (.o(n248393),
	.a(n247094),
	.b(n252195));
   no02f01 U266826 (.o(n248392),
	.a(n247094),
	.b(n251053));
   no02f01 U266827 (.o(n248151),
	.a(n247094),
	.b(FE_OFN28_n251337));
   no02f01 U266828 (.o(n247092),
	.a(n247094),
	.b(FE_OFN22_n250202));
   ao22s01 U266831 (.o(n247096),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1370]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[346]));
   no02f01 U266832 (.o(n248153),
	.a(n247094),
	.b(FE_OFN33_n251904));
   no02f01 U266833 (.o(n248152),
	.a(n247094),
	.b(n250770));
   ao22s01 U266834 (.o(n247095),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1882]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[858]));
   no02f01 U266835 (.o(n248159),
	.a(n247101),
	.b(n251621));
   no02f01 U266836 (.o(n248158),
	.a(n247101),
	.b(FE_OFN24_n250486));
   ao22s01 U266837 (.o(n247105),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1178]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[154]));
   no02f01 U266838 (.o(n248399),
	.a(n247101),
	.b(n252195));
   no02f01 U266839 (.o(n248398),
	.a(n247101),
	.b(n251053));
   ao22s01 U266840 (.o(n247104),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1690]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[666]));
   no02f01 U266841 (.o(n248160),
	.a(n247101),
	.b(FE_OFN28_n251337));
   no02f01 U266842 (.o(n247099),
	.a(n247101),
	.b(FE_OFN22_n250202));
   ao22f01 U266844 (.o(n247103),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1434]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[410]));
   no02f01 U266845 (.o(n248162),
	.a(n247101),
	.b(FE_OFN32_n251904));
   no02f10 U266846 (.o(n248161),
	.a(n247101),
	.b(n250770));
   ao22s01 U266847 (.o(n247102),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1946]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[922]));
   no02f01 U266848 (.o(n248405),
	.a(n247109),
	.b(n251621));
   no02f01 U266849 (.o(n248404),
	.a(n247109),
	.b(FE_OFN24_n250486));
   ao22s01 U266850 (.o(n247113),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1242]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[218]));
   no02f01 U266851 (.o(n248407),
	.a(n247109),
	.b(n252195));
   no02f01 U266852 (.o(n248406),
	.a(n247109),
	.b(n251053));
   ao22s01 U266853 (.o(n247112),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1754]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[730]));
   no02f01 U266854 (.o(n247107),
	.a(n247109),
	.b(FE_OFN22_n250202));
   ao22s01 U266857 (.o(n247111),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1498]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[474]));
   no02f10 U266858 (.o(n248168),
	.a(n247109),
	.b(FE_OFN33_n251904));
   ao22s01 U266859 (.o(n247110),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2010]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[986]));
   no02f01 U266860 (.o(n248173),
	.a(n251621),
	.b(n247114));
   no02f01 U266861 (.o(n248413),
	.a(FE_OFN24_n250486),
	.b(n247114));
   ao22s01 U266862 (.o(n247118),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1050]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[26]));
   no02f01 U266863 (.o(n248415),
	.a(n252195),
	.b(n247114));
   no02f01 U266864 (.o(n248414),
	.a(n251053),
	.b(n247114));
   ao22s01 U266865 (.o(n247117),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1562]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[538]));
   no02f01 U266866 (.o(n248174),
	.a(FE_OFN28_n251337),
	.b(n247114));
   no02f01 U266867 (.o(n247531),
	.a(FE_OFN22_n250202),
	.b(n247114));
   ao22s01 U266868 (.o(n247116),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1306]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[282]));
   no02f01 U266869 (.o(n248176),
	.a(FE_OFN32_n251904),
	.b(n247114));
   no02f01 U266870 (.o(n248175),
	.a(n250770),
	.b(n247114));
   ao22s01 U266871 (.o(n247115),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1818]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[794]));
   na04f01 U266872 (.o(n247119),
	.a(n247118),
	.b(n247117),
	.c(n247116),
	.d(n247115));
   na02f01 U266873 (.o(regtop_w1_hdi00_q[26]),
	.a(n247124),
	.b(FE_OFN368_n247123));
   no02s01 U266874 (.o(n247130),
	.a(vldtop_vld_syndec_UREG[21]),
	.b(n247591));
   na02s01 U266875 (.o(n247128),
	.a(g_swrst_r_n),
	.b(n247127));
   no02s01 U266876 (.o(n247134),
	.a(vldtop_vld_syndec_UREG[25]),
	.b(n247591));
   na02s01 U266877 (.o(n247132),
	.a(g_swrst_r_n),
	.b(n247131));
   in01s01 U266878 (.o(n247135),
	.a(vldtop_vld_syndec_vld_seqhed_state_0_));
   na02s01 U266879 (.o(n247136),
	.a(v_seqstrt_r),
	.b(n247135));
   no02s01 U266880 (.o(n247137),
	.a(n246370),
	.b(n247136));
   na02s01 U266881 (.o(n247138),
	.a(n249064),
	.b(vldtop_vld_syndec_vld_seqhed_state_0_));
   no02s01 U266882 (.o(n247142),
	.a(vldtop_vld_syndec_UREG[6]),
	.b(FE_OFN68_n247591));
   na02s01 U266883 (.o(n247140),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247139));
   ao12f01 U266884 (.o(n247152),
	.a(FE_OFN68_n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[7]));
   ao22f01 U266885 (.o(n247153),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[25]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[25]));
   no02s01 U266886 (.o(n247158),
	.a(vldtop_vld_syndec_UREG[12]),
	.b(FE_OFN68_n247591));
   na02s01 U266887 (.o(n247156),
	.a(FE_OFN2_g_swrst_r_n),
	.b(FE_OFN540_vldtop_vld_syndec_vld_vlfeed_lower_12_));
   no02s01 U266888 (.o(n247162),
	.a(vldtop_vld_syndec_UREG[31]),
	.b(FE_OFN68_n247591));
   na02s01 U266889 (.o(n247160),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247159));
   no02s01 U266890 (.o(n247166),
	.a(vldtop_vld_syndec_UREG[30]),
	.b(FE_OFN68_n247591));
   na02s01 U266891 (.o(n247164),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247163));
   ao12f01 U266892 (.o(n247168),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[29]));
   no02s01 U266893 (.o(n247172),
	.a(vldtop_vld_syndec_UREG[13]),
	.b(FE_OFN68_n247591));
   in01s01 U266894 (.o(n247169),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[13]));
   no02s01 U266895 (.o(n247176),
	.a(vldtop_vld_syndec_UREG[20]),
	.b(FE_OFN68_n247591));
   na02s01 U266896 (.o(n247174),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247173));
   ao22f01 U266897 (.o(n247177),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[20]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[20]));
   no02s01 U266898 (.o(n247182),
	.a(vldtop_vld_syndec_UREG[4]),
	.b(FE_OFN68_n247591));
   in01s01 U266899 (.o(n247179),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[4]));
   na02s01 U266900 (.o(n247180),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247179));
   no02s01 U266901 (.o(n247186),
	.a(vldtop_vld_syndec_UREG[16]),
	.b(FE_OFN68_n247591));
   na02s01 U266902 (.o(n247184),
	.a(FE_OFN2_g_swrst_r_n),
	.b(FE_OFN525_vldtop_vld_syndec_vld_vlfeed_lower_16_));
   ao22f01 U266903 (.o(n247187),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[21]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[21]));
   ao12f01 U266904 (.o(n247190),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[0]));
   ao22f01 U266905 (.o(n247189),
	.a(FE_OFN14_n247150),
	.b(vldtop_vld_syndec_vld_vlfeed_temporal[0]),
	.c(vldtop_vld_syndec_vld_vlfeed_lower[0]),
	.d(FE_OFN577_n247126));
   in01s01 U266906 (.o(n247191),
	.a(y1_bs_data[19]));
   no03f01 U266907 (.o(n247193),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[19]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no02m01 U266908 (.o(n253051),
	.a(n247194),
	.b(n247193));
   no02s01 U266909 (.o(n247198),
	.a(vldtop_vld_syndec_UREG[17]),
	.b(FE_OFN68_n247591));
   in01s01 U266910 (.o(n247195),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[17]));
   na02f01 U266911 (.o(n247196),
	.a(g_swrst_r_n),
	.b(n247195));
   no02s01 U266912 (.o(n247202),
	.a(vldtop_vld_syndec_UREG[15]),
	.b(n247591));
   in01s01 U266913 (.o(n247199),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[15]));
   na02s01 U266914 (.o(n247200),
	.a(g_swrst_r_n),
	.b(n247199));
   ao22f01 U266915 (.o(n247204),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[24]),
	.b(n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[24]));
   ao22f01 U266916 (.o(n247206),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[12]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[12]));
   ao22f01 U266917 (.o(n247208),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[18]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[18]));
   no02s01 U266918 (.o(n247213),
	.a(vldtop_vld_syndec_UREG[27]),
	.b(FE_OFN68_n247591));
   na02s01 U266919 (.o(n247211),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247210));
   no02s01 U266920 (.o(n247217),
	.a(vldtop_vld_syndec_UREG[7]),
	.b(FE_OFN68_n247591));
   in01s01 U266921 (.o(n247214),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[7]));
   na02s01 U266922 (.o(n247215),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247214));
   ao12f01 U266923 (.o(n247219),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[30]));
   ao22f01 U266924 (.o(n247220),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[14]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[14]));
   no02s01 U266925 (.o(n247225),
	.a(vldtop_vld_syndec_UREG[10]),
	.b(FE_OFN68_n247591));
   na02s01 U266926 (.o(n247223),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247222));
   ao12f01 U266927 (.o(n247227),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[8]));
   no02s01 U266928 (.o(n247231),
	.a(vldtop_vld_syndec_UREG[5]),
	.b(n247591));
   in01s01 U266929 (.o(n247228),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[5]));
   na02s01 U266930 (.o(n247229),
	.a(g_swrst_r_n),
	.b(n247228));
   in01s01 U266931 (.o(n247232),
	.a(y1_bs_data[3]));
   in01s01 U266932 (.o(n247236),
	.a(y1_bs_data[10]));
   no03m01 U266933 (.o(n247238),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[10]),
	.b(n247494),
	.c(FE_OFN68_n247591));
   no02s01 U266934 (.o(n247243),
	.a(vldtop_vld_syndec_UREG[26]),
	.b(FE_OFN68_n247591));
   na02s01 U266935 (.o(n247241),
	.a(FE_OFN2_g_swrst_r_n),
	.b(FE_OFN543_vldtop_vld_syndec_vld_vlfeed_lower_26_));
   ao12f01 U266936 (.o(n247245),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[1]));
   ao22f01 U266937 (.o(n247244),
	.a(FE_OFN14_n247150),
	.b(vldtop_vld_syndec_vld_vlfeed_temporal[1]),
	.c(vldtop_vld_syndec_vld_vlfeed_lower[1]),
	.d(FE_OFN577_n247126));
   ao12f01 U266938 (.o(n247247),
	.a(FE_OFN68_n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[16]));
   ao22f01 U266939 (.o(n247246),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[16]),
	.b(n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[16]));
   ao12f01 U266940 (.o(n247249),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[13]));
   ao22f01 U266941 (.o(n247248),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[13]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[13]));
   ao12f01 U266942 (.o(n247251),
	.a(FE_OFN68_n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[22]));
   ao22f01 U266943 (.o(n247250),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[22]),
	.b(n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[22]));
   in01s01 U266944 (.o(n247255),
	.a(vldtop_vld_syndec_vld_seqhed_pre_SHIFT[3]));
   ao22f01 U266945 (.o(n247256),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[27]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[27]));
   no02s01 U266946 (.o(n247261),
	.a(vldtop_vld_syndec_UREG[8]),
	.b(FE_OFN68_n247591));
   in01s01 U266947 (.o(n247258),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[8]));
   na02s01 U266948 (.o(n247259),
	.a(g_swrst_r_n),
	.b(n247258));
   no02s01 U266949 (.o(n247267),
	.a(vldtop_vld_syndec_UREG[9]),
	.b(FE_OFN68_n247591));
   in01s01 U266950 (.o(n247264),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[9]));
   na02s01 U266951 (.o(n247265),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247264));
   ao22f01 U266952 (.o(n247268),
	.a(FE_OFN14_n247150),
	.b(vldtop_vld_syndec_vld_vlfeed_temporal[2]),
	.c(vldtop_vld_syndec_vld_vlfeed_lower[2]),
	.d(FE_OFN577_n247126));
   no02s01 U266953 (.o(n247275),
	.a(vldtop_vld_syndec_UREG[18]),
	.b(FE_OFN68_n247591));
   na02s01 U266954 (.o(n247273),
	.a(FE_OFN2_g_swrst_r_n),
	.b(FE_OFN537_vldtop_vld_syndec_vld_vlfeed_lower_18_));
   no02s01 U266955 (.o(n247279),
	.a(vldtop_vld_syndec_UREG[22]),
	.b(FE_OFN68_n247591));
   na02s01 U266956 (.o(n247277),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247276));
   no03f01 U266957 (.o(n247281),
	.a(n247591),
	.b(n247441),
	.c(y1_bs_data[27]));
   no03f01 U266958 (.o(n247280),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[27]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   in01s01 U266959 (.o(n247282),
	.a(y1_bs_data[31]));
   no03f01 U266960 (.o(n247284),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[31]),
	.b(n247494),
	.c(FE_OFN68_n247591));
   no02s01 U266961 (.o(n247288),
	.a(vldtop_vld_syndec_UREG[1]),
	.b(FE_OFN68_n247591));
   no03f01 U266962 (.o(n247286),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[1]),
	.b(n247126),
	.c(FE_OFN68_n247591));
   no02s01 U266963 (.o(n247292),
	.a(vldtop_vld_syndec_UREG[29]),
	.b(FE_OFN68_n247591));
   na02s01 U266964 (.o(n247290),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247289));
   no02s01 U266965 (.o(n247296),
	.a(vldtop_vld_syndec_UREG[23]),
	.b(n247591));
   na02s01 U266966 (.o(n247294),
	.a(g_swrst_r_n),
	.b(n247293));
   no02s01 U266967 (.o(n247298),
	.a(vldtop_vld_syndec_UREG[0]),
	.b(FE_OFN68_n247591));
   no03f01 U266968 (.o(n247297),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[0]),
	.b(n247126),
	.c(FE_OFN68_n247591));
   ao22f01 U266969 (.o(n247299),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[9]),
	.b(n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[9]));
   ao22f01 U266970 (.o(n247301),
	.a(FE_OFN14_n247150),
	.b(vldtop_vld_syndec_vld_vlfeed_temporal[3]),
	.c(vldtop_vld_syndec_vld_vlfeed_lower[3]),
	.d(FE_OFN577_n247126));
   ao22f01 U266971 (.o(n247304),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[23]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[23]));
   ao12f01 U266972 (.o(n247307),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[10]));
   no02s01 U266973 (.o(n247311),
	.a(vldtop_vld_syndec_UREG[2]),
	.b(FE_OFN68_n247591));
   in01s01 U266974 (.o(n247308),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[2]));
   na02s01 U266975 (.o(n247309),
	.a(g_swrst_r_n),
	.b(n247308));
   no02s01 U266976 (.o(n247315),
	.a(vldtop_vld_syndec_UREG[11]),
	.b(n247591));
   in01s01 U266977 (.o(n247312),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[11]));
   na02s01 U266978 (.o(n247313),
	.a(g_swrst_r_n),
	.b(n247312));
   no02s01 U266979 (.o(n247319),
	.a(vldtop_vld_syndec_UREG[14]),
	.b(FE_OFN68_n247591));
   na02s01 U266980 (.o(n247317),
	.a(FE_OFN2_g_swrst_r_n),
	.b(FE_OFN530_vldtop_vld_syndec_vld_vlfeed_lower_14_));
   in01s01 U266981 (.o(n247320),
	.a(y1_bs_data[5]));
   in01s01 U266982 (.o(n247323),
	.a(n247321));
   no03f01 U266983 (.o(n247322),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[5]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no02m01 U266984 (.o(n253065),
	.a(n247323),
	.b(n247322));
   in01s01 U266985 (.o(n247324),
	.a(y1_bs_data[15]));
   no03m01 U266986 (.o(n247326),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[15]),
	.b(n247494),
	.c(FE_OFN68_n247591));
   no02m01 U266987 (.o(n253055),
	.a(n247327),
	.b(n247326));
   ao12f01 U266988 (.o(n247329),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[5]));
   ao22f01 U266989 (.o(n247330),
	.a(FE_OFN14_n247150),
	.b(vldtop_vld_syndec_vld_vlfeed_temporal[4]),
	.c(vldtop_vld_syndec_vld_vlfeed_lower[4]),
	.d(n247126));
   no02s01 U266990 (.o(n247335),
	.a(vldtop_vld_syndec_UREG[28]),
	.b(FE_OFN68_n247591));
   na02s01 U266991 (.o(n247333),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247332));
   ao22f01 U266992 (.o(n247336),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[6]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[6]));
   in01s01 U266993 (.o(n247338),
	.a(y1_bs_data[13]));
   in01s01 U266994 (.o(n247341),
	.a(n247339));
   no03f01 U266995 (.o(n247340),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[13]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   in01s01 U266996 (.o(n247342),
	.a(y1_bs_data[7]));
   in01s01 U266997 (.o(n247345),
	.a(n247343));
   no03f01 U266998 (.o(n247344),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[7]),
	.b(FE_OFN18_n247494),
	.c(FE_OFN68_n247591));
   no02m01 U266999 (.o(n253063),
	.a(n247345),
	.b(n247344));
   in01s01 U267000 (.o(n247346),
	.a(y1_bs_data[30]));
   na03m02 U267001 (.o(n247347),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247346));
   in01s01 U267002 (.o(n247349),
	.a(n247347));
   no03f01 U267003 (.o(n247348),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[30]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no02m01 U267004 (.o(n253040),
	.a(n247349),
	.b(n247348));
   ao12f01 U267005 (.o(n247355),
	.a(n247591),
	.b(FE_OFN16_n247350),
	.c(y1_bs_data[17]));
   ao22f01 U267006 (.o(n247354),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[17]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[17]));
   in01s01 U267007 (.o(n247356),
	.a(y1_bs_data[23]));
   na03f01 U267008 (.o(n247357),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247356));
   no03f01 U267009 (.o(n247358),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[23]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   in01s01 U267010 (.o(n247360),
	.a(y1_bs_data[14]));
   in01s01 U267011 (.o(n247363),
	.a(n247361));
   no03f01 U267012 (.o(n247362),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[14]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no02m01 U267013 (.o(n253056),
	.a(n247363),
	.b(n247362));
   no02s01 U267014 (.o(n247367),
	.a(vldtop_vld_syndec_UREG[19]),
	.b(FE_OFN68_n247591));
   na02s01 U267015 (.o(n247365),
	.a(g_swrst_r_n),
	.b(n247364));
   no02s01 U267016 (.o(n247371),
	.a(vldtop_vld_syndec_UREG[24]),
	.b(FE_OFN68_n247591));
   na02s01 U267017 (.o(n247369),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247368));
   in01s01 U267018 (.o(n247374),
	.a(y1_bs_data[0]));
   ao22f01 U267019 (.o(n247382),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[15]),
	.b(FE_OFN577_n247126),
	.c(FE_OFN14_n247150),
	.d(vldtop_vld_syndec_vld_vlfeed_temporal[15]));
   no02s01 U267020 (.o(n247385),
	.a(vldtop_vld_syndec_UREG[3]),
	.b(FE_OFN68_n247591));
   no03f01 U267021 (.o(n247384),
	.a(vldtop_vld_syndec_vld_vlfeed_lower[3]),
	.b(n247126),
	.c(FE_OFN68_n247591));
   in01s01 U267022 (.o(n247386),
	.a(y1_bs_data[28]));
   na03m02 U267023 (.o(n247387),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247386));
   in01s01 U267024 (.o(n247389),
	.a(n247387));
   no03f01 U267025 (.o(n247388),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[28]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no02m01 U267026 (.o(n253042),
	.a(n247389),
	.b(n247388));
   in01s01 U267027 (.o(n247390),
	.a(y1_bs_data[22]));
   in01s01 U267028 (.o(n247393),
	.a(n247391));
   no03f01 U267029 (.o(n247392),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[22]),
	.b(n247494),
	.c(FE_OFN68_n247591));
   no02m01 U267030 (.o(n253048),
	.a(n247393),
	.b(n247392));
   ao22s01 U267032 (.o(n247398),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1145]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[121]));
   ao22s01 U267033 (.o(n247397),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1657]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[633]));
   ao22s01 U267034 (.o(n247396),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1401]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[377]));
   ao22s01 U267035 (.o(n247395),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1913]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[889]));
   ao22s01 U267037 (.o(n247403),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1209]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[185]));
   ao22s01 U267038 (.o(n247402),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1721]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[697]));
   ao22s01 U267039 (.o(n247401),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1465]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[441]));
   ao22s01 U267040 (.o(n247400),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1977]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[953]));
   ao22s01 U267041 (.o(n247407),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1273]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[249]));
   ao22s01 U267042 (.o(n247406),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1785]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[761]));
   ao22s01 U267043 (.o(n247405),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1529]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[505]));
   ao22s01 U267044 (.o(n247404),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2041]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1017]));
   ao22s01 U267046 (.o(n247412),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1081]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[57]));
   ao22s01 U267047 (.o(n247411),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1593]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[569]));
   ao22s01 U267048 (.o(n247410),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1337]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[313]));
   ao22s01 U267049 (.o(n247409),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1849]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[825]));
   ao22s01 U267051 (.o(n247421),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1113]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[89]));
   ao22s01 U267052 (.o(n247420),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1625]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[601]));
   ao22s01 U267053 (.o(n247419),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1369]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[345]));
   ao22s01 U267054 (.o(n247425),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1177]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[153]));
   ao22s01 U267055 (.o(n247424),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1689]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[665]));
   ao22s01 U267056 (.o(n247423),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1433]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[409]));
   ao22s01 U267057 (.o(n247422),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1945]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[921]));
   ao22s01 U267058 (.o(n247429),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1241]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[217]));
   ao22s01 U267059 (.o(n247428),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1753]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[729]));
   ao22s01 U267060 (.o(n247427),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1497]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[473]));
   ao22s01 U267061 (.o(n247426),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2009]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[985]));
   ao22s01 U267063 (.o(n247434),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1049]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[25]));
   ao22s01 U267064 (.o(n247433),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1561]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[537]));
   ao22s01 U267065 (.o(n247432),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1305]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[281]));
   ao22s01 U267066 (.o(n247431),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1817]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[793]));
   na02f04 U267067 (.o(regtop_w1_hdi00_q[25]),
	.a(n247440),
	.b(n247439));
   no03f01 U267068 (.o(n247444),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[11]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no03f01 U267069 (.o(n247448),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[25]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   in01s01 U267070 (.o(n247450),
	.a(y1_bs_data[26]));
   in01s01 U267071 (.o(n247454),
	.a(n247451));
   no03f01 U267072 (.o(n247453),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[26]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no02m01 U267073 (.o(n253044),
	.a(n247454),
	.b(n247453));
   in01s01 U267074 (.o(n247455),
	.a(y1_bs_data[8]));
   no03f01 U267075 (.o(n247457),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[8]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   in01s01 U267076 (.o(n247459),
	.a(y1_bs_data[16]));
   in01s01 U267077 (.o(n247462),
	.a(n247460));
   no03f01 U267078 (.o(n247461),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[16]),
	.b(n247494),
	.c(FE_OFN68_n247591));
   no02f01 U267079 (.o(n253054),
	.a(n247462),
	.b(n247461));
   in01s01 U267080 (.o(n247463),
	.a(y1_bs_data[24]));
   no03m01 U267081 (.o(n247465),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[24]),
	.b(n247494),
	.c(FE_OFN68_n247591));
   in01s01 U267082 (.o(n247467),
	.a(y1_bs_data[29]));
   na03m02 U267083 (.o(n247468),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247467));
   in01s01 U267084 (.o(n247470),
	.a(n247468));
   no03f01 U267085 (.o(n247469),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[29]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no02m01 U267086 (.o(n253041),
	.a(n247470),
	.b(n247469));
   in01s01 U267087 (.o(n247471),
	.a(y1_bs_data[17]));
   na03f01 U267088 (.o(n247472),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247471));
   no03f01 U267089 (.o(n247473),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[17]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no02m01 U267090 (.o(n253053),
	.a(n247474),
	.b(n247473));
   in01s01 U267091 (.o(n247475),
	.a(y1_bs_data[20]));
   na03f01 U267092 (.o(n247476),
	.a(FE_OFN2_g_swrst_r_n),
	.b(n247494),
	.c(n247475));
   no03f01 U267093 (.o(n247477),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[20]),
	.b(n247494),
	.c(FE_OFN68_n247591));
   no02m01 U267094 (.o(n253050),
	.a(n247478),
	.b(n247477));
   in01s01 U267095 (.o(n247479),
	.a(y1_bs_data[4]));
   no03f01 U267096 (.o(n247481),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[4]),
	.b(n247494),
	.c(FE_OFN68_n247591));
   in01s01 U267097 (.o(n247483),
	.a(y1_bs_data[12]));
   in01s01 U267098 (.o(n247486),
	.a(n247484));
   no03f01 U267099 (.o(n247485),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[12]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no02m01 U267100 (.o(n253058),
	.a(n247486),
	.b(n247485));
   in01s01 U267101 (.o(n247487),
	.a(y1_bs_data[6]));
   in01s01 U267102 (.o(n247491),
	.a(n247489));
   no03f01 U267103 (.o(n247490),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[6]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no02m01 U267104 (.o(n253064),
	.a(n247491),
	.b(n247490));
   in01s01 U267105 (.o(n247492),
	.a(y1_bs_data[18]));
   na03f01 U267106 (.o(n247493),
	.a(g_swrst_r_n),
	.b(FE_OFN18_n247494),
	.c(n247492));
   no03m02 U267107 (.o(n247495),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[18]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no02m01 U267108 (.o(n253052),
	.a(n247496),
	.b(n247495));
   ao22s01 U267109 (.o(n247499),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1659]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[635]));
   ao22s01 U267110 (.o(n247498),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1403]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[379]));
   ao22s01 U267111 (.o(n247497),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1915]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[891]));
   ao22s01 U267112 (.o(n247504),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1211]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[187]));
   ao22s01 U267113 (.o(n247503),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1723]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[699]));
   ao22s01 U267114 (.o(n247502),
	.a(FE_OFN81_n248127),
	.b(regtop_dchdi_w1_hdi00[1467]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[443]));
   ao22s01 U267115 (.o(n247501),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1979]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[955]));
   ao22s01 U267116 (.o(n247508),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1275]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[251]));
   ao22s01 U267117 (.o(n247507),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1787]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[763]));
   ao22s01 U267118 (.o(n247506),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1531]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[507]));
   ao22s01 U267119 (.o(n247505),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2043]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1019]));
   ao22s01 U267120 (.o(n247514),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1083]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[59]));
   ao22s01 U267121 (.o(n247513),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1595]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[571]));
   ao22s01 U267124 (.o(n247512),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1339]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[315]));
   ao22s01 U267125 (.o(n247522),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1115]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[91]));
   ao22s01 U267126 (.o(n247521),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1627]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[603]));
   ao22s01 U267127 (.o(n247520),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1371]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[347]));
   ao22s01 U267128 (.o(n247519),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1883]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[859]));
   ao22s01 U267129 (.o(n247526),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1179]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[155]));
   ao22s01 U267130 (.o(n247525),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1691]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[667]));
   ao22s01 U267131 (.o(n247524),
	.a(FE_OFN108_n248160),
	.b(regtop_dchdi_w1_hdi00[1435]),
	.c(n247099),
	.d(regtop_dchdi_w1_hdi00[411]));
   ao22s01 U267132 (.o(n247523),
	.a(FE_OFN113_n248162),
	.b(regtop_dchdi_w1_hdi00[1947]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[923]));
   ao22s01 U267133 (.o(n247530),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1243]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[219]));
   ao22s01 U267134 (.o(n247529),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1755]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[731]));
   ao22s01 U267135 (.o(n247528),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1499]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[475]));
   ao22s01 U267136 (.o(n247527),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2011]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[987]));
   ao22s01 U267137 (.o(n247536),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1051]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[27]));
   ao22s01 U267138 (.o(n247535),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1563]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[539]));
   ao22s01 U267141 (.o(n247533),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1819]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[795]));
   na02f03 U267142 (.o(regtop_w1_hdi00_q[27]),
	.a(n247542),
	.b(FE_OFN567_n247541));
   ao22s01 U267143 (.o(n247546),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1148]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[124]));
   ao22s01 U267144 (.o(n247545),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1660]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[636]));
   ao22s01 U267145 (.o(n247544),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1404]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[380]));
   ao22s01 U267146 (.o(n247543),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1916]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[892]));
   ao22s01 U267147 (.o(n247550),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1212]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[188]));
   ao22s01 U267148 (.o(n247549),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1724]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[700]));
   ao22s01 U267149 (.o(n247548),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1468]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[444]));
   ao22s01 U267150 (.o(n247547),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1980]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[956]));
   ao22s01 U267151 (.o(n247554),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1276]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[252]));
   ao22s01 U267152 (.o(n247553),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1788]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[764]));
   ao22s01 U267153 (.o(n247552),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1532]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[508]));
   ao22f01 U267154 (.o(n247551),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2044]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1020]));
   ao22s01 U267155 (.o(n247558),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1084]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[60]));
   ao22s01 U267156 (.o(n247556),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1340]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[316]));
   ao22s01 U267157 (.o(n247555),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1852]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[828]));
   ao22f01 U267158 (.o(n247566),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1116]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[92]));
   ao22s01 U267159 (.o(n247565),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1628]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[604]));
   ao22s01 U267160 (.o(n247564),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1372]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[348]));
   ao22s01 U267161 (.o(n247563),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1884]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[860]));
   ao22s01 U267162 (.o(n247570),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1180]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[156]));
   ao22s01 U267163 (.o(n247569),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1692]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[668]));
   ao22s01 U267164 (.o(n247568),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1436]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[412]));
   ao22s01 U267165 (.o(n247567),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1948]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[924]));
   ao22s01 U267166 (.o(n247574),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1244]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[220]));
   ao22s01 U267167 (.o(n247573),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1756]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[732]));
   ao22s01 U267168 (.o(n247572),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1500]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[476]));
   ao22s01 U267169 (.o(n247571),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2012]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[988]));
   ao22s01 U267170 (.o(n247577),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1564]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[540]));
   ao22s01 U267171 (.o(n247576),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1308]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[284]));
   ao22s01 U267172 (.o(n247575),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1820]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[796]));
   na02f03 U267173 (.o(regtop_w1_hdi00_q[28]),
	.a(n247584),
	.b(n247583));
   in01s01 U267174 (.o(n247585),
	.a(y1_bs_data[2]));
   in01s01 U267175 (.o(n247589),
	.a(y1_bs_data[21]));
   no03f01 U267176 (.o(n247592),
	.a(vldtop_vld_syndec_vld_vlfeed_temporal[21]),
	.b(FE_OFN18_n247494),
	.c(n247591));
   no02f02 U267177 (.o(n247602),
	.a(n247603),
	.b(regtop_g_hclr_r_s));
   in01s01 U267178 (.o(n186690),
	.a(n247597));
   in01s01 U267179 (.o(n186689),
	.a(n247598));
   in01s01 U267180 (.o(n186691),
	.a(n247599));
   in01s01 U267181 (.o(n186687),
	.a(n247600));
   in01s01 U267182 (.o(n186686),
	.a(n247601));
   in01s01 U267183 (.o(n186688),
	.a(n247604));
   ao22s01 U267185 (.o(n247614),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1138]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[114]));
   ao22s01 U267188 (.o(n247613),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1650]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[626]));
   ao22s01 U267190 (.o(n247612),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1394]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[370]));
   ao22s01 U267193 (.o(n247611),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1906]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[882]));
   ao22s01 U267195 (.o(n247624),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1202]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[178]));
   ao22s01 U267198 (.o(n247623),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1714]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[690]));
   ao22s01 U267200 (.o(n247622),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1458]),
	.c(FE_OFN54_n247067),
	.d(regtop_dchdi_w1_hdi00[434]));
   ao22s01 U267203 (.o(n247621),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1970]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[946]));
   ao22s01 U267206 (.o(n247635),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1266]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[242]));
   ao22s01 U267209 (.o(n247634),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1778]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[754]));
   ao22s01 U267211 (.o(n247633),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1522]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[498]));
   ao22s01 U267214 (.o(n247632),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2034]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1010]));
   ao22s01 U267216 (.o(n247645),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1074]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[50]));
   ao22s01 U267219 (.o(n247644),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1586]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[562]));
   ao22s01 U267220 (.o(n247643),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1330]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[306]));
   ao22s01 U267223 (.o(n247642),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1842]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[818]));
   ao22s01 U267225 (.o(n247659),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1106]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[82]));
   ao22s01 U267228 (.o(n247658),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1618]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[594]));
   ao22s01 U267230 (.o(n247657),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1362]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[338]));
   ao22s01 U267233 (.o(n247656),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1874]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[850]));
   ao22s01 U267236 (.o(n247670),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1170]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[146]));
   ao22s01 U267238 (.o(n247669),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1682]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[658]));
   ao22s01 U267240 (.o(n247668),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1426]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[402]));
   ao22s01 U267243 (.o(n247667),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1938]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[914]));
   ao22s01 U267246 (.o(n247681),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1234]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[210]));
   ao22s01 U267249 (.o(n247680),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1746]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[722]));
   ao22s01 U267251 (.o(n247679),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1490]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[466]));
   ao22s01 U267254 (.o(n247678),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2002]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[978]));
   ao22s01 U267256 (.o(n247691),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1042]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[18]));
   ao22s01 U267258 (.o(n247690),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1554]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[530]));
   ao22s01 U267260 (.o(n247689),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1298]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[274]));
   ao22s01 U267263 (.o(n247688),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1810]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[786]));
   na02f01 U267264 (.o(regtop_w1_hdi00_q[18]),
	.a(n247697),
	.b(FE_OFN524_n247696));
   ao22s01 U267265 (.o(n247701),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1137]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[113]));
   ao22s01 U267266 (.o(n247700),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1649]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[625]));
   ao22s01 U267267 (.o(n247699),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1393]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[369]));
   ao22s01 U267268 (.o(n247698),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1905]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[881]));
   ao22f01 U267269 (.o(n247705),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1201]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[177]));
   ao22s01 U267270 (.o(n247704),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1713]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[689]));
   ao22s01 U267271 (.o(n247703),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1457]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[433]));
   ao22s01 U267272 (.o(n247702),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1969]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[945]));
   ao22s01 U267273 (.o(n247709),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1265]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[241]));
   ao22s01 U267274 (.o(n247708),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1777]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[753]));
   ao22s01 U267275 (.o(n247707),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1521]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[497]));
   ao22s01 U267276 (.o(n247706),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2033]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1009]));
   ao22s01 U267277 (.o(n247713),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1073]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[49]));
   ao22s01 U267278 (.o(n247712),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1585]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[561]));
   ao22s01 U267279 (.o(n247711),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1329]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[305]));
   ao22s01 U267280 (.o(n247710),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1841]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[817]));
   ao22s01 U267281 (.o(n247721),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1105]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[81]));
   ao22s01 U267282 (.o(n247720),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1617]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[593]));
   ao22s01 U267283 (.o(n247719),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1361]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[337]));
   ao22s01 U267284 (.o(n247718),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1873]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[849]));
   ao22s01 U267285 (.o(n247725),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1169]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[145]));
   ao22s01 U267286 (.o(n247724),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1681]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[657]));
   ao22s01 U267287 (.o(n247723),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1425]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[401]));
   ao22s01 U267288 (.o(n247722),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1937]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[913]));
   ao22s01 U267289 (.o(n247729),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1233]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[209]));
   ao22s01 U267290 (.o(n247728),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1745]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[721]));
   ao22s01 U267291 (.o(n247727),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1489]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[465]));
   ao22s01 U267292 (.o(n247726),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2001]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[977]));
   ao22s01 U267293 (.o(n247733),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1041]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[17]));
   ao22s01 U267294 (.o(n247732),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1553]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[529]));
   ao22s01 U267295 (.o(n247731),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1297]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[273]));
   ao22s01 U267296 (.o(n247730),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1809]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[785]));
   na02s01 U267297 (.o(regtop_w1_hdi00_q[17]),
	.a(n247739),
	.b(FE_OFN565_n247738));
   ao22s01 U267298 (.o(n247743),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1136]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[112]));
   ao22s01 U267299 (.o(n247742),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1648]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[624]));
   ao22s01 U267300 (.o(n247741),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1392]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[368]));
   ao22s01 U267301 (.o(n247740),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1904]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[880]));
   ao22s01 U267302 (.o(n247747),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1200]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[176]));
   ao22s01 U267303 (.o(n247746),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1712]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[688]));
   ao22s01 U267304 (.o(n247745),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1456]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[432]));
   ao22s01 U267305 (.o(n247744),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1968]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[944]));
   ao22s01 U267306 (.o(n247751),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1264]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[240]));
   ao22s01 U267307 (.o(n247750),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1776]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[752]));
   ao22s01 U267308 (.o(n247749),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1520]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[496]));
   ao22s01 U267309 (.o(n247748),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2032]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1008]));
   ao22s01 U267310 (.o(n247755),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1072]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[48]));
   ao22s01 U267311 (.o(n247754),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1584]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[560]));
   ao22s01 U267312 (.o(n247753),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1328]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[304]));
   ao22s01 U267313 (.o(n247752),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1840]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[816]));
   ao22s01 U267314 (.o(n247763),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1104]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[80]));
   ao22s01 U267315 (.o(n247762),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1616]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[592]));
   ao22s01 U267316 (.o(n247761),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1360]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[336]));
   ao22s01 U267317 (.o(n247760),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1872]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[848]));
   ao22s01 U267318 (.o(n247767),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1168]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[144]));
   ao22s01 U267319 (.o(n247766),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1680]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[656]));
   ao22s01 U267320 (.o(n247765),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1424]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[400]));
   ao22s01 U267321 (.o(n247764),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1936]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[912]));
   ao22s01 U267322 (.o(n247771),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1232]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[208]));
   ao22s01 U267323 (.o(n247770),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1744]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[720]));
   ao22s01 U267324 (.o(n247769),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1488]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[464]));
   ao22s01 U267325 (.o(n247768),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2000]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[976]));
   ao22s01 U267326 (.o(n247775),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1040]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[16]));
   ao22s01 U267327 (.o(n247774),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1552]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[528]));
   ao22s01 U267328 (.o(n247773),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1296]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[272]));
   ao22s01 U267329 (.o(n247772),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1808]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[784]));
   na02s01 U267330 (.o(regtop_w1_hdi00_q[16]),
	.a(n247781),
	.b(FE_OFN569_n247780));
   ao22s01 U267331 (.o(n247785),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1135]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[111]));
   ao22s01 U267332 (.o(n247784),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1647]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[623]));
   ao22s01 U267333 (.o(n247783),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1391]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[367]));
   ao22s01 U267334 (.o(n247782),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1903]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[879]));
   ao22s01 U267335 (.o(n247789),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1199]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[175]));
   ao22s01 U267336 (.o(n247788),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1711]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[687]));
   ao22s01 U267337 (.o(n247787),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1455]),
	.c(FE_OFN54_n247067),
	.d(regtop_dchdi_w1_hdi00[431]));
   ao22s01 U267338 (.o(n247786),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1967]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[943]));
   ao22s01 U267339 (.o(n247793),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1263]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[239]));
   ao22f01 U267340 (.o(n247792),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1775]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[751]));
   ao22s01 U267341 (.o(n247791),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1519]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[495]));
   ao22s01 U267342 (.o(n247790),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2031]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1007]));
   ao22s01 U267343 (.o(n247797),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1071]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[47]));
   ao22s01 U267344 (.o(n247796),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1583]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[559]));
   ao22f02 U267345 (.o(n247795),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1327]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[303]));
   ao22s01 U267346 (.o(n247794),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1839]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[815]));
   ao22s01 U267347 (.o(n247805),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1103]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[79]));
   ao22s01 U267348 (.o(n247804),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1615]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[591]));
   ao22s01 U267349 (.o(n247803),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1359]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[335]));
   ao22s01 U267350 (.o(n247802),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1871]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[847]));
   ao22s01 U267351 (.o(n247809),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1167]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[143]));
   ao22s01 U267352 (.o(n247808),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1679]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[655]));
   ao22s01 U267353 (.o(n247807),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1423]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[399]));
   ao22s01 U267354 (.o(n247806),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1935]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[911]));
   ao22s01 U267355 (.o(n247813),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1231]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[207]));
   ao22f01 U267356 (.o(n247812),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1743]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[719]));
   ao22s01 U267357 (.o(n247811),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1487]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[463]));
   ao22s01 U267358 (.o(n247810),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1999]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[975]));
   ao22s01 U267359 (.o(n247817),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1039]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[15]));
   ao22s01 U267360 (.o(n247816),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1551]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[527]));
   ao22s01 U267361 (.o(n247815),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1295]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[271]));
   ao22s01 U267362 (.o(n247814),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1807]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[783]));
   na02f03 U267363 (.o(regtop_w1_hdi00_q[15]),
	.a(n247823),
	.b(n247822));
   ao22s01 U267364 (.o(n247827),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1143]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[119]));
   ao22s01 U267365 (.o(n247826),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1655]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[631]));
   ao22s01 U267366 (.o(n247825),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1399]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[375]));
   ao22s01 U267367 (.o(n247824),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1911]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[887]));
   ao22s01 U267368 (.o(n247831),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1207]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[183]));
   ao22s01 U267369 (.o(n247830),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1719]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[695]));
   ao22s01 U267370 (.o(n247829),
	.a(FE_OFN81_n248127),
	.b(regtop_dchdi_w1_hdi00[1463]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[439]));
   ao22s01 U267371 (.o(n247828),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1975]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[951]));
   ao22s01 U267372 (.o(n247835),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1271]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[247]));
   ao22s01 U267373 (.o(n247834),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1783]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[759]));
   ao22s01 U267374 (.o(n247833),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1527]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[503]));
   ao22s01 U267375 (.o(n247832),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2039]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1015]));
   ao22f01 U267376 (.o(n247839),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1079]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[55]));
   ao22s01 U267377 (.o(n247838),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1591]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[567]));
   ao22s01 U267378 (.o(n247837),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1335]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[311]));
   ao22f02 U267379 (.o(n247836),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1847]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[823]));
   ao22s01 U267380 (.o(n247847),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1111]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[87]));
   ao22s01 U267381 (.o(n247846),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1623]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[599]));
   ao22s01 U267382 (.o(n247845),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1367]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[343]));
   ao22s01 U267383 (.o(n247844),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1879]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[855]));
   ao22s01 U267384 (.o(n247851),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1175]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[151]));
   ao22s01 U267385 (.o(n247850),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1687]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[663]));
   ao22s01 U267386 (.o(n247849),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1431]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[407]));
   ao22s01 U267387 (.o(n247848),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1943]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[919]));
   ao22s01 U267388 (.o(n247855),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1239]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[215]));
   ao22s01 U267389 (.o(n247854),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1751]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[727]));
   ao22f01 U267390 (.o(n247853),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1495]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[471]));
   ao22s01 U267391 (.o(n247852),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2007]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[983]));
   ao22s01 U267392 (.o(n247859),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1047]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[23]));
   ao22s01 U267393 (.o(n247858),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1559]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[535]));
   ao22s01 U267394 (.o(n247857),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1303]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[279]));
   ao22s01 U267395 (.o(n247856),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1815]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[791]));
   na02f03 U267396 (.o(regtop_w1_hdi00_q[23]),
	.a(n247865),
	.b(n247864));
   ao22s01 U267397 (.o(n247869),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1134]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[110]));
   ao22s01 U267398 (.o(n247868),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1646]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[622]));
   ao22s01 U267399 (.o(n247867),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1390]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[366]));
   ao22s01 U267400 (.o(n247866),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1902]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[878]));
   ao22s01 U267401 (.o(n247873),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1198]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[174]));
   ao22s01 U267402 (.o(n247872),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1710]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[686]));
   ao22s01 U267403 (.o(n247871),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1454]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[430]));
   ao22s01 U267404 (.o(n247870),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1966]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[942]));
   ao22s01 U267405 (.o(n247877),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1262]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[238]));
   ao22f01 U267406 (.o(n247876),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1774]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[750]));
   ao22f01 U267407 (.o(n247875),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1518]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[494]));
   ao22s01 U267408 (.o(n247881),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1070]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[46]));
   ao22f01 U267409 (.o(n247880),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1582]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[558]));
   ao22s01 U267410 (.o(n247879),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1326]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[302]));
   ao22s01 U267411 (.o(n247878),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1838]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[814]));
   ao22s01 U267412 (.o(n247889),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1102]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[78]));
   ao22f01 U267413 (.o(n247888),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1614]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[590]));
   ao22s01 U267414 (.o(n247887),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1358]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[334]));
   ao22s01 U267415 (.o(n247886),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1870]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[846]));
   ao22s01 U267416 (.o(n247893),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1166]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[142]));
   ao22s01 U267417 (.o(n247892),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1678]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[654]));
   ao22s01 U267418 (.o(n247891),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1422]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[398]));
   ao22s01 U267419 (.o(n247890),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1934]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[910]));
   ao22s01 U267420 (.o(n247897),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1230]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[206]));
   ao22s01 U267421 (.o(n247896),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1742]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[718]));
   ao22s01 U267422 (.o(n247895),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1486]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[462]));
   ao22s01 U267423 (.o(n247894),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1998]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[974]));
   ao22s01 U267424 (.o(n247901),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1038]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[14]));
   ao22s01 U267425 (.o(n247900),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1550]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[526]));
   ao22s01 U267426 (.o(n247899),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1294]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[270]));
   ao22s01 U267427 (.o(n247898),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1806]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[782]));
   na02f02 U267428 (.o(regtop_w1_hdi00_q[14]),
	.a(n247907),
	.b(n247906));
   ao22s01 U267429 (.o(n247911),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1133]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[109]));
   ao22s01 U267430 (.o(n247910),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1645]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[621]));
   ao22s01 U267431 (.o(n247909),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1389]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[365]));
   ao22s01 U267432 (.o(n247908),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1901]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[877]));
   ao22s01 U267433 (.o(n247915),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1197]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[173]));
   ao22s01 U267434 (.o(n247914),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1709]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[685]));
   ao22s01 U267435 (.o(n247913),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1453]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[429]));
   ao22s01 U267436 (.o(n247912),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1965]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[941]));
   ao22f01 U267437 (.o(n247919),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1261]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[237]));
   ao22s01 U267438 (.o(n247918),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1773]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[749]));
   ao22s01 U267439 (.o(n247917),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1517]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[493]));
   ao22s01 U267440 (.o(n247916),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2029]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1005]));
   ao22s01 U267441 (.o(n247923),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1069]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[45]));
   ao22s01 U267442 (.o(n247921),
	.a(n248139),
	.b(regtop_dchdi_w1_hdi00[1325]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[301]));
   ao22s01 U267443 (.o(n247920),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1837]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[813]));
   ao22s01 U267444 (.o(n247931),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1101]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[77]));
   ao22s01 U267445 (.o(n247930),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1613]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[589]));
   ao22s01 U267446 (.o(n247929),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1357]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[333]));
   ao22s01 U267447 (.o(n247928),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1869]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[845]));
   ao22s01 U267448 (.o(n247935),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1165]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[141]));
   ao22s01 U267449 (.o(n247934),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1677]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[653]));
   ao22s01 U267450 (.o(n247933),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1421]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[397]));
   ao22s01 U267451 (.o(n247932),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1933]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[909]));
   ao22s01 U267452 (.o(n247939),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1229]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[205]));
   ao22s01 U267453 (.o(n247938),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1741]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[717]));
   ao22s01 U267454 (.o(n247937),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1485]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[461]));
   ao22s01 U267455 (.o(n247936),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1997]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[973]));
   ao22s01 U267456 (.o(n247942),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1549]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[525]));
   ao22s01 U267457 (.o(n247941),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1293]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[269]));
   ao22s01 U267458 (.o(n247940),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1805]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[781]));
   na02f03 U267459 (.o(regtop_w1_hdi00_q[13]),
	.a(n247949),
	.b(n247948));
   ao22s01 U267460 (.o(n247953),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1139]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[115]));
   ao22s01 U267461 (.o(n247952),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1651]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[627]));
   ao22s01 U267462 (.o(n247951),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1395]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[371]));
   ao22s01 U267463 (.o(n247950),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1907]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[883]));
   ao22s01 U267464 (.o(n247957),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1203]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[179]));
   ao22s01 U267465 (.o(n247956),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1715]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[691]));
   ao22s01 U267466 (.o(n247955),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1459]),
	.c(FE_OFN54_n247067),
	.d(regtop_dchdi_w1_hdi00[435]));
   ao22s01 U267467 (.o(n247954),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1971]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[947]));
   ao22s01 U267468 (.o(n247961),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1267]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[243]));
   ao22s01 U267469 (.o(n247960),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1779]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[755]));
   ao22s01 U267470 (.o(n247959),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1523]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[499]));
   ao22s01 U267471 (.o(n247958),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2035]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1011]));
   ao22s01 U267472 (.o(n247965),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1075]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[51]));
   ao22s01 U267473 (.o(n247964),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1587]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[563]));
   ao22s01 U267474 (.o(n247963),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1331]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[307]));
   ao22s01 U267475 (.o(n247962),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1843]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[819]));
   ao22s01 U267476 (.o(n247973),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1107]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[83]));
   ao22s01 U267477 (.o(n247972),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1619]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[595]));
   ao22s01 U267478 (.o(n247971),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1363]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[339]));
   ao22s01 U267479 (.o(n247970),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1875]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[851]));
   ao22s01 U267480 (.o(n247977),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1171]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[147]));
   ao22s01 U267481 (.o(n247976),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1683]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[659]));
   ao22s01 U267482 (.o(n247975),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1427]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[403]));
   ao22s01 U267483 (.o(n247974),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1939]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[915]));
   ao22s01 U267484 (.o(n247981),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1235]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[211]));
   ao22s01 U267485 (.o(n247980),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1747]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[723]));
   ao22s01 U267486 (.o(n247979),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1491]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[467]));
   ao22s01 U267487 (.o(n247978),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2003]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[979]));
   ao22f01 U267488 (.o(n247985),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1043]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[19]));
   ao22f02 U267489 (.o(n247984),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1555]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[531]));
   ao22f01 U267490 (.o(n247983),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1299]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[275]));
   ao22s01 U267491 (.o(n247982),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1811]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[787]));
   na02f01 U267492 (.o(regtop_w1_hdi00_q[19]),
	.a(n247991),
	.b(n247990));
   ao22s01 U267493 (.o(n247995),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1122]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[98]));
   ao22s01 U267494 (.o(n247994),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1634]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[610]));
   ao22s01 U267495 (.o(n247993),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1378]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[354]));
   ao22s01 U267496 (.o(n247992),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1890]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[866]));
   ao22s01 U267497 (.o(n247999),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1186]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[162]));
   ao22s01 U267498 (.o(n247997),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1442]),
	.c(FE_OFN54_n247067),
	.d(regtop_dchdi_w1_hdi00[418]));
   ao22s01 U267499 (.o(n247996),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1954]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[930]));
   ao22s01 U267500 (.o(n248003),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1250]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[226]));
   ao22s01 U267501 (.o(n248002),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1762]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[738]));
   ao22s01 U267502 (.o(n248001),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1506]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[482]));
   ao22s01 U267503 (.o(n248000),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2018]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[994]));
   ao22s01 U267504 (.o(n248007),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1058]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[34]));
   ao22s01 U267505 (.o(n248006),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1570]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[546]));
   ao22s01 U267506 (.o(n248005),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1314]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[290]));
   ao22s01 U267507 (.o(n248004),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1826]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[802]));
   ao22s01 U267508 (.o(n248015),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1090]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[66]));
   ao22s01 U267509 (.o(n248014),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1602]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[578]));
   ao22s01 U267510 (.o(n248013),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1346]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[322]));
   ao22s01 U267511 (.o(n248012),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1858]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[834]));
   ao22s01 U267512 (.o(n248018),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1666]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[642]));
   ao22s01 U267513 (.o(n248017),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1410]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[386]));
   ao22s01 U267514 (.o(n248016),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1922]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[898]));
   ao22s01 U267515 (.o(n248023),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1218]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[194]));
   ao22f01 U267516 (.o(n248022),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1730]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[706]));
   ao22s01 U267517 (.o(n248021),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1474]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[450]));
   ao22s01 U267518 (.o(n248020),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1986]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[962]));
   ao22s01 U267519 (.o(n248027),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1026]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[2]));
   ao22f01 U267520 (.o(n248026),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1538]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[514]));
   ao22s01 U267521 (.o(n248025),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1282]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[258]));
   ao22s01 U267522 (.o(n248024),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1794]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[770]));
   na02s01 U267523 (.o(regtop_w1_hdi00_q[2]),
	.a(n248033),
	.b(n248032));
   ao22s01 U267524 (.o(n248037),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1131]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[107]));
   ao22s01 U267525 (.o(n248036),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1643]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[619]));
   ao22s01 U267526 (.o(n248035),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1387]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[363]));
   ao22s01 U267527 (.o(n248034),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1899]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[875]));
   ao22f01 U267528 (.o(n248041),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1195]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[171]));
   ao22s01 U267529 (.o(n248040),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1707]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[683]));
   ao22s01 U267530 (.o(n248039),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1451]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[427]));
   ao22s01 U267531 (.o(n248038),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1963]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[939]));
   ao22f01 U267532 (.o(n248045),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1259]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[235]));
   ao22s01 U267533 (.o(n248044),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1771]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[747]));
   ao22s01 U267534 (.o(n248043),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1515]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[491]));
   ao22s01 U267535 (.o(n248042),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2027]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1003]));
   ao22s01 U267536 (.o(n248049),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1067]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[43]));
   ao22s01 U267537 (.o(n248048),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1579]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[555]));
   ao22s01 U267538 (.o(n248047),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1323]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[299]));
   ao22s01 U267539 (.o(n248046),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1835]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[811]));
   ao22s01 U267540 (.o(n248057),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1099]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[75]));
   ao22s01 U267541 (.o(n248055),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1355]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[331]));
   ao22s01 U267542 (.o(n248054),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1867]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[843]));
   ao22s01 U267543 (.o(n248061),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1163]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[139]));
   ao22s01 U267544 (.o(n248060),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1675]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[651]));
   ao22s01 U267545 (.o(n248059),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1419]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[395]));
   ao22s01 U267546 (.o(n248058),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1931]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[907]));
   ao22s01 U267547 (.o(n248065),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1227]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[203]));
   ao22s01 U267548 (.o(n248064),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1739]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[715]));
   ao22s01 U267549 (.o(n248063),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1483]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[459]));
   ao22s01 U267550 (.o(n248062),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1995]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[971]));
   ao22s01 U267551 (.o(n248069),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1035]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[11]));
   ao22s01 U267552 (.o(n248068),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1547]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[523]));
   ao22s01 U267553 (.o(n248067),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1291]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[267]));
   ao22s01 U267554 (.o(n248066),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1803]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[779]));
   na02f01 U267555 (.o(regtop_w1_hdi00_q[11]),
	.a(n248075),
	.b(FE_OFN571_n248074));
   ao22s01 U267556 (.o(n248079),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1130]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[106]));
   ao22s01 U267557 (.o(n248078),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1642]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[618]));
   ao22s01 U267558 (.o(n248077),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1386]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[362]));
   ao22s01 U267559 (.o(n248076),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1898]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[874]));
   ao22s01 U267560 (.o(n248082),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1706]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[682]));
   ao22s01 U267561 (.o(n248081),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1450]),
	.c(FE_OFN54_n247067),
	.d(regtop_dchdi_w1_hdi00[426]));
   ao22s01 U267562 (.o(n248080),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1962]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[938]));
   ao22s01 U267563 (.o(n248087),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1258]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[234]));
   ao22s01 U267564 (.o(n248086),
	.a(FE_OFN146_n248372),
	.b(regtop_dchdi_w1_hdi00[1770]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[746]));
   ao22s01 U267565 (.o(n248085),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1514]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[490]));
   ao22s01 U267566 (.o(n248084),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2026]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1002]));
   ao22s01 U267567 (.o(n248091),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1066]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[42]));
   ao22s01 U267568 (.o(n248090),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1578]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[554]));
   ao22s01 U267569 (.o(n248089),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1322]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[298]));
   ao22s01 U267570 (.o(n248088),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1834]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[810]));
   ao22s01 U267571 (.o(n248099),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1098]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[74]));
   ao22s01 U267572 (.o(n248098),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1610]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[586]));
   ao22s01 U267573 (.o(n248097),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1354]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[330]));
   ao22s01 U267574 (.o(n248103),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1162]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[138]));
   ao22s01 U267575 (.o(n248102),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1674]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[650]));
   ao22s01 U267576 (.o(n248101),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1418]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[394]));
   ao22s01 U267577 (.o(n248100),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1930]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[906]));
   ao22s01 U267578 (.o(n248107),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1226]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[202]));
   ao22s01 U267579 (.o(n248106),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1738]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[714]));
   ao22f02 U267580 (.o(n248105),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1482]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[458]));
   ao22s01 U267581 (.o(n248104),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1994]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[970]));
   ao22s01 U267582 (.o(n248111),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1034]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[10]));
   ao22s01 U267583 (.o(n248110),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1546]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[522]));
   ao22s01 U267584 (.o(n248109),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1290]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[266]));
   ao22s01 U267585 (.o(n248108),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1802]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[778]));
   na02f02 U267586 (.o(regtop_w1_hdi00_q[10]),
	.a(n248117),
	.b(n248116));
   ao22s01 U267587 (.o(n248125),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1149]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[125]));
   ao22s01 U267588 (.o(n248124),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1661]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[637]));
   ao22s01 U267589 (.o(n248123),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1405]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[381]));
   ao22s01 U267590 (.o(n248122),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1917]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[893]));
   ao22s01 U267591 (.o(n248133),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1213]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[189]));
   ao22s01 U267592 (.o(n248132),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1725]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[701]));
   ao22s01 U267593 (.o(n248131),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1469]),
	.c(FE_OFN54_n247067),
	.d(regtop_dchdi_w1_hdi00[445]));
   ao22s01 U267594 (.o(n248130),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1981]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[957]));
   ao22s01 U267595 (.o(n248137),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1277]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[253]));
   ao22s01 U267596 (.o(n248136),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1789]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[765]));
   ao22s01 U267597 (.o(n248135),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1533]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[509]));
   ao22s01 U267598 (.o(n248134),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2045]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1021]));
   ao22s01 U267599 (.o(n248145),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1085]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[61]));
   ao22s01 U267600 (.o(n248144),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1597]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[573]));
   ao22s01 U267601 (.o(n248143),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1341]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[317]));
   ao22s01 U267602 (.o(n248142),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1853]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[829]));
   ao22s01 U267603 (.o(n248157),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1117]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[93]));
   ao22s01 U267604 (.o(n248156),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1629]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[605]));
   ao22s01 U267605 (.o(n248155),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1373]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[349]));
   ao22s01 U267606 (.o(n248154),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1885]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[861]));
   ao22s01 U267607 (.o(n248166),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1181]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[157]));
   ao22s01 U267608 (.o(n248165),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1693]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[669]));
   ao22s01 U267609 (.o(n248164),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1437]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[413]));
   ao22s01 U267610 (.o(n248163),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1949]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[925]));
   ao22s01 U267611 (.o(n248172),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1245]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[221]));
   ao22f01 U267612 (.o(n248171),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1757]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[733]));
   ao22f01 U267613 (.o(n248170),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1501]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[477]));
   ao22s01 U267614 (.o(n248169),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2013]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[989]));
   ao22s01 U267615 (.o(n248180),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1053]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[29]));
   ao22s01 U267616 (.o(n248179),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1565]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[541]));
   ao22s01 U267617 (.o(n248178),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1309]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[285]));
   ao22s01 U267618 (.o(n248177),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1821]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[797]));
   na02f03 U267619 (.o(regtop_w1_hdi00_q[29]),
	.a(n248186),
	.b(n248185));
   ao22s01 U267620 (.o(n248190),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1120]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[96]));
   ao22s01 U267621 (.o(n248189),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1632]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[608]));
   ao22s01 U267622 (.o(n248188),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1376]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[352]));
   ao22s01 U267623 (.o(n248187),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1888]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[864]));
   ao22s01 U267624 (.o(n248194),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1184]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[160]));
   ao22s01 U267625 (.o(n248193),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1696]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[672]));
   ao22s01 U267626 (.o(n248192),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1440]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[416]));
   ao22s01 U267627 (.o(n248191),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1952]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[928]));
   ao22s01 U267628 (.o(n248198),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1248]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[224]));
   ao22s01 U267629 (.o(n248196),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1504]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[480]));
   ao22s01 U267630 (.o(n248195),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2016]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[992]));
   ao22s01 U267631 (.o(n248202),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1056]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[32]));
   ao22s01 U267632 (.o(n248201),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1568]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[544]));
   ao22s01 U267633 (.o(n248200),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1312]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[288]));
   ao22s01 U267634 (.o(n248199),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1824]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[800]));
   ao22f01 U267635 (.o(n248210),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1088]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[64]));
   ao22s01 U267636 (.o(n248209),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1600]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[576]));
   ao22s01 U267637 (.o(n248208),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1344]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[320]));
   ao22s01 U267638 (.o(n248207),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1856]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[832]));
   ao22s01 U267639 (.o(n248214),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1152]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[128]));
   ao22s01 U267640 (.o(n248213),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1664]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[640]));
   ao22s01 U267641 (.o(n248212),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1408]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[384]));
   ao22s01 U267642 (.o(n248211),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1920]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[896]));
   ao22f01 U267643 (.o(n248217),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1728]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[704]));
   ao22s01 U267644 (.o(n248216),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1472]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[448]));
   ao22s01 U267645 (.o(n248215),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1984]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[960]));
   ao22s01 U267646 (.o(n248222),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1024]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[0]));
   ao22s01 U267647 (.o(n248221),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1536]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[512]));
   ao22s01 U267648 (.o(n248220),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1280]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[256]));
   ao22s01 U267649 (.o(n248219),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1792]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[768]));
   na02f03 U267650 (.o(regtop_w1_hdi00_q[0]),
	.a(n248228),
	.b(n248227));
   ao22s01 U267651 (.o(n248232),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1150]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[126]));
   ao22s01 U267652 (.o(n248231),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1662]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[638]));
   ao22s01 U267653 (.o(n248230),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1406]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[382]));
   ao22s01 U267654 (.o(n248229),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1918]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[894]));
   ao22m02 U267655 (.o(n248236),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1214]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[190]));
   ao22s01 U267656 (.o(n248235),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1726]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[702]));
   ao22s01 U267657 (.o(n248234),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1470]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[446]));
   ao22s01 U267658 (.o(n248233),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1982]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[958]));
   ao22s01 U267659 (.o(n248240),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1278]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[254]));
   ao22s01 U267660 (.o(n248239),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1790]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[766]));
   ao22s01 U267661 (.o(n248238),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1534]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[510]));
   ao22f01 U267662 (.o(n248237),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2046]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1022]));
   ao22s01 U267663 (.o(n248244),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1086]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[62]));
   ao22s01 U267664 (.o(n248243),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1598]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[574]));
   ao22s01 U267665 (.o(n248242),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1342]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[318]));
   ao22s01 U267666 (.o(n248241),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1854]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[830]));
   ao22s01 U267667 (.o(n248252),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1118]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[94]));
   ao22s01 U267668 (.o(n248251),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1630]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[606]));
   ao22s01 U267669 (.o(n248250),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1374]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[350]));
   ao22s01 U267670 (.o(n248249),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1886]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[862]));
   ao22s01 U267671 (.o(n248256),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1182]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[158]));
   ao22s01 U267672 (.o(n248255),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1694]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[670]));
   ao22s01 U267673 (.o(n248254),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1438]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[414]));
   ao22s01 U267674 (.o(n248253),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1950]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[926]));
   ao22s01 U267675 (.o(n248260),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1246]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[222]));
   ao22s01 U267676 (.o(n248259),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1758]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[734]));
   ao22f02 U267677 (.o(n248258),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1502]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[478]));
   ao22s01 U267678 (.o(n248257),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2014]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[990]));
   ao22s01 U267679 (.o(n248264),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1054]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[30]));
   ao22s01 U267680 (.o(n248263),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1566]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[542]));
   ao22s01 U267681 (.o(n248262),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1310]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[286]));
   ao22s01 U267682 (.o(n248261),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1822]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[798]));
   na02f01 U267683 (.o(regtop_w1_hdi00_q[30]),
	.a(n248270),
	.b(n248269));
   ao22s01 U267684 (.o(n248274),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1142]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[118]));
   ao22s01 U267685 (.o(n248273),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1654]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[630]));
   ao22s01 U267686 (.o(n248272),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1398]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[374]));
   ao22s01 U267687 (.o(n248271),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1910]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[886]));
   ao22f01 U267688 (.o(n248278),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1206]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[182]));
   ao22s01 U267689 (.o(n248277),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1718]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[694]));
   ao22s01 U267690 (.o(n248276),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1462]),
	.c(FE_OFN54_n247067),
	.d(regtop_dchdi_w1_hdi00[438]));
   ao22s01 U267691 (.o(n248275),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1974]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[950]));
   ao22s01 U267692 (.o(n248282),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1270]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[246]));
   ao22s01 U267693 (.o(n248281),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1782]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[758]));
   ao22s01 U267694 (.o(n248280),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1526]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[502]));
   ao22s01 U267695 (.o(n248279),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2038]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1014]));
   ao22s01 U267696 (.o(n248286),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1078]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[54]));
   ao22s01 U267697 (.o(n248285),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1590]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[566]));
   ao22s01 U267698 (.o(n248284),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1334]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[310]));
   ao22s01 U267699 (.o(n248283),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1846]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[822]));
   ao22s01 U267700 (.o(n248294),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1110]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[86]));
   ao22s01 U267701 (.o(n248293),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1622]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[598]));
   ao22s01 U267702 (.o(n248292),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1366]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[342]));
   ao22s01 U267703 (.o(n248291),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1878]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[854]));
   ao22s01 U267704 (.o(n248298),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1174]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[150]));
   ao22s01 U267705 (.o(n248297),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1686]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[662]));
   ao22s01 U267706 (.o(n248296),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1430]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[406]));
   ao22s01 U267707 (.o(n248295),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1942]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[918]));
   ao22s01 U267708 (.o(n248302),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1238]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[214]));
   ao22s01 U267709 (.o(n248301),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1750]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[726]));
   ao22s01 U267710 (.o(n248300),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1494]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[470]));
   ao22s01 U267711 (.o(n248299),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2006]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[982]));
   ao22s01 U267712 (.o(n248306),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1046]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[22]));
   ao22s01 U267713 (.o(n248305),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1558]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[534]));
   ao22s01 U267714 (.o(n248304),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1302]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[278]));
   ao22s01 U267715 (.o(n248303),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1814]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[790]));
   na02f02 U267716 (.o(regtop_w1_hdi00_q[22]),
	.a(n248312),
	.b(FE_OFN374_n248311));
   ao22s01 U267717 (.o(n248316),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1127]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[103]));
   ao22s01 U267718 (.o(n248315),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1639]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[615]));
   ao22s01 U267719 (.o(n248314),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1383]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[359]));
   ao22s01 U267720 (.o(n248313),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1895]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[871]));
   ao22s01 U267721 (.o(n248320),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1191]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[167]));
   ao22s01 U267722 (.o(n248319),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1703]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[679]));
   ao22s01 U267723 (.o(n248318),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1447]),
	.c(FE_OFN54_n247067),
	.d(regtop_dchdi_w1_hdi00[423]));
   ao22s01 U267724 (.o(n248317),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1959]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[935]));
   ao22s01 U267725 (.o(n248324),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1255]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[231]));
   ao22f06 U267726 (.o(n248323),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1767]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[743]));
   ao22s01 U267727 (.o(n248322),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1511]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[487]));
   ao22f04 U267728 (.o(n248321),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2023]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[999]));
   ao22s01 U267729 (.o(n248328),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1063]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[39]));
   ao22s01 U267730 (.o(n248327),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1575]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[551]));
   ao22s01 U267731 (.o(n248326),
	.a(n248139),
	.b(regtop_dchdi_w1_hdi00[1319]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[295]));
   ao22s01 U267732 (.o(n248325),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1831]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[807]));
   ao22s01 U267733 (.o(n248336),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1095]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[71]));
   ao22s01 U267734 (.o(n248335),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1607]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[583]));
   ao22s01 U267735 (.o(n248334),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1351]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[327]));
   ao22s01 U267736 (.o(n248333),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1863]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[839]));
   ao22s01 U267737 (.o(n248340),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1159]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[135]));
   ao22s01 U267738 (.o(n248339),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1671]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[647]));
   ao22s01 U267739 (.o(n248338),
	.a(FE_OFN108_n248160),
	.b(regtop_dchdi_w1_hdi00[1415]),
	.c(n247099),
	.d(regtop_dchdi_w1_hdi00[391]));
   ao22s01 U267740 (.o(n248337),
	.a(FE_OFN113_n248162),
	.b(regtop_dchdi_w1_hdi00[1927]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[903]));
   ao22s01 U267741 (.o(n248344),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1223]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[199]));
   ao22s01 U267742 (.o(n248342),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1479]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[455]));
   ao22s01 U267743 (.o(n248341),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1991]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[967]));
   ao22f01 U267744 (.o(n248348),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1031]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[7]));
   ao22s01 U267745 (.o(n248347),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1543]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[519]));
   ao22s01 U267746 (.o(n248346),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1287]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[263]));
   ao22s01 U267747 (.o(n248345),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1799]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[775]));
   na02f02 U267748 (.o(regtop_w1_hdi00_q[7]),
	.a(n248354),
	.b(n248353));
   ao22s01 U267749 (.o(n248361),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1144]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[120]));
   ao22s01 U267750 (.o(n248360),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1656]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[632]));
   ao22s01 U267751 (.o(n248359),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1400]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[376]));
   ao22s01 U267752 (.o(n248358),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1912]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[888]));
   ao22s01 U267753 (.o(n248368),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1208]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[184]));
   ao22s01 U267754 (.o(n248367),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1720]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[696]));
   ao22s01 U267755 (.o(n248366),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1464]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[440]));
   ao22s01 U267756 (.o(n248365),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1976]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[952]));
   ao22s01 U267757 (.o(n248379),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1272]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[248]));
   ao22s01 U267758 (.o(n248378),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1784]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[760]));
   ao22s01 U267759 (.o(n248377),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1528]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[504]));
   ao22s01 U267760 (.o(n248376),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2040]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1016]));
   ao22s01 U267761 (.o(n248386),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1080]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[56]));
   ao22s01 U267762 (.o(n248385),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1592]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[568]));
   ao22s01 U267763 (.o(n248384),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1336]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[312]));
   ao22s01 U267764 (.o(n248383),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1848]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[824]));
   ao22s01 U267765 (.o(n248397),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1112]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[88]));
   ao22s01 U267766 (.o(n248396),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1624]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[600]));
   ao22s01 U267767 (.o(n248395),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1368]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[344]));
   ao22s01 U267768 (.o(n248394),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1880]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[856]));
   ao22s01 U267769 (.o(n248403),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1176]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[152]));
   ao22s01 U267770 (.o(n248401),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1432]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[408]));
   ao22s01 U267771 (.o(n248400),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1944]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[920]));
   ao22s01 U267772 (.o(n248412),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1240]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[216]));
   ao22s01 U267773 (.o(n248411),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1752]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[728]));
   ao22s01 U267774 (.o(n248410),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1496]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[472]));
   ao22s01 U267775 (.o(n248409),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2008]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[984]));
   ao22s01 U267776 (.o(n248419),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1048]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[24]));
   ao22s01 U267777 (.o(n248418),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1560]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[536]));
   ao22s01 U267778 (.o(n248417),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1304]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[280]));
   ao22s01 U267779 (.o(n248416),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1816]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[792]));
   na02f03 U267780 (.o(regtop_w1_hdi00_q[24]),
	.a(n248425),
	.b(FE_OFN542_n248424));
   ao22s01 U267781 (.o(n248428),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1644]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[620]));
   ao22s01 U267782 (.o(n248427),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1388]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[364]));
   ao22s01 U267783 (.o(n248426),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1900]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[876]));
   ao22s01 U267784 (.o(n248433),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1196]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[172]));
   ao22f02 U267785 (.o(n248432),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1708]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[684]));
   ao22s01 U267786 (.o(n248431),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1452]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[428]));
   ao22s01 U267787 (.o(n248430),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1964]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[940]));
   ao22s01 U267788 (.o(n248437),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1260]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[236]));
   ao22s01 U267789 (.o(n248436),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1772]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[748]));
   ao22s01 U267790 (.o(n248435),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1516]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[492]));
   ao22s01 U267791 (.o(n248434),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2028]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1004]));
   ao22s01 U267792 (.o(n248441),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1068]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[44]));
   ao22s01 U267793 (.o(n248440),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1580]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[556]));
   ao22s01 U267794 (.o(n248439),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1324]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[300]));
   ao22s01 U267795 (.o(n248449),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1100]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[76]));
   ao22s01 U267796 (.o(n248448),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1612]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[588]));
   ao22s01 U267797 (.o(n248447),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1356]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[332]));
   ao22s01 U267798 (.o(n248446),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1868]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[844]));
   ao22s01 U267799 (.o(n248453),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1164]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[140]));
   ao22s01 U267800 (.o(n248452),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1676]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[652]));
   ao22s01 U267801 (.o(n248451),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1420]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[396]));
   ao22s01 U267802 (.o(n248450),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1932]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[908]));
   ao22s01 U267803 (.o(n248457),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1228]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[204]));
   ao22s01 U267804 (.o(n248456),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1740]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[716]));
   ao22s01 U267805 (.o(n248455),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1484]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[460]));
   ao22s01 U267806 (.o(n248454),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1996]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[972]));
   ao22s01 U267807 (.o(n248461),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1036]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[12]));
   ao22s01 U267808 (.o(n248460),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1548]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[524]));
   ao22s01 U267809 (.o(n248458),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1804]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[780]));
   na02f01 U267810 (.o(regtop_w1_hdi00_q[12]),
	.a(n248467),
	.b(n248466));
   ao22s01 U267811 (.o(n248471),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1140]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[116]));
   ao22s01 U267812 (.o(n248470),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1652]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[628]));
   ao22s01 U267813 (.o(n248469),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1396]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[372]));
   ao22s01 U267814 (.o(n248468),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1908]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[884]));
   ao22s01 U267815 (.o(n248475),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1204]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[180]));
   ao22s01 U267816 (.o(n248474),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1716]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[692]));
   ao22s01 U267817 (.o(n248473),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1460]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[436]));
   ao22s01 U267818 (.o(n248472),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1972]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[948]));
   ao22s01 U267819 (.o(n248479),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1268]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[244]));
   ao22s01 U267820 (.o(n248478),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1780]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[756]));
   ao22s01 U267821 (.o(n248477),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1524]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[500]));
   ao22f01 U267822 (.o(n248476),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2036]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1012]));
   ao22s01 U267823 (.o(n248483),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1076]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[52]));
   ao22s01 U267824 (.o(n248482),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1588]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[564]));
   ao22s01 U267825 (.o(n248480),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1844]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[820]));
   ao22s01 U267826 (.o(n248491),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1108]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[84]));
   ao22s01 U267827 (.o(n248490),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1620]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[596]));
   ao22s01 U267828 (.o(n248489),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1364]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[340]));
   ao22s01 U267829 (.o(n248488),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1876]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[852]));
   ao22s01 U267830 (.o(n248495),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1172]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[148]));
   ao22s01 U267831 (.o(n248494),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1684]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[660]));
   ao22s01 U267832 (.o(n248493),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1428]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[404]));
   ao22s01 U267833 (.o(n248492),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1940]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[916]));
   ao22s01 U267834 (.o(n248499),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1236]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[212]));
   ao22s01 U267835 (.o(n248498),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1748]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[724]));
   ao22s01 U267836 (.o(n248497),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1492]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[468]));
   ao22s01 U267837 (.o(n248496),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2004]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[980]));
   ao22s01 U267838 (.o(n248503),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1044]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[20]));
   ao22s01 U267839 (.o(n248502),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1556]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[532]));
   ao22s01 U267840 (.o(n248501),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1300]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[276]));
   ao22s01 U267841 (.o(n248500),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1812]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[788]));
   ao22s01 U267842 (.o(n248513),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1123]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[99]));
   ao22s01 U267843 (.o(n248512),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1635]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[611]));
   ao22s01 U267844 (.o(n248511),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1379]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[355]));
   ao22s01 U267845 (.o(n248517),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1187]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[163]));
   ao22s01 U267846 (.o(n248516),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1699]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[675]));
   ao22s01 U267847 (.o(n248515),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1443]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[419]));
   ao22s01 U267848 (.o(n248514),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1955]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[931]));
   ao22s01 U267849 (.o(n248521),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1251]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[227]));
   ao22s01 U267850 (.o(n248520),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1763]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[739]));
   ao22s01 U267851 (.o(n248519),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1507]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[483]));
   ao22s01 U267852 (.o(n248518),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2019]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[995]));
   ao22s01 U267853 (.o(n248525),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1059]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[35]));
   ao22s01 U267854 (.o(n248524),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1571]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[547]));
   ao22s01 U267855 (.o(n248523),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1315]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[291]));
   ao22s01 U267856 (.o(n248522),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1827]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[803]));
   ao22s01 U267857 (.o(n248533),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1091]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[67]));
   ao22s01 U267858 (.o(n248532),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1603]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[579]));
   ao22s01 U267859 (.o(n248531),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1347]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[323]));
   ao22s01 U267860 (.o(n248530),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1859]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[835]));
   ao22s01 U267861 (.o(n248537),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1155]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[131]));
   ao22s01 U267862 (.o(n248536),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1667]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[643]));
   ao22s01 U267863 (.o(n248535),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1411]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[387]));
   ao22s01 U267864 (.o(n248534),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1923]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[899]));
   ao22s01 U267865 (.o(n248541),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1219]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[195]));
   ao22s01 U267866 (.o(n248540),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1731]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[707]));
   ao22s01 U267867 (.o(n248539),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1475]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[451]));
   ao22s01 U267868 (.o(n248538),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1987]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[963]));
   ao22s01 U267869 (.o(n248545),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1027]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[3]));
   ao22f01 U267870 (.o(n248544),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1539]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[515]));
   ao22s01 U267871 (.o(n248543),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1283]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[259]));
   ao22s01 U267872 (.o(n248542),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1795]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[771]));
   na02s01 U267873 (.o(regtop_w1_hdi00_q[3]),
	.a(n248551),
	.b(n248550));
   ao22s01 U267874 (.o(n248555),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1124]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[100]));
   ao22s01 U267875 (.o(n248553),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1380]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[356]));
   ao22s01 U267876 (.o(n248552),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1892]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[868]));
   ao22f01 U267877 (.o(n248559),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1188]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[164]));
   ao22s01 U267878 (.o(n248558),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1700]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[676]));
   ao22s01 U267879 (.o(n248557),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1444]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[420]));
   ao22s01 U267880 (.o(n248556),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1956]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[932]));
   ao22s01 U267881 (.o(n248563),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1252]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[228]));
   ao22s01 U267882 (.o(n248562),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1764]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[740]));
   ao22s01 U267883 (.o(n248561),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1508]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[484]));
   ao22s01 U267884 (.o(n248560),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2020]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[996]));
   ao22s01 U267885 (.o(n248567),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1060]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[36]));
   ao22s01 U267886 (.o(n248566),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1572]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[548]));
   ao22s01 U267887 (.o(n248565),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1316]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[292]));
   ao22s01 U267888 (.o(n248564),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1828]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[804]));
   ao22s01 U267889 (.o(n248574),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1604]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[580]));
   ao22s01 U267890 (.o(n248573),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1348]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[324]));
   ao22s01 U267891 (.o(n248572),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1860]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[836]));
   ao22s01 U267892 (.o(n248579),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1156]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[132]));
   ao22s01 U267893 (.o(n248578),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1668]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[644]));
   ao22s01 U267894 (.o(n248577),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1412]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[388]));
   ao22s01 U267895 (.o(n248576),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1924]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[900]));
   ao22s01 U267896 (.o(n248583),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1220]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[196]));
   ao22s01 U267897 (.o(n248582),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1732]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[708]));
   ao22s01 U267898 (.o(n248581),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1476]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[452]));
   ao22s01 U267899 (.o(n248580),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1988]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[964]));
   ao22s01 U267900 (.o(n248587),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1028]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[4]));
   ao22s01 U267901 (.o(n248586),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1540]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[516]));
   ao22s01 U267902 (.o(n248585),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1284]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[260]));
   na02s01 U267903 (.o(regtop_w1_hdi00_q[4]),
	.a(n248593),
	.b(n248592));
   ao22s01 U267904 (.o(n248597),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1121]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[97]));
   ao22s01 U267905 (.o(n248596),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1633]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[609]));
   ao22s01 U267906 (.o(n248595),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1377]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[353]));
   ao22s01 U267907 (.o(n248594),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1889]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[865]));
   ao22s01 U267908 (.o(n248601),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1185]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[161]));
   ao22s01 U267909 (.o(n248600),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1697]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[673]));
   ao22s01 U267910 (.o(n248599),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1441]),
	.c(FE_OFN54_n247067),
	.d(regtop_dchdi_w1_hdi00[417]));
   ao22s01 U267911 (.o(n248605),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1249]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[225]));
   ao22s01 U267912 (.o(n248604),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1761]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[737]));
   ao22s01 U267913 (.o(n248603),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1505]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[481]));
   ao22s01 U267914 (.o(n248602),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2017]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[993]));
   ao22s01 U267915 (.o(n248609),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1057]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[33]));
   ao22s01 U267916 (.o(n248608),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1569]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[545]));
   ao22s01 U267917 (.o(n248607),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1313]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[289]));
   ao22s01 U267918 (.o(n248606),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1825]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[801]));
   ao22s01 U267919 (.o(n248617),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1089]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[65]));
   ao22s01 U267920 (.o(n248616),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1601]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[577]));
   ao22s01 U267921 (.o(n248615),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1345]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[321]));
   ao22s01 U267922 (.o(n248614),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1857]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[833]));
   ao22s01 U267923 (.o(n248621),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1153]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[129]));
   ao22s01 U267924 (.o(n248620),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1665]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[641]));
   ao22s01 U267925 (.o(n248619),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1409]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[385]));
   ao22s01 U267926 (.o(n248618),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1921]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[897]));
   ao22s01 U267927 (.o(n248625),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1217]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[193]));
   ao22s01 U267928 (.o(n248624),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1729]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[705]));
   ao22s01 U267929 (.o(n248623),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1473]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[449]));
   ao22s01 U267930 (.o(n248622),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1985]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[961]));
   ao22s01 U267931 (.o(n248629),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1025]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[1]));
   ao22f02 U267932 (.o(n248628),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1537]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[513]));
   ao22s01 U267933 (.o(n248627),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1281]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[257]));
   ao22s01 U267934 (.o(n248626),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1793]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[769]));
   na02s01 U267935 (.o(regtop_w1_hdi00_q[1]),
	.a(n248635),
	.b(FE_OFN512_n248634));
   ao22s01 U267936 (.o(n248639),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1125]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[101]));
   ao22s01 U267937 (.o(n248638),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1637]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[613]));
   ao22s01 U267938 (.o(n248637),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1381]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[357]));
   ao22s01 U267939 (.o(n248636),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1893]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[869]));
   ao22s01 U267940 (.o(n248643),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1189]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[165]));
   ao22s01 U267941 (.o(n248642),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1701]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[677]));
   ao22s01 U267942 (.o(n248641),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1445]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[421]));
   ao22s01 U267943 (.o(n248640),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1957]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[933]));
   ao22s01 U267944 (.o(n248647),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1253]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[229]));
   ao22s01 U267945 (.o(n248646),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1765]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[741]));
   ao22s01 U267946 (.o(n248645),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1509]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[485]));
   ao22s01 U267947 (.o(n248644),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2021]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[997]));
   ao22s01 U267948 (.o(n248651),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1061]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[37]));
   ao22s01 U267949 (.o(n248650),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1573]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[549]));
   ao22s01 U267950 (.o(n248648),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1829]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[805]));
   ao22s01 U267951 (.o(n248659),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1093]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[69]));
   ao22f02 U267952 (.o(n248658),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1605]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[581]));
   ao22s01 U267953 (.o(n248657),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1349]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[325]));
   ao22s01 U267954 (.o(n248656),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1861]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[837]));
   ao22s01 U267955 (.o(n248663),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1157]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[133]));
   ao22s01 U267956 (.o(n248662),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1669]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[645]));
   ao22s01 U267957 (.o(n248661),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1413]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[389]));
   ao22s01 U267958 (.o(n248660),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1925]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[901]));
   ao22s01 U267959 (.o(n248667),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1221]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[197]));
   ao22s01 U267960 (.o(n248666),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1733]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[709]));
   ao22s01 U267961 (.o(n248665),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1477]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[453]));
   ao22s01 U267962 (.o(n248664),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1989]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[965]));
   ao22s01 U267963 (.o(n248671),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1029]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[5]));
   ao22s01 U267964 (.o(n248669),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1285]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[261]));
   ao22s01 U267965 (.o(n248668),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1797]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[773]));
   ao22s01 U267966 (.o(n248681),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1129]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[105]));
   ao22s01 U267967 (.o(n248680),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1641]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[617]));
   ao22s01 U267968 (.o(n248679),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1385]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[361]));
   ao22s01 U267969 (.o(n248678),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1897]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[873]));
   ao22s01 U267970 (.o(n248685),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1193]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[169]));
   ao22s01 U267971 (.o(n248684),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1705]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[681]));
   ao22s01 U267972 (.o(n248683),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1449]),
	.c(FE_OFN54_n247067),
	.d(regtop_dchdi_w1_hdi00[425]));
   ao22s01 U267973 (.o(n248682),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1961]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[937]));
   ao22s01 U267974 (.o(n248689),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1257]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[233]));
   ao22s01 U267975 (.o(n248688),
	.a(FE_OFN146_n248372),
	.b(regtop_dchdi_w1_hdi00[1769]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[745]));
   ao22s01 U267976 (.o(n248687),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1513]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[489]));
   ao22s01 U267977 (.o(n248686),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2025]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1001]));
   ao22s01 U267978 (.o(n248693),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1065]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[41]));
   ao22s01 U267979 (.o(n248692),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1577]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[553]));
   ao22s01 U267980 (.o(n248691),
	.a(n248139),
	.b(regtop_dchdi_w1_hdi00[1321]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[297]));
   ao22s01 U267981 (.o(n248690),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1833]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[809]));
   ao22s01 U267982 (.o(n248701),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1097]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[73]));
   ao22f01 U267983 (.o(n248700),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1609]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[585]));
   ao22s01 U267984 (.o(n248699),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1353]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[329]));
   ao22s01 U267985 (.o(n248698),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1865]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[841]));
   ao22s01 U267986 (.o(n248705),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1161]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[137]));
   ao22s01 U267987 (.o(n248703),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1417]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[393]));
   ao22s01 U267988 (.o(n248702),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1929]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[905]));
   ao22s01 U267989 (.o(n248709),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1225]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[201]));
   ao22s01 U267990 (.o(n248708),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1737]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[713]));
   ao22s01 U267991 (.o(n248707),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1481]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[457]));
   ao22f01 U267992 (.o(n248706),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1993]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[969]));
   ao22s01 U267993 (.o(n248713),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1033]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[9]));
   ao22s01 U267994 (.o(n248712),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1545]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[521]));
   ao22s01 U267995 (.o(n248711),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1289]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[265]));
   ao22s01 U267996 (.o(n248710),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1801]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[777]));
   na02f03 U267997 (.o(regtop_w1_hdi00_q[9]),
	.a(n248719),
	.b(n248718));
   ao22s01 U267998 (.o(n248723),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1128]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[104]));
   ao22s01 U267999 (.o(n248722),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1640]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[616]));
   ao22s01 U268000 (.o(n248721),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1384]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[360]));
   ao22s01 U268001 (.o(n248720),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1896]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[872]));
   ao22f01 U268002 (.o(n248727),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1192]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[168]));
   ao22s01 U268003 (.o(n248726),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1704]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[680]));
   ao22s01 U268004 (.o(n248725),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1448]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[424]));
   ao22s01 U268005 (.o(n248724),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1960]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[936]));
   ao22s01 U268006 (.o(n248730),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1768]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[744]));
   ao22s01 U268007 (.o(n248729),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1512]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[488]));
   ao22f01 U268008 (.o(n248728),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2024]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1000]));
   ao22s01 U268009 (.o(n248735),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1064]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[40]));
   ao22s01 U268010 (.o(n248734),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1576]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[552]));
   ao22s01 U268011 (.o(n248733),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1320]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[296]));
   ao22s01 U268012 (.o(n248732),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1832]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[808]));
   ao22s01 U268013 (.o(n248743),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1096]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[72]));
   ao22s01 U268014 (.o(n248742),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1608]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[584]));
   ao22s01 U268015 (.o(n248741),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1352]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[328]));
   ao22s01 U268016 (.o(n248740),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1864]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[840]));
   ao22s01 U268017 (.o(n248747),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1160]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[136]));
   ao22s01 U268018 (.o(n248746),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1672]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[648]));
   ao22s01 U268019 (.o(n248745),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1416]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[392]));
   ao22s01 U268020 (.o(n248751),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1224]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[200]));
   ao22s01 U268021 (.o(n248750),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1736]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[712]));
   ao22s01 U268022 (.o(n248749),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1480]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[456]));
   ao22s01 U268023 (.o(n248748),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[1992]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[968]));
   ao22s01 U268024 (.o(n248755),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1032]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[8]));
   ao22s01 U268025 (.o(n248754),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1544]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[520]));
   ao22s01 U268026 (.o(n248753),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1288]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[264]));
   ao22s01 U268027 (.o(n248752),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1800]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[776]));
   na02s01 U268028 (.o(regtop_w1_hdi00_q[8]),
	.a(n248761),
	.b(FE_OFN386_n248760));
   ao22s01 U268029 (.o(n248765),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1126]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[102]));
   ao22s01 U268030 (.o(n248764),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1638]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[614]));
   ao22s01 U268031 (.o(n248763),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1382]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[358]));
   ao22s01 U268032 (.o(n248762),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1894]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[870]));
   ao22s01 U268033 (.o(n248769),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1190]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[166]));
   ao22s01 U268034 (.o(n248768),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1702]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[678]));
   ao22s01 U268035 (.o(n248767),
	.a(FE_OFN81_n248127),
	.b(regtop_dchdi_w1_hdi00[1446]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[422]));
   ao22s01 U268036 (.o(n248766),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1958]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[934]));
   ao22s01 U268037 (.o(n248773),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1254]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[230]));
   ao22s01 U268038 (.o(n248772),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1766]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[742]));
   ao22s01 U268039 (.o(n248771),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1510]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[486]));
   ao22f01 U268040 (.o(n248770),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2022]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[998]));
   ao22s01 U268041 (.o(n248776),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1574]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[550]));
   ao22s01 U268042 (.o(n248775),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1318]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[294]));
   ao22s01 U268043 (.o(n248774),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1830]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[806]));
   ao22s01 U268044 (.o(n248785),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1094]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[70]));
   ao22s01 U268045 (.o(n248784),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1606]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[582]));
   ao22s01 U268046 (.o(n248783),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1350]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[326]));
   ao22s01 U268047 (.o(n248782),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1862]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[838]));
   ao22s01 U268048 (.o(n248789),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1158]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[134]));
   ao22f02 U268049 (.o(n248788),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1670]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[646]));
   ao22s01 U268050 (.o(n248787),
	.a(FE_OFN108_n248160),
	.b(regtop_dchdi_w1_hdi00[1414]),
	.c(n247099),
	.d(regtop_dchdi_w1_hdi00[390]));
   ao22s01 U268051 (.o(n248786),
	.a(FE_OFN113_n248162),
	.b(regtop_dchdi_w1_hdi00[1926]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[902]));
   ao22s01 U268052 (.o(n248793),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1222]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[198]));
   ao22s01 U268053 (.o(n248792),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1734]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[710]));
   ao22s01 U268054 (.o(n248791),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1478]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[454]));
   ao22s01 U268055 (.o(n248797),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1030]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[6]));
   ao22s01 U268056 (.o(n248796),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1542]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[518]));
   ao22s01 U268057 (.o(n248795),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1286]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[262]));
   ao22s01 U268058 (.o(n248794),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1798]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[774]));
   na02f03 U268059 (.o(regtop_w1_hdi00_q[6]),
	.a(n248803),
	.b(n248802));
   ao22s01 U268060 (.o(n248807),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1151]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[127]));
   ao22s01 U268061 (.o(n248806),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1663]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[639]));
   ao22s01 U268062 (.o(n248805),
	.a(FE_OFN72_n248119),
	.b(regtop_dchdi_w1_hdi00[1407]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[383]));
   ao22s01 U268063 (.o(n248804),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1919]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[895]));
   ao22s01 U268064 (.o(n248811),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1215]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[191]));
   ao22s01 U268065 (.o(n248810),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1727]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[703]));
   ao22s01 U268066 (.o(n248809),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1471]),
	.c(FE_OFN54_n247067),
	.d(regtop_dchdi_w1_hdi00[447]));
   ao22s01 U268067 (.o(n248808),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1983]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[959]));
   ao22s01 U268068 (.o(n248815),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1279]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[255]));
   ao22s01 U268069 (.o(n248814),
	.a(FE_OFN146_n248372),
	.b(regtop_dchdi_w1_hdi00[1791]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[767]));
   ao22s01 U268070 (.o(n248813),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1535]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[511]));
   ao22s01 U268071 (.o(n248812),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2047]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1023]));
   ao22s01 U268072 (.o(n248819),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1087]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[63]));
   ao22s01 U268073 (.o(n248818),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1599]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[575]));
   ao22s01 U268074 (.o(n248817),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1343]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[319]));
   ao22s01 U268075 (.o(n248816),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1855]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[831]));
   ao22s01 U268076 (.o(n248827),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1119]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[95]));
   ao22s01 U268077 (.o(n248826),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1631]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[607]));
   ao22s01 U268078 (.o(n248825),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1375]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[351]));
   ao22s01 U268079 (.o(n248824),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1887]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[863]));
   ao22s01 U268080 (.o(n248831),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1183]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[159]));
   ao22s01 U268081 (.o(n248830),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1695]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[671]));
   ao22s01 U268082 (.o(n248829),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1439]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[415]));
   ao22s01 U268083 (.o(n248828),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1951]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[927]));
   ao22s01 U268084 (.o(n248835),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1247]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[223]));
   ao22s01 U268085 (.o(n248834),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1759]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[735]));
   ao22s01 U268086 (.o(n248833),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1503]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[479]));
   ao22s01 U268087 (.o(n248832),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2015]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[991]));
   ao22f02 U268088 (.o(n248839),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1055]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[31]));
   ao22s01 U268089 (.o(n248838),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1567]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[543]));
   ao22s01 U268090 (.o(n248837),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1311]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[287]));
   ao22s01 U268091 (.o(n248836),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1823]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[799]));
   ao22s01 U268092 (.o(n248857),
	.a(FE_OFN70_n248118),
	.b(regtop_dchdi_w1_hdi00[1141]),
	.c(FE_OFN128_n248355),
	.d(regtop_dchdi_w1_hdi00[117]));
   ao22s01 U268093 (.o(n248856),
	.a(FE_OFN132_n248357),
	.b(regtop_dchdi_w1_hdi00[1653]),
	.c(FE_OFN130_n248356),
	.d(regtop_dchdi_w1_hdi00[629]));
   ao22s01 U268094 (.o(n248855),
	.a(FE_OFN73_n248119),
	.b(regtop_dchdi_w1_hdi00[1397]),
	.c(FE_OFN51_n247057),
	.d(regtop_dchdi_w1_hdi00[373]));
   ao22s01 U268095 (.o(n248854),
	.a(FE_OFN77_n248121),
	.b(regtop_dchdi_w1_hdi00[1909]),
	.c(FE_OFN75_n248120),
	.d(regtop_dchdi_w1_hdi00[885]));
   ao22s01 U268096 (.o(n248869),
	.a(FE_OFN79_n248126),
	.b(regtop_dchdi_w1_hdi00[1205]),
	.c(FE_OFN134_n248362),
	.d(regtop_dchdi_w1_hdi00[181]));
   ao22s01 U268097 (.o(n248868),
	.a(FE_OFN138_n248364),
	.b(regtop_dchdi_w1_hdi00[1717]),
	.c(FE_OFN136_n248363),
	.d(regtop_dchdi_w1_hdi00[693]));
   ao22s01 U268098 (.o(n248867),
	.a(FE_OFN82_n248127),
	.b(regtop_dchdi_w1_hdi00[1461]),
	.c(FE_OFN53_n247067),
	.d(regtop_dchdi_w1_hdi00[437]));
   ao22s01 U268099 (.o(n248866),
	.a(FE_OFN86_n248129),
	.b(regtop_dchdi_w1_hdi00[1973]),
	.c(FE_OFN84_n248128),
	.d(regtop_dchdi_w1_hdi00[949]));
   ao22s01 U268100 (.o(n248881),
	.a(FE_OFN142_n248370),
	.b(regtop_dchdi_w1_hdi00[1269]),
	.c(FE_OFN140_n248369),
	.d(regtop_dchdi_w1_hdi00[245]));
   ao22s01 U268101 (.o(n248880),
	.a(FE_OFN147_n248372),
	.b(regtop_dchdi_w1_hdi00[1781]),
	.c(FE_OFN144_n248371),
	.d(regtop_dchdi_w1_hdi00[757]));
   ao22s01 U268102 (.o(n248879),
	.a(FE_OFN149_n248373),
	.b(regtop_dchdi_w1_hdi00[1525]),
	.c(FE_OFN56_n247074),
	.d(regtop_dchdi_w1_hdi00[501]));
   ao22f01 U268103 (.o(n248878),
	.a(FE_OFN153_n248375),
	.b(regtop_dchdi_w1_hdi00[2037]),
	.c(FE_OFN151_n248374),
	.d(regtop_dchdi_w1_hdi00[1013]));
   ao22f01 U268104 (.o(n248893),
	.a(FE_OFN88_n248138),
	.b(regtop_dchdi_w1_hdi00[1077]),
	.c(FE_OFN155_n248380),
	.d(regtop_dchdi_w1_hdi00[53]));
   ao22s01 U268105 (.o(n248892),
	.a(FE_OFN159_n248382),
	.b(regtop_dchdi_w1_hdi00[1589]),
	.c(FE_OFN157_n248381),
	.d(regtop_dchdi_w1_hdi00[565]));
   ao22s01 U268106 (.o(n248891),
	.a(FE_OFN90_n248139),
	.b(regtop_dchdi_w1_hdi00[1333]),
	.c(FE_OFN64_n247509),
	.d(regtop_dchdi_w1_hdi00[309]));
   ao22f02 U268107 (.o(n248890),
	.a(FE_OFN94_n248141),
	.b(regtop_dchdi_w1_hdi00[1845]),
	.c(n248140),
	.d(regtop_dchdi_w1_hdi00[821]));
   ao22s01 U268108 (.o(n248909),
	.a(FE_OFN96_n248150),
	.b(regtop_dchdi_w1_hdi00[1109]),
	.c(FE_OFN161_n248391),
	.d(regtop_dchdi_w1_hdi00[85]));
   ao22f02 U268109 (.o(n248908),
	.a(FE_OFN165_n248393),
	.b(regtop_dchdi_w1_hdi00[1621]),
	.c(FE_OFN163_n248392),
	.d(regtop_dchdi_w1_hdi00[597]));
   ao22s01 U268110 (.o(n248907),
	.a(FE_OFN98_n248151),
	.b(regtop_dchdi_w1_hdi00[1365]),
	.c(FE_OFN58_n247092),
	.d(regtop_dchdi_w1_hdi00[341]));
   ao22s01 U268111 (.o(n248906),
	.a(FE_OFN102_n248153),
	.b(regtop_dchdi_w1_hdi00[1877]),
	.c(FE_OFN100_n248152),
	.d(regtop_dchdi_w1_hdi00[853]));
   ao22s01 U268112 (.o(n248921),
	.a(FE_OFN106_n248159),
	.b(regtop_dchdi_w1_hdi00[1173]),
	.c(FE_OFN104_n248158),
	.d(regtop_dchdi_w1_hdi00[149]));
   ao22s01 U268113 (.o(n248920),
	.a(FE_OFN169_n248399),
	.b(regtop_dchdi_w1_hdi00[1685]),
	.c(FE_OFN167_n248398),
	.d(regtop_dchdi_w1_hdi00[661]));
   ao22s01 U268114 (.o(n248919),
	.a(FE_OFN109_n248160),
	.b(regtop_dchdi_w1_hdi00[1429]),
	.c(FE_OFN60_n247099),
	.d(regtop_dchdi_w1_hdi00[405]));
   ao22s01 U268115 (.o(n248918),
	.a(FE_OFN114_n248162),
	.b(regtop_dchdi_w1_hdi00[1941]),
	.c(n248161),
	.d(regtop_dchdi_w1_hdi00[917]));
   ao22s01 U268116 (.o(n248933),
	.a(FE_OFN173_n248405),
	.b(regtop_dchdi_w1_hdi00[1237]),
	.c(FE_OFN171_n248404),
	.d(regtop_dchdi_w1_hdi00[213]));
   ao22s01 U268117 (.o(n248932),
	.a(FE_OFN177_n248407),
	.b(regtop_dchdi_w1_hdi00[1749]),
	.c(FE_OFN175_n248406),
	.d(regtop_dchdi_w1_hdi00[725]));
   ao22s01 U268118 (.o(n248931),
	.a(FE_OFN179_n248408),
	.b(regtop_dchdi_w1_hdi00[1493]),
	.c(FE_OFN62_n247107),
	.d(regtop_dchdi_w1_hdi00[469]));
   ao22s01 U268119 (.o(n248930),
	.a(n248168),
	.b(regtop_dchdi_w1_hdi00[2005]),
	.c(FE_OFN116_n248167),
	.d(regtop_dchdi_w1_hdi00[981]));
   ao22s01 U268120 (.o(n248945),
	.a(FE_OFN120_n248173),
	.b(regtop_dchdi_w1_hdi00[1045]),
	.c(FE_OFN181_n248413),
	.d(regtop_dchdi_w1_hdi00[21]));
   ao22s01 U268121 (.o(n248944),
	.a(FE_OFN185_n248415),
	.b(regtop_dchdi_w1_hdi00[1557]),
	.c(FE_OFN183_n248414),
	.d(regtop_dchdi_w1_hdi00[533]));
   ao22s01 U268122 (.o(n248943),
	.a(FE_OFN122_n248174),
	.b(regtop_dchdi_w1_hdi00[1301]),
	.c(FE_OFN66_n247531),
	.d(regtop_dchdi_w1_hdi00[277]));
   ao22s01 U268123 (.o(n248942),
	.a(FE_OFN126_n248176),
	.b(regtop_dchdi_w1_hdi00[1813]),
	.c(FE_OFN124_n248175),
	.d(regtop_dchdi_w1_hdi00[789]));
   na02s01 U268124 (.o(regtop_w1_hdi00_q[21]),
	.a(n248951),
	.b(n248950));
   ao22s01 U268125 (.o(n248958),
	.a(n248978),
	.b(regtop_g_usrd_r[27]),
	.c(n248977),
	.d(regtop_g_atscd_r[27]));
   in01s01 U268126 (.o(n248955),
	.a(n248952));
   in01s01 U268127 (.o(n248954),
	.a(n248953));
   ao22s01 U268128 (.o(n248961),
	.a(n248978),
	.b(regtop_g_usrd_r[31]),
	.c(n248977),
	.d(regtop_g_atscd_r[31]));
   ao22s01 U268129 (.o(n248964),
	.a(n248978),
	.b(regtop_g_usrd_r[24]),
	.c(n248977),
	.d(regtop_g_atscd_r[24]));
   ao22s01 U268130 (.o(n248967),
	.a(n248978),
	.b(regtop_g_usrd_r[28]),
	.c(n248977),
	.d(regtop_g_atscd_r[28]));
   ao22s01 U268131 (.o(n248970),
	.a(n248978),
	.b(regtop_g_usrd_r[29]),
	.c(n248977),
	.d(regtop_g_atscd_r[29]));
   ao22s01 U268132 (.o(n248973),
	.a(n248978),
	.b(regtop_g_usrd_r[30]),
	.c(n248977),
	.d(regtop_g_atscd_r[30]));
   ao22f01 U268133 (.o(n248976),
	.a(n248978),
	.b(regtop_g_usrd_r[26]),
	.c(n248977),
	.d(regtop_g_atscd_r[26]));
   ao22s01 U268134 (.o(n248983),
	.a(n248978),
	.b(regtop_g_usrd_r[25]),
	.c(n248977),
	.d(regtop_g_atscd_r[25]));
   na02s01 U268136 (.o(n248986),
	.a(n249113),
	.b(n252731));
   na02s01 U268137 (.o(n248987),
	.a(n249242),
	.b(n248986));
   in01s01 U268138 (.o(n244986),
	.a(n248989));
   in01f02 U268140 (.o(n249106),
	.a(n248996));
   na02s01 U268141 (.o(n249000),
	.a(n246670),
	.b(n248999));
   in01s01 U268142 (.o(n249010),
	.a(n249000));
   in01s01 U268143 (.o(n249002),
	.a(vldtop_vld_syndec_UREG[7]));
   in01s01 U268144 (.o(n249009),
	.a(n249008));
   no02s01 U268145 (.o(n249017),
	.a(n249016),
	.b(n249015));
   na02s01 U268146 (.o(n249024),
	.a(n246964),
	.b(n249023));
   in01s01 U268147 (.o(n249025),
	.a(n249024));
   ao22f02 U268148 (.o(n249030),
	.a(n249066),
	.b(n249029),
	.c(regtop_g_adb_r[4]),
	.d(n249041));
   in01f02 U268149 (.o(n249038),
	.a(n249030));
   no02f01 U268150 (.o(n249033),
	.a(n249031),
	.b(n249038));
   na02f03 U268151 (.o(n249052),
	.a(n249031),
	.b(n249038));
   no02f01 U268152 (.o(n249034),
	.a(n249033),
	.b(n249032));
   ao22f04 U268153 (.o(n249037),
	.a(n249036),
	.b(n249066),
	.c(regtop_g_adb_r[5]),
	.d(n249041));
   in01f02 U268154 (.o(n249051),
	.a(n249037));
   no02f04 U268155 (.o(n249045),
	.a(n249040),
	.b(n249039));
   in01f01 U268156 (.o(n249043),
	.a(n249044));
   no02f01 U268157 (.o(n249047),
	.a(n249045),
	.b(n249043));
   na02f04 U268158 (.o(n249067),
	.a(n249045),
	.b(n249043));
   in01f01 U268159 (.o(n249046),
	.a(n249067));
   na02f02 U268160 (.o(n249053),
	.a(n249052),
	.b(n249037));
   ao12f02 U268161 (.o(n249058),
	.a(n249072),
	.b(n249057),
	.c(n249073));
   no02s01 U268162 (.o(n249062),
	.a(n249061),
	.b(n249060));
   ao22f01 U268163 (.o(n249065),
	.a(n249064),
	.b(vldtop_vld_syndec_vld_vscdet_v_search_1st_r),
	.c(n249063),
	.d(n249062));
   in01s01 U268164 (.o(n212488),
	.a(n249065));
   in01s01 U268165 (.o(n249069),
	.a(n249066));
   na02f04 U268166 (.o(n249068),
	.a(n249067),
	.b(n249069));
   na02f01 U268167 (.o(n249071),
	.a(n249067),
	.b(n249068));
   na02f02 U268168 (.o(n249070),
	.a(n249069),
	.b(n249068));
   na02f02 U268169 (.o(n249074),
	.a(n249071),
	.b(n249070));
   in01s01 U268170 (.o(n249080),
	.a(n252597));
   na02m01 U268171 (.o(n249086),
	.a(regtop_g_paramdata_r[24]),
	.b(n249132));
   na02s01 U268172 (.o(n249090),
	.a(n249128),
	.b(regtop_g_usrd_r[19]));
   na02s01 U268173 (.o(n249096),
	.a(n249128),
	.b(regtop_g_usrd_r[17]));
   na02s01 U268174 (.o(n249098),
	.a(n249097),
	.b(n249096));
   na02s01 U268175 (.o(n249101),
	.a(n249128),
	.b(regtop_g_usrd_r[20]));
   na02s01 U268176 (.o(n249103),
	.a(n249102),
	.b(n249101));
   oa22f01 U268177 (.o(n249112),
	.a(n249107),
	.b(n252664),
	.c(n249106),
	.d(n252660));
   in01s01 U268178 (.o(n249111),
	.a(n249108));
   na02s01 U268179 (.o(n249110),
	.a(n252684),
	.b(n249109));
   in01s01 U268180 (.o(n249115),
	.a(n249114));
   na02s01 U268181 (.o(n249116),
	.a(n249128),
	.b(regtop_g_usrd_r[16]));
   na02s01 U268182 (.o(n249121),
	.a(n249128),
	.b(regtop_g_usrd_r[21]));
   na02f01 U268183 (.o(n249123),
	.a(n249122),
	.b(n249121));
   na02s01 U268184 (.o(n249129),
	.a(n249128),
	.b(regtop_g_usrd_r[18]));
   in01s01 U268185 (.o(n249136),
	.a(n249135));
   na02s01 U268186 (.o(n252782),
	.a(regtop_g_paramdata_r[18]),
	.b(n249241));
   no02s01 U268187 (.o(n249144),
	.a(n252658),
	.b(n249247));
   na02s01 U268189 (.o(n249141),
	.a(FE_OFN551_n249140),
	.b(regtop_g_atscd_r[9]));
   in01f01 U268190 (.o(n252646),
	.a(regtop_g_paramdata_r[12]));
   ao22s01 U268191 (.o(n249149),
	.a(n249211),
	.b(regtop_g_paramdata_r[10]),
	.c(regtop_g_paramdata_r[23]),
	.d(n249210));
   oa12s01 U268192 (.o(n249150),
	.a(n249149),
	.b(FE_OFN573_n249242),
	.c(n252646));
   in01f01 U268193 (.o(n252644),
	.a(regtop_g_paramdata_r[11]));
   ao22s01 U268194 (.o(n249154),
	.a(n249211),
	.b(regtop_g_paramdata_r[9]),
	.c(regtop_g_paramdata_r[22]),
	.d(n249210));
   oa12s01 U268195 (.o(n249155),
	.a(n249154),
	.b(FE_OFN573_n249242),
	.c(n252644));
   ao22s01 U268196 (.o(n249159),
	.a(n249211),
	.b(regtop_g_paramdata_r[8]),
	.c(regtop_g_paramdata_r[21]),
	.d(n249210));
   oa12s01 U268197 (.o(n249160),
	.a(n249159),
	.b(FE_OFN573_n249242),
	.c(n252670));
   ao22s01 U268198 (.o(n249164),
	.a(n249211),
	.b(regtop_g_paramdata_r[7]),
	.c(regtop_g_paramdata_r[20]),
	.d(n249210));
   oa12s01 U268199 (.o(n249166),
	.a(n249164),
	.b(FE_OFN573_n249242),
	.c(n249165));
   in01s01 U268200 (.o(n249171),
	.a(regtop_g_paramdata_r[8]));
   ao22s01 U268201 (.o(n249170),
	.a(n249211),
	.b(regtop_g_paramdata_r[6]),
	.c(regtop_g_paramdata_r[19]),
	.d(n249210));
   oa12s01 U268202 (.o(n249172),
	.a(n249170),
	.b(FE_OFN573_n249242),
	.c(n249171));
   in01s01 U268203 (.o(n249177),
	.a(regtop_g_paramdata_r[7]));
   ao22s01 U268204 (.o(n249176),
	.a(n249211),
	.b(regtop_g_paramdata_r[5]),
	.c(regtop_g_paramdata_r[18]),
	.d(n249210));
   oa12f01 U268205 (.o(n249178),
	.a(n249176),
	.b(n249242),
	.c(n249177));
   no02f01 U268206 (.o(n249186),
	.a(n249189),
	.b(n252658));
   in01s01 U268207 (.o(n249184),
	.a(regtop_g_paramdata_r[6]));
   ao22s01 U268208 (.o(n249183),
	.a(n249211),
	.b(regtop_g_paramdata_r[4]),
	.c(regtop_g_paramdata_r[17]),
	.d(n249210));
   oa12s01 U268209 (.o(n249185),
	.a(n249183),
	.b(FE_OFN573_n249242),
	.c(n249184));
   in01s01 U268210 (.o(n249191),
	.a(regtop_g_paramdata_r[5]));
   ao22s01 U268211 (.o(n249190),
	.a(n249211),
	.b(regtop_g_paramdata_r[3]),
	.c(n249210),
	.d(regtop_g_paramdata_r[16]));
   oa12s01 U268212 (.o(n249192),
	.a(n249190),
	.b(n249242),
	.c(n249191));
   na02s01 U268213 (.o(n252798),
	.a(regtop_g_paramdata_r[22]),
	.b(n249241));
   in01f02 U268214 (.o(n252654),
	.a(regtop_g_paramdata_r[16]));
   oa22f01 U268215 (.o(n249196),
	.a(FE_OFN483_n249211),
	.b(n252654),
	.c(n249242),
	.d(n252658));
   ao12m01 U268216 (.o(n249197),
	.a(n249196),
	.b(FE_OFN551_n249140),
	.c(regtop_g_atscd_r[13]));
   oa12m01 U268217 (.o(n249198),
	.a(n249197),
	.b(n252666),
	.c(n249247));
   na02s01 U268218 (.o(n252806),
	.a(regtop_g_paramdata_r[24]),
	.b(n249241));
   na02s01 U268219 (.o(n252810),
	.a(regtop_g_paramdata_r[17]),
	.b(n249241));
   in01f02 U268220 (.o(n252648),
	.a(regtop_g_paramdata_r[13]));
   na02s01 U268221 (.o(n252802),
	.a(regtop_g_paramdata_r[23]),
	.b(n249241));
   na02s01 U268222 (.o(n252786),
	.a(regtop_g_paramdata_r[19]),
	.b(n249241));
   in01f02 U268223 (.o(n252652),
	.a(regtop_g_paramdata_r[15]));
   na02s01 U268224 (.o(n252790),
	.a(regtop_g_paramdata_r[20]),
	.b(n249241));
   in01f02 U268225 (.o(n252650),
	.a(regtop_g_paramdata_r[14]));
   na02s01 U268226 (.o(n252794),
	.a(regtop_g_paramdata_r[21]),
	.b(n249241));
   no02s01 U268227 (.o(n253037),
	.a(n249255),
	.b(FE_OFN68_n247591));
   no02s01 U268228 (.o(n249256),
	.a(busrtop_b_rreq_vrh_add1_r[6]),
	.b(busrtop_b_rreq_vrh_add1_r[7]));
   no02s01 U268229 (.o(n249260),
	.a(busrtop_b_rreq_vrh_add1_r[4]),
	.b(busrtop_b_rreq_vrh_add1_r[5]));
   na02s01 U268230 (.o(n249258),
	.a(n249256),
	.b(n249260));
   no02s01 U268231 (.o(n249257),
	.a(busrtop_b_rreq_vrh_add1_r[2]),
	.b(busrtop_b_rreq_vrh_add1_r[3]));
   no02s01 U268232 (.o(n249259),
	.a(n249258),
	.b(n249282));
   in01s01 U268233 (.o(n249272),
	.a(n249259));
   in01s01 U268234 (.o(n249263),
	.a(n249282));
   na02s01 U268235 (.o(n249276),
	.a(n249263),
	.b(n249260));
   no02s01 U268236 (.o(n249277),
	.a(n249276),
	.b(busrtop_b_rreq_vrh_add1_r[6]));
   in01s01 U268237 (.o(n249261),
	.a(n249277));
   na02s01 U268238 (.o(n249262),
	.a(busrtop_b_rreq_vrh_add1_r[7]),
	.b(n249261));
   na02s01 U268239 (.o(busrtop_b_rreq_N429),
	.a(n249272),
	.b(n249262));
   in01s01 U268240 (.o(n249888),
	.a(busrtop_b_rreq_vrh_add1_r[4]));
   na02s01 U268241 (.o(n249265),
	.a(n249263),
	.b(n249888));
   na02s01 U268242 (.o(n249264),
	.a(busrtop_b_rreq_vrh_add1_r[4]),
	.b(n249282));
   na02s01 U268243 (.o(busrtop_b_rreq_N426),
	.a(n249265),
	.b(n249264));
   in01s01 U268244 (.o(n249266),
	.a(n249276));
   no02s01 U268245 (.o(n249268),
	.a(n249265),
	.b(n249266));
   no02s01 U268246 (.o(n249267),
	.a(busrtop_b_rreq_vrh_add1_r[5]),
	.b(n249266));
   no02s01 U268247 (.o(busrtop_b_rreq_N427),
	.a(n249268),
	.b(n249267));
   na02s01 U268248 (.o(n249269),
	.a(n249273),
	.b(busrtop_b_rreq_vrh_add1_r[9]));
   na02s01 U268249 (.o(n249270),
	.a(busrtop_b_rreq_vrh_add1_r[9]),
	.b(n249269));
   na02s01 U268250 (.o(busrtop_b_rreq_N431),
	.a(n249271),
	.b(n249270));
   no02s01 U268251 (.o(n249275),
	.a(n249273),
	.b(n249272));
   no02s01 U268252 (.o(n249274),
	.a(busrtop_b_rreq_vrh_add1_r[8]),
	.b(n249273));
   no02s01 U268253 (.o(busrtop_b_rreq_N430),
	.a(n249275),
	.b(n249274));
   no02s01 U268254 (.o(n249279),
	.a(n249276),
	.b(n249277));
   no02s01 U268255 (.o(n249278),
	.a(busrtop_b_rreq_vrh_add1_r[6]),
	.b(n249277));
   in01s01 U268256 (.o(n249283),
	.a(n249287));
   no02s01 U268257 (.o(n249284),
	.a(n249283),
	.b(busrtop_b_rreq_vrh_add1_r[2]));
   in01s01 U268258 (.o(n249280),
	.a(n249284));
   na02s01 U268259 (.o(n249281),
	.a(busrtop_b_rreq_vrh_add1_r[3]),
	.b(n249280));
   na02s01 U268260 (.o(busrtop_b_rreq_N425),
	.a(n249282),
	.b(n249281));
   no02s01 U268261 (.o(n249286),
	.a(n249284),
	.b(n249283));
   no02s01 U268262 (.o(n249285),
	.a(busrtop_b_rreq_vrh_add1_r[2]),
	.b(n249284));
   no02s01 U268263 (.o(busrtop_b_rreq_N424),
	.a(n249286),
	.b(n249285));
   no02s01 U268264 (.o(n249289),
	.a(busrtop_b_rreq_vrh_add1_r[1]),
	.b(n249287));
   no02s01 U268265 (.o(busrtop_b_rreq_N423),
	.a(n249289),
	.b(n249288));
   in01s01 U268266 (.o(n253124),
	.a(n249290));
   in01s01 U268267 (.o(n253123),
	.a(n249291));
   in01s01 U268268 (.o(n253121),
	.a(n249293));
   in01s01 U268269 (.o(n253120),
	.a(n249294));
   in01s01 U268270 (.o(n253119),
	.a(n249295));
   in01s01 U268271 (.o(n253118),
	.a(n249296));
   in01s01 U268272 (.o(n253117),
	.a(n249297));
   in01s01 U268273 (.o(n253116),
	.a(n249298));
   in01s01 U268274 (.o(n253115),
	.a(n249299));
   in01s01 U268275 (.o(n253114),
	.a(n249300));
   in01s01 U268276 (.o(n253113),
	.a(n249301));
   in01s01 U268277 (.o(n253112),
	.a(n249302));
   in01s01 U268278 (.o(n253111),
	.a(n249303));
   in01s01 U268279 (.o(n253110),
	.a(n249304));
   in01s01 U268280 (.o(n253108),
	.a(n249306));
   in01s01 U268281 (.o(n253107),
	.a(n249307));
   in01s01 U268282 (.o(n253106),
	.a(n249308));
   in01s01 U268283 (.o(n253105),
	.a(n249309));
   in01s01 U268284 (.o(n253104),
	.a(n249310));
   in01s01 U268285 (.o(n253103),
	.a(n249311));
   in01s01 U268296 (.o(n249312),
	.a(cntrltop_ctmg_ctpedet_c_tmg_ferr_pre));
   no02s01 U268297 (.o(cntrltop_ctmg_ctpedet_N22),
	.a(cntrltop_ctmg_ctpedet_c_tmg_ferr_pre_d1_r),
	.b(n249312));
   no02s01 U268298 (.o(regtop_N1267),
	.a(n249925),
	.b(n252305));
   in01s01 U268299 (.o(n252308),
	.a(n249317));
   no02s01 U268300 (.o(regtop_N1279),
	.a(n252309),
	.b(n252308));
   in01s01 U268301 (.o(n249320),
	.a(busiftop_vmem_ch_r));
   no02s01 U268302 (.o(n249318),
	.a(n249320),
	.b(y1_bs_data_r[21]));
   ao22f03 U268303 (.o(n249321),
	.a(n249320),
	.b(busiftop_status_b_current_0_),
	.c(n249319),
	.d(n249318));
   in01s01 U268304 (.o(busiftop_N35),
	.a(n249321));
   in01s01 U268305 (.o(regtop_N1993),
	.a(n249322));
   na02s01 U268306 (.o(n249323),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[1]));
   in01s01 U268307 (.o(regtop_N1994),
	.a(n249323));
   na02s01 U268308 (.o(n249324),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[2]));
   in01s01 U268309 (.o(regtop_N1995),
	.a(n249324));
   na02s01 U268310 (.o(n249325),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[3]));
   in01s01 U268311 (.o(regtop_N1996),
	.a(n249325));
   na02f03 U268312 (.o(n249326),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[4]));
   na02s01 U268313 (.o(n249327),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[5]));
   in01s01 U268314 (.o(regtop_N1998),
	.a(n249327));
   na02s01 U268315 (.o(n249328),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[6]));
   in01s01 U268316 (.o(regtop_N1999),
	.a(n249328));
   na02s01 U268317 (.o(n249329),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[7]));
   in01s01 U268318 (.o(regtop_N2000),
	.a(n249329));
   na02s01 U268319 (.o(n249330),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[8]));
   in01s01 U268320 (.o(regtop_N2001),
	.a(n249330));
   na02f02 U268321 (.o(n249331),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[9]));
   in01s01 U268322 (.o(regtop_N2002),
	.a(n249331));
   na02s01 U268323 (.o(n249332),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[10]));
   in01s01 U268324 (.o(regtop_N2003),
	.a(n249332));
   na02f02 U268325 (.o(n249333),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[11]));
   in01s01 U268326 (.o(regtop_N2004),
	.a(n249333));
   na02s01 U268327 (.o(n249334),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[12]));
   in01s01 U268328 (.o(regtop_N2005),
	.a(n249334));
   na02s01 U268329 (.o(n249335),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[13]));
   in01s01 U268330 (.o(regtop_N2006),
	.a(n249335));
   na02s01 U268331 (.o(n249336),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[14]));
   in01s01 U268332 (.o(regtop_N2007),
	.a(n249336));
   in01s01 U268333 (.o(regtop_N2008),
	.a(n249337));
   na02s01 U268334 (.o(n249338),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[16]));
   in01s01 U268335 (.o(regtop_N2009),
	.a(n249338));
   na02s01 U268336 (.o(n249339),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[17]));
   in01s01 U268337 (.o(regtop_N2010),
	.a(n249339));
   na02f02 U268338 (.o(n249340),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[18]));
   in01s01 U268339 (.o(regtop_N2011),
	.a(n249340));
   na02f02 U268340 (.o(n249341),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[19]));
   na02f02 U268341 (.o(n249342),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[20]));
   in01f01 U268342 (.o(regtop_N2013),
	.a(n249342));
   na02f02 U268343 (.o(n249343),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[21]));
   in01s01 U268344 (.o(regtop_N2014),
	.a(n249343));
   na02f02 U268345 (.o(n249344),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[22]));
   in01s01 U268346 (.o(regtop_N2015),
	.a(n249344));
   na02s01 U268347 (.o(n249345),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[23]));
   in01s01 U268348 (.o(regtop_N2016),
	.a(n249345));
   na02f03 U268349 (.o(n249346),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[24]));
   in01s01 U268350 (.o(regtop_N2017),
	.a(n249346));
   na02s01 U268351 (.o(n249347),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[25]));
   in01s01 U268352 (.o(regtop_N2018),
	.a(n249347));
   na02s01 U268353 (.o(n249348),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[26]));
   in01s01 U268354 (.o(regtop_N2019),
	.a(n249348));
   na02s01 U268355 (.o(n249349),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[27]));
   in01s01 U268356 (.o(regtop_N2020),
	.a(n249349));
   na02s01 U268357 (.o(n249350),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[28]));
   in01s01 U268358 (.o(regtop_N2021),
	.a(n249350));
   na02f80 U268359 (.o(n249351),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[29]));
   in01s01 U268360 (.o(regtop_N2022),
	.a(n249351));
   in01s01 U268361 (.o(regtop_N2023),
	.a(n249352));
   na02s01 U268362 (.o(n249353),
	.a(regtop_g_rd_en2_r),
	.b(regtop_g_mem_rd_r[31]));
   in01s01 U268363 (.o(regtop_N2024),
	.a(n249353));
   in01s01 U268364 (.o(n249357),
	.a(n252873));
   oa12s01 U268365 (.o(n245111),
	.a(n252377),
	.b(regtop_g_init_cnt_r[0]),
	.c(n249357));
   oa12s01 U268366 (.o(n245110),
	.a(n252377),
	.b(n249355),
	.c(n249354));
   ao12s01 U268367 (.o(n249356),
	.a(n249355),
	.b(regtop_g_init_cnt_r[0]),
	.c(regtop_g_init_cnt_r[1]));
   oa12s01 U268368 (.o(n245109),
	.a(n252377),
	.b(n249357),
	.c(n249356));
   no04s01 U268369 (.o(n249358),
	.a(regtop_g_isfb_r),
	.b(regtop_g_isfp_r),
	.c(regtop_g_issr_r),
	.d(regtop_g_issw_r));
   in01s01 U268370 (.o(n249359),
	.a(n249358));
   no04f03 U268371 (.o(n245091),
	.a(regtop_g_isnf_r),
	.b(regtop_g_isdc_r),
	.c(regtop_g_isuc_r),
	.d(n249359));
   no03f06 U268372 (.o(n245090),
	.a(regtop_g_isph_r),
	.b(regtop_g_ispi_r),
	.c(regtop_g_issh_r));
   ao22s01 U268373 (.o(n249366),
	.a(n249813),
	.b(regtop_g_vf_r[2]),
	.c(FE_OFN400_n249836),
	.d(g_field_start_add_r[30]));
   ao22s01 U268374 (.o(n249365),
	.a(FE_OFN527_n249828),
	.b(regtop_g_fcho2_r[14]),
	.c(FE_OFN546_n245460),
	.d(regtop_g_ari_r[2]));
   ao22f01 U268375 (.o(n249364),
	.a(n249838),
	.b(regtop_g_fcho1_r[14]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcho0_r[14]));
   na02s01 U268376 (.o(n249361),
	.a(FE_OFN552_n245462),
	.b(regtop_g_pct_r[2]));
   ao12s01 U268377 (.o(n249360),
	.a(n249825),
	.b(n249786),
	.c(g_hsdc_r[6]));
   na02s01 U268378 (.o(n249362),
	.a(n249361),
	.b(n249360));
   ao12s01 U268379 (.o(n249363),
	.a(n249362),
	.b(regtop_g_mem_rd2_r[30]),
	.c(regtop_g_memr_ok_r));
   na02s01 U268380 (.o(n249374),
	.a(n249824),
	.b(regtop_g_dhs_r[13]));
   ao22s01 U268381 (.o(n249373),
	.a(FE_OFN546_n245460),
	.b(regtop_g_ari_r[1]),
	.c(FE_OFN400_n249836),
	.d(g_field_start_add_r[29]));
   ao22s01 U268382 (.o(n249372),
	.a(FE_OFN527_n249828),
	.b(regtop_g_fcho2_r[13]),
	.c(FE_OFN552_n245462),
	.d(regtop_g_pct_r[1]));
   in01s01 U268383 (.o(n252418),
	.a(regtop_g_fcho0_r[13]));
   ao12s01 U268384 (.o(n249367),
	.a(n249825),
	.b(regtop_g_mem_rd2_r[29]),
	.c(regtop_g_memr_ok_r));
   oa12s01 U268385 (.o(n249370),
	.a(n249367),
	.b(n249763),
	.c(n252418));
   in01s01 U268386 (.o(n252504),
	.a(regtop_g_fcho1_r[13]));
   ao22s01 U268387 (.o(n249368),
	.a(g_hsdc_r[5]),
	.b(n249786),
	.c(n249813),
	.d(regtop_g_vf_r[1]));
   oa12s01 U268388 (.o(n249369),
	.a(n249368),
	.b(n249375),
	.c(n252504));
   no02s01 U268389 (.o(n249371),
	.a(n249370),
	.b(n249369));
   ao22s01 U268390 (.o(n249383),
	.a(n249823),
	.b(regtop_g_hsv_r[10]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcho0_r[10]));
   na02s01 U268391 (.o(n249382),
	.a(FE_OFN400_n249836),
	.b(g_field_start_add_r[26]));
   ao22s01 U268392 (.o(n249381),
	.a(FE_OFN546_n245460),
	.b(regtop_g_frc_r[2]),
	.c(n249824),
	.d(regtop_g_dhs_r[10]));
   ao12f01 U268393 (.o(n249378),
	.a(n249825),
	.b(g_pcut_r[10]),
	.c(n249811));
   in01s01 U268394 (.o(n252394),
	.a(regtop_g_fcho2_r[10]));
   in01s01 U268395 (.o(n252501),
	.a(regtop_g_fcho1_r[10]));
   oa22s01 U268396 (.o(n249376),
	.a(n249828),
	.b(n252394),
	.c(n249375),
	.d(n252501));
   ao12s01 U268397 (.o(n249377),
	.a(n249376),
	.b(g_hsdc_r[2]),
	.c(n249786));
   na02s01 U268398 (.o(n249379),
	.a(FE_OFN462_n249378),
	.b(n249377));
   na02s01 U268399 (.o(n249387),
	.a(n249628),
	.b(regtop_g_hsv_r[9]));
   ao22f01 U268400 (.o(n249386),
	.a(n252944),
	.b(g_vldmode_r[0]),
	.c(n249768),
	.d(regtop_g_pis_r[1]));
   ao22f01 U268401 (.o(n249385),
	.a(FE_OFN396_n249640),
	.b(regtop_g_fcho0_r[9]),
	.c(n249639),
	.d(regtop_g_fcho2_r[9]));
   ao22f01 U268402 (.o(n249384),
	.a(FE_OFN392_n249635),
	.b(regtop_g_dhs_r[9]),
	.c(FE_OFN264_n249636),
	.d(regtop_g_tr_r[9]));
   ao22f01 U268403 (.o(n249391),
	.a(g_hsdc_r[1]),
	.b(FE_OFN398_n249646),
	.c(n252874),
	.d(g_pcut_r[9]));
   in01f03 U268404 (.o(n249543),
	.a(n249388));
   ao12s01 U268405 (.o(n249390),
	.a(n249543),
	.b(regtop_g_frc_r[1]),
	.c(n249629));
   ao22f02 U268406 (.o(n249389),
	.a(n249637),
	.b(regtop_g_fcho1_r[9]),
	.c(n252972),
	.d(g_field_start_add_r[25]));
   no02s01 U268407 (.o(n249395),
	.a(n249393),
	.b(n249392));
   na02f02 U268408 (.o(n249394),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[25]));
   oa12f01 U268409 (.o(n244982),
	.a(FE_OFN20_n249394),
	.b(FE_OFN575_n245444),
	.c(n249395));
   ao22s01 U268410 (.o(n249400),
	.a(FE_OFN396_n249640),
	.b(regtop_g_fcho0_r[6]),
	.c(n249637),
	.d(regtop_g_fcho1_r[6]));
   in01f04 U268411 (.o(n249634),
	.a(n249396));
   ao22s01 U268412 (.o(n249399),
	.a(FE_OFN392_n249635),
	.b(regtop_g_dhs_r[6]),
	.c(n249634),
	.d(regtop_g_tmc_r[22]));
   ao22s01 U268413 (.o(n249398),
	.a(FE_OFN264_n249636),
	.b(regtop_g_tr_r[6]),
	.c(n249639),
	.d(regtop_g_fcho2_r[6]));
   ao22f08 U268414 (.o(n249397),
	.a(regtop_g_nfst_r[22]),
	.b(n249584),
	.c(g_vsdc_r[6]),
	.d(FE_OFN398_n249646));
   ao12f02 U268415 (.o(n249404),
	.a(n249543),
	.b(g_pcut_r[6]),
	.c(n252874));
   ao22s01 U268416 (.o(n249403),
	.a(n249638),
	.b(regtop_g_cp_r[6]),
	.c(n249787),
	.d(regtop_g_fs_r[2]));
   na02s01 U268417 (.o(n249402),
	.a(n249628),
	.b(regtop_g_hsv_r[6]));
   na02f01 U268418 (.o(n249401),
	.a(n252972),
	.b(g_field_start_add_r[22]));
   na02f80 U268419 (.o(n249407),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[22]));
   ao22s01 U268420 (.o(n249412),
	.a(FE_OFN396_n249640),
	.b(regtop_g_fcho0_r[5]),
	.c(n249637),
	.d(regtop_g_fcho1_r[5]));
   ao22s01 U268421 (.o(n249411),
	.a(FE_OFN392_n249635),
	.b(regtop_g_dhs_r[5]),
	.c(n249634),
	.d(regtop_g_tmc_r[21]));
   ao22s01 U268422 (.o(n249410),
	.a(FE_OFN264_n249636),
	.b(regtop_g_tr_r[5]),
	.c(n249639),
	.d(regtop_g_fcho2_r[5]));
   na02f01 U268423 (.o(n249409),
	.a(g_vsdc_r[5]),
	.b(FE_OFN398_n249646));
   ao12f02 U268424 (.o(n249416),
	.a(n249543),
	.b(g_pcut_r[5]),
	.c(n252874));
   ao22f01 U268425 (.o(n249415),
	.a(n249638),
	.b(regtop_g_cp_r[5]),
	.c(FE_OFN266_n249787),
	.d(regtop_g_fs_r[1]));
   na02s01 U268426 (.o(n249414),
	.a(n249628),
	.b(regtop_g_hsv_r[5]));
   na02s01 U268427 (.o(n249413),
	.a(n252972),
	.b(g_field_start_add_r[21]));
   no02f02 U268428 (.o(n249420),
	.a(n249418),
	.b(n249417));
   na02f02 U268429 (.o(n249419),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[21]));
   oa12f02 U268430 (.o(n244980),
	.a(n249419),
	.b(FE_OFN575_n245444),
	.c(n249420));
   ao22s01 U268431 (.o(n249424),
	.a(n249639),
	.b(regtop_g_fcho2_r[2]),
	.c(n249637),
	.d(regtop_g_fcho1_r[2]));
   ao22s01 U268432 (.o(n249423),
	.a(FE_OFN392_n249635),
	.b(regtop_g_dhs_r[2]),
	.c(n249634),
	.d(regtop_g_tmc_r[18]));
   ao22s01 U268433 (.o(n249422),
	.a(g_vsdc_r[2]),
	.b(FE_OFN398_n249646),
	.c(FE_OFN264_n249636),
	.d(regtop_g_tr_r[2]));
   ao22f08 U268434 (.o(n249421),
	.a(n252874),
	.b(g_pcut_r[2]),
	.c(n249584),
	.d(regtop_g_nfst_r[18]));
   ao12s01 U268435 (.o(n249427),
	.a(n249543),
	.b(g_field_start_add_r[18]),
	.c(n252972));
   ao22s01 U268436 (.o(n249426),
	.a(n249638),
	.b(regtop_g_cp_r[2]),
	.c(FE_OFN396_n249640),
	.d(regtop_g_fcho0_r[2]));
   na02s01 U268437 (.o(n249425),
	.a(n249628),
	.b(regtop_g_hsv_r[2]));
   na02f03 U268438 (.o(n249431),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[18]));
   oa12f02 U268439 (.o(n244979),
	.a(n249431),
	.b(n245444),
	.c(n249432));
   na02s01 U268440 (.o(n249439),
	.a(g_vsdc_r[1]),
	.b(FE_OFN398_n249646));
   ao22s01 U268441 (.o(n249438),
	.a(g_fcyc_r[17]),
	.b(n252912),
	.c(n249584),
	.d(regtop_g_nfst_r[17]));
   ao12s01 U268442 (.o(n249437),
	.a(n249543),
	.b(regtop_g_cf_r[1]),
	.c(n249769));
   ao22f01 U268443 (.o(n249434),
	.a(n249628),
	.b(regtop_g_hsv_r[1]),
	.c(FE_OFN392_n249635),
	.d(regtop_g_dhs_r[1]));
   ao22f01 U268444 (.o(n249433),
	.a(n249634),
	.b(regtop_g_tmc_r[17]),
	.c(FE_OFN396_n249640),
	.d(regtop_g_fcho0_r[1]));
   na02f02 U268445 (.o(n249435),
	.a(n249434),
	.b(n249433));
   ao12f01 U268446 (.o(n249436),
	.a(n249435),
	.b(g_pcut_r[1]),
	.c(n252874));
   ao22s01 U268447 (.o(n249443),
	.a(n249639),
	.b(regtop_g_fcho2_r[1]),
	.c(n249637),
	.d(regtop_g_fcho1_r[1]));
   ao22f02 U268448 (.o(n249441),
	.a(n249663),
	.b(regtop_g_isfb_r),
	.c(regtop_g_icfb_r),
	.d(n249547));
   ao22s01 U268449 (.o(n249440),
	.a(FE_OFN264_n249636),
	.b(regtop_g_tr_r[1]),
	.c(n252972),
	.d(g_field_start_add_r[17]));
   ao22f01 U268450 (.o(n249456),
	.a(n249813),
	.b(regtop_g_tc_r[7]),
	.c(n249838),
	.d(regtop_g_fcvo1_r[15]));
   ao22s01 U268451 (.o(n249455),
	.a(n249812),
	.b(regtop_g_tmc_r[15]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcvo0_r[15]));
   ao22f01 U268452 (.o(n249449),
	.a(g_fcyc_r[15]),
	.b(n252912),
	.c(n252972),
	.d(g_field_start_add_r[15]));
   ao12s01 U268453 (.o(n249452),
	.a(n245444),
	.b(n249449),
	.c(n249448));
   in01s01 U268454 (.o(n252891),
	.a(g_mbc_en_r));
   ao22f01 U268455 (.o(n249450),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[15]),
	.c(FE_OFN527_n249828),
	.d(regtop_g_fcvo2_r[15]));
   oa12f01 U268456 (.o(n249451),
	.a(n249450),
	.b(n249827),
	.c(n252891));
   no02f02 U268457 (.o(n249453),
	.a(n249452),
	.b(n249451));
   ao22s01 U268458 (.o(n249460),
	.a(n249634),
	.b(regtop_g_tmc_r[14]),
	.c(n249637),
	.d(regtop_g_fcvo1_r[14]));
   ao22f01 U268459 (.o(n249459),
	.a(n249638),
	.b(regtop_g_tc_r[6]),
	.c(FE_OFN266_n249787),
	.d(regtop_g_ba_r[6]));
   ao22s01 U268460 (.o(n249458),
	.a(FE_OFN264_n249636),
	.b(regtop_g_vd_r[14]),
	.c(n249639),
	.d(regtop_g_fcvo2_r[14]));
   ao22f01 U268461 (.o(n249457),
	.a(g_hs60p_r[6]),
	.b(FE_OFN398_n249646),
	.c(n249652),
	.d(regtop_g_embh_adr_r[6]));
   ao22f02 U268462 (.o(n249463),
	.a(g_fcyc_r[14]),
	.b(n252912),
	.c(n249584),
	.d(regtop_g_nfst_r[14]));
   ao22s01 U268463 (.o(n249461),
	.a(n249629),
	.b(regtop_g_brv_r[14]),
	.c(FE_OFN396_n249640),
	.d(regtop_g_fcvo0_r[14]));
   no02s01 U268464 (.o(n249467),
	.a(n249465),
	.b(n249464));
   na02f03 U268465 (.o(n249466),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[14]));
   oa12f01 U268466 (.o(n244976),
	.a(n249466),
	.b(FE_OFN575_n245444),
	.c(n249467));
   ao22f01 U268467 (.o(n249471),
	.a(n249638),
	.b(regtop_g_tc_r[5]),
	.c(n249637),
	.d(regtop_g_fcvo1_r[13]));
   ao22s01 U268468 (.o(n249470),
	.a(FE_OFN396_n249640),
	.b(regtop_g_fcvo0_r[13]),
	.c(FE_OFN266_n249787),
	.d(regtop_g_ba_r[5]));
   ao22s01 U268469 (.o(n249469),
	.a(n252912),
	.b(g_fcyc_r[13]),
	.c(FE_OFN264_n249636),
	.d(regtop_g_vd_r[13]));
   ao22f01 U268470 (.o(n249468),
	.a(n249652),
	.b(regtop_g_embh_adr_r[5]),
	.c(n249584),
	.d(regtop_g_nfst_r[13]));
   ao22s01 U268471 (.o(n249474),
	.a(n249629),
	.b(regtop_g_brv_r[13]),
	.c(n249639),
	.d(regtop_g_fcvo2_r[13]));
   na02s01 U268472 (.o(n249472),
	.a(n252972),
	.b(g_field_start_add_r[13]));
   oa12s01 U268473 (.o(n244975),
	.a(n249478),
	.b(FE_OFN575_n245444),
	.c(n249479));
   ao22s01 U268474 (.o(n249483),
	.a(FE_OFN266_n249787),
	.b(regtop_g_ba_r[4]),
	.c(n249639),
	.d(regtop_g_fcvo2_r[12]));
   ao22s01 U268475 (.o(n249482),
	.a(FE_OFN396_n249640),
	.b(regtop_g_fcvo0_r[12]),
	.c(FE_OFN264_n249636),
	.d(regtop_g_vd_r[12]));
   ao22s01 U268476 (.o(n249481),
	.a(g_hs60p_r[4]),
	.b(FE_OFN398_n249646),
	.c(n252912),
	.d(g_fcyc_r[12]));
   ao22f01 U268477 (.o(n249480),
	.a(n249652),
	.b(regtop_g_embh_adr_r[4]),
	.c(n249584),
	.d(regtop_g_nfst_r[12]));
   na02f01 U268478 (.o(n249486),
	.a(n252972),
	.b(g_field_start_add_r[12]));
   ao22s01 U268479 (.o(n249485),
	.a(FE_OFN392_n249635),
	.b(regtop_g_dvs_r[12]),
	.c(n249637),
	.d(regtop_g_fcvo1_r[12]));
   ao22s01 U268480 (.o(n249484),
	.a(n249629),
	.b(regtop_g_brv_r[12]),
	.c(n249634),
	.d(regtop_g_tmc_r[12]));
   na02f02 U268481 (.o(n249490),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[12]));
   oa12f01 U268482 (.o(n244974),
	.a(n249490),
	.b(FE_OFN575_n245444),
	.c(n249491));
   ao22s01 U268483 (.o(n249494),
	.a(n249663),
	.b(regtop_g_isdc_r),
	.c(n252972),
	.d(g_field_start_add_r[11]));
   ao22f02 U268484 (.o(n249492),
	.a(g_hs60p_r[3]),
	.b(FE_OFN398_n249646),
	.c(g_fcyc_r[11]),
	.d(n252912));
   ao22s01 U268485 (.o(n249498),
	.a(n252998),
	.b(g_field_offset_r[11]),
	.c(n253014),
	.d(g_cbcr_offset_r[11]));
   ao22s01 U268486 (.o(n249497),
	.a(n249628),
	.b(regtop_g_vsv_r[11]),
	.c(n249629),
	.d(regtop_g_brv_r[11]));
   na02s01 U268487 (.o(n249496),
	.a(n249634),
	.b(regtop_g_tmc_r[11]));
   ao22s01 U268488 (.o(n249495),
	.a(n249635),
	.b(regtop_g_dvs_r[11]),
	.c(n249787),
	.d(regtop_g_ba_r[3]));
   ao22s01 U268489 (.o(n249502),
	.a(n249638),
	.b(regtop_g_tc_r[3]),
	.c(n249639),
	.d(regtop_g_fcvo2_r[11]));
   ao22s01 U268490 (.o(n249501),
	.a(n249640),
	.b(regtop_g_fcvo0_r[11]),
	.c(FE_OFN264_n249636),
	.d(regtop_g_vd_r[11]));
   ao22s01 U268491 (.o(n249500),
	.a(n249637),
	.b(regtop_g_fcvo1_r[11]),
	.c(n249584),
	.d(regtop_g_nfst_r[11]));
   ao22s01 U268492 (.o(n249499),
	.a(n249652),
	.b(regtop_g_embh_adr_r[3]),
	.c(n252874),
	.d(g_mbc_r[11]));
   na02s01 U268493 (.o(n249506),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[11]));
   oa12s01 U268494 (.o(n244973),
	.a(n249506),
	.b(n245444),
	.c(n249507));
   ao22f01 U268495 (.o(n249510),
	.a(n249663),
	.b(regtop_g_isuc_r),
	.c(n252998),
	.d(g_field_offset_r[10]));
   ao22s01 U268496 (.o(n249509),
	.a(n253014),
	.b(g_cbcr_offset_r[10]),
	.c(n249634),
	.d(regtop_g_tmc_r[10]));
   ao22s01 U268497 (.o(n249508),
	.a(n249628),
	.b(regtop_g_vsv_r[10]),
	.c(n249635),
	.d(regtop_g_dvs_r[10]));
   na02s01 U268498 (.o(n249515),
	.a(n249629),
	.b(regtop_g_brv_r[10]));
   ao22s01 U268499 (.o(n249514),
	.a(n249787),
	.b(regtop_g_ba_r[2]),
	.c(n249639),
	.d(regtop_g_fcvo2_r[10]));
   ao22s01 U268500 (.o(n249513),
	.a(n249638),
	.b(regtop_g_tc_r[2]),
	.c(FE_OFN264_n249636),
	.d(regtop_g_vd_r[10]));
   ao22s01 U268501 (.o(n249512),
	.a(n249640),
	.b(regtop_g_fcvo0_r[10]),
	.c(n249637),
	.d(regtop_g_fcvo1_r[10]));
   ao22s01 U268502 (.o(n249519),
	.a(g_fcyc_r[10]),
	.b(n252912),
	.c(n249547),
	.d(regtop_g_icuc_r));
   ao22s01 U268503 (.o(n249518),
	.a(n252874),
	.b(g_mbc_r[10]),
	.c(n249584),
	.d(regtop_g_nfst_r[10]));
   na02s01 U268504 (.o(n249517),
	.a(n249652),
	.b(regtop_g_embh_adr_r[2]));
   na02f02 U268505 (.o(n249516),
	.a(g_hs60p_r[2]),
	.b(FE_OFN398_n249646));
   na02f01 U268506 (.o(n249523),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[10]));
   ao22s01 U268507 (.o(n249528),
	.a(FE_OFN264_n249636),
	.b(regtop_g_vd_r[9]),
	.c(n249637),
	.d(regtop_g_fcvo1_r[9]));
   ao22f02 U268508 (.o(n249527),
	.a(n249663),
	.b(regtop_g_issw_r),
	.c(n249547),
	.d(regtop_g_icsw_r));
   na02f01 U268509 (.o(n249525),
	.a(n249584),
	.b(regtop_g_nfst_r[9]));
   ao22s01 U268510 (.o(n249532),
	.a(n252998),
	.b(g_field_offset_r[9]),
	.c(n249628),
	.d(regtop_g_vsv_r[9]));
   na02s01 U268511 (.o(n249531),
	.a(n249634),
	.b(regtop_g_tmc_r[9]));
   ao22s01 U268512 (.o(n249530),
	.a(n249630),
	.b(regtop_g_vbsv_r[9]),
	.c(n249629),
	.d(regtop_g_brv_r[9]));
   ao22f02 U268513 (.o(n249529),
	.a(FE_OFN392_n249635),
	.b(regtop_g_dvs_r[9]),
	.c(n249787),
	.d(regtop_g_ba_r[1]));
   ao22f01 U268514 (.o(n249536),
	.a(FE_OFN396_n249640),
	.b(regtop_g_fcvo0_r[9]),
	.c(n249639),
	.d(regtop_g_fcvo2_r[9]));
   ao22f01 U268515 (.o(n249535),
	.a(g_hs60p_r[1]),
	.b(FE_OFN398_n249646),
	.c(n249638),
	.d(regtop_g_tc_r[1]));
   ao22f01 U268516 (.o(n249534),
	.a(n249582),
	.b(regtop_g_fbst_r[9]),
	.c(n252874),
	.d(g_mbc_r[9]));
   ao22f01 U268517 (.o(n249533),
	.a(n252912),
	.b(g_fcyc_r[9]),
	.c(n249652),
	.d(regtop_g_embh_adr_r[1]));
   na04f03 U268518 (.o(n249537),
	.a(n249536),
	.b(n249535),
	.c(n249534),
	.d(n249533));
   na02s01 U268519 (.o(n249540),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[9]));
   ao22s01 U268520 (.o(n249546),
	.a(g_hs60p_r[0]),
	.b(FE_OFN398_n249646),
	.c(g_init_vld_r_s),
	.d(n249542));
   ao22s01 U268521 (.o(n249545),
	.a(regtop_g_dmod_r),
	.b(n252944),
	.c(n249543),
	.d(regtop_g_vldstatus_r[4]));
   na02s01 U268522 (.o(n249544),
	.a(n252912),
	.b(g_fcyc_r[8]));
   na03f03 U268523 (.o(n249564),
	.a(n249546),
	.b(n249545),
	.c(n249544));
   ao22f02 U268524 (.o(n249552),
	.a(n249663),
	.b(regtop_g_issr_r),
	.c(n249547),
	.d(regtop_g_icsr_r));
   ao22f02 U268525 (.o(n249551),
	.a(regtop_g_rff_r),
	.b(n249768),
	.c(n252998),
	.d(g_field_offset_r[8]));
   na02s01 U268526 (.o(n249549),
	.a(regtop_g_vsv_r[8]),
	.b(n249628));
   ao22s01 U268527 (.o(n249556),
	.a(regtop_g_vbsv_r[8]),
	.b(n249630),
	.c(regtop_g_dvs_r[8]),
	.d(n249635));
   ao22s01 U268528 (.o(n249555),
	.a(regtop_g_brv_r[8]),
	.b(n249629),
	.c(regtop_g_ld_r),
	.d(n249769));
   ao22s01 U268529 (.o(n249554),
	.a(regtop_g_tmc_r[8]),
	.b(n249634),
	.c(regtop_g_tc_r[0]),
	.d(n249638));
   ao22s01 U268530 (.o(n249553),
	.a(regtop_g_fcvo0_r[8]),
	.b(n249640),
	.c(regtop_g_ba_r[0]),
	.d(n249787));
   na02s01 U268531 (.o(n249559),
	.a(regtop_g_fcvo1_r[8]),
	.b(n249637));
   na02s01 U268532 (.o(n249558),
	.a(regtop_g_embh_adr_r[0]),
	.b(n249652));
   ao22s01 U268533 (.o(n249557),
	.a(n252874),
	.b(g_mbc_r[8]),
	.c(regtop_g_nfst_r[8]),
	.d(n249584));
   na02f01 U268534 (.o(n249565),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[8]));
   in01f01 U268535 (.o(n249589),
	.a(n253014));
   no02s01 U268536 (.o(n249579),
	.a(n249589),
	.b(n253022));
   in01s01 U268537 (.o(n252930),
	.a(g_fcyc_r[7]));
   na02s01 U268538 (.o(n249567),
	.a(n249584),
	.b(regtop_g_nfst_r[7]));
   oa12f02 U268539 (.o(n249578),
	.a(n249567),
	.b(n252930),
	.c(FE_OFN544_n252912));
   ao22s01 U268540 (.o(n249571),
	.a(n249787),
	.b(regtop_g_scp_r[7]),
	.c(FE_OFN264_n249636),
	.d(regtop_g_vd_r[7]));
   ao22s01 U268541 (.o(n249570),
	.a(n249635),
	.b(regtop_g_dvs_r[7]),
	.c(n249638),
	.d(regtop_g_mc_r[7]));
   ao22s01 U268542 (.o(n249569),
	.a(n249639),
	.b(regtop_g_fcvo2_r[7]),
	.c(n249637),
	.d(regtop_g_fcvo1_r[7]));
   na02f01 U268543 (.o(n249568),
	.a(n252998),
	.b(g_field_offset_r[7]));
   ao22s01 U268544 (.o(n249575),
	.a(n249630),
	.b(regtop_g_vbsv_r[7]),
	.c(n249629),
	.d(regtop_g_brv_r[7]));
   ao22s01 U268545 (.o(n249574),
	.a(n249628),
	.b(regtop_g_vsv_r[7]),
	.c(n249640),
	.d(regtop_g_fcvo0_r[7]));
   ao22s01 U268546 (.o(n249573),
	.a(n249769),
	.b(regtop_g_pali_r[7]),
	.c(n249634),
	.d(regtop_g_tmc_r[7]));
   ao22f02 U268547 (.o(n249572),
	.a(n249582),
	.b(regtop_g_fbst_r[7]),
	.c(n252874),
	.d(g_mbc_r[7]));
   na02s01 U268548 (.o(n249580),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[7]));
   oa12f03 U268549 (.o(n244969),
	.a(n249580),
	.b(n245444),
	.c(n249581));
   ao22s01 U268550 (.o(n249606),
	.a(g_vs60p_r[6]),
	.b(n249786),
	.c(FE_OFN527_n249828),
	.d(regtop_g_fcvo2_r[6]));
   in01f01 U268551 (.o(n249649),
	.a(n249582));
   no02f02 U268552 (.o(n249744),
	.a(n245444),
	.b(n249649));
   na02s01 U268553 (.o(n249615),
	.a(FE_OFN4_n245443),
	.b(n249652));
   in01f01 U268554 (.o(n249746),
	.a(n249615));
   ao22f02 U268555 (.o(n249605),
	.a(regtop_g_fbst_r[6]),
	.b(n249744),
	.c(n249746),
	.d(regtop_g_embv_adr_r[6]));
   in01s01 U268556 (.o(n252884),
	.a(g_mbc_r[6]));
   na02s01 U268557 (.o(n249585),
	.a(FE_OFN4_n245443),
	.b(n249584));
   in01f01 U268558 (.o(n249713),
	.a(n249585));
   ao22s01 U268559 (.o(n249586),
	.a(g_fcyc_r[6]),
	.b(n249841),
	.c(n249713),
	.d(regtop_g_nfst_r[6]));
   in01s01 U268560 (.o(n249602),
	.a(n249586));
   na02s01 U268561 (.o(n249587),
	.a(FE_OFN4_n245443),
	.b(n249630));
   in01f01 U268562 (.o(n249733),
	.a(n249587));
   ao22s01 U268563 (.o(n249595),
	.a(n249729),
	.b(regtop_g_udb_cpu_r[6]),
	.c(n249733),
	.d(regtop_g_vbsv_r[6]));
   na02s01 U268564 (.o(n249594),
	.a(n249728),
	.b(regtop_g_adb_cpu_r[6]));
   in01f01 U268565 (.o(n249627),
	.a(n252998));
   no02f02 U268566 (.o(n249732),
	.a(n245444),
	.b(n249589));
   ao22s01 U268567 (.o(n249593),
	.a(n249731),
	.b(g_field_offset_r[6]),
	.c(n249732),
	.d(g_cbcr_offset_r[6]));
   na02s01 U268568 (.o(n249590),
	.a(FE_OFN4_n245443),
	.b(n249769));
   in01f01 U268569 (.o(n249739),
	.a(n249590));
   na02f01 U268570 (.o(n249591),
	.a(FE_OFN4_n245443),
	.b(FE_OFN266_n249787));
   in01f02 U268571 (.o(n249757),
	.a(n249591));
   ao22f01 U268572 (.o(n249592),
	.a(n249739),
	.b(regtop_g_pali_r[6]),
	.c(n249757),
	.d(regtop_g_scp_r[6]));
   ao22s01 U268573 (.o(n249598),
	.a(n249813),
	.b(regtop_g_mc_r[6]),
	.c(n249823),
	.d(regtop_g_vsv_r[6]));
   ao22f01 U268574 (.o(n249597),
	.a(FE_OFN545_n245460),
	.b(regtop_g_brv_r[6]),
	.c(n249824),
	.d(regtop_g_dvs_r[6]));
   ao22f01 U268575 (.o(n249596),
	.a(n249838),
	.b(regtop_g_fcvo1_r[6]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcvo0_r[6]));
   ao22s01 U268576 (.o(n249626),
	.a(g_vs60p_r[5]),
	.b(n249786),
	.c(g_fcyc_r[5]),
	.d(n249841));
   na02s01 U268577 (.o(n249696),
	.a(FE_OFN4_n245443),
	.b(n249647));
   in01s01 U268578 (.o(n249712),
	.a(n249696));
   ao22f01 U268579 (.o(n249625),
	.a(regtop_g_fbst_r[5]),
	.b(n249744),
	.c(regtop_g_fpst_r[5]),
	.d(n249712));
   ao22f02 U268580 (.o(n249609),
	.a(regtop_g_adb_cpu_r[5]),
	.b(n249728),
	.c(regtop_g_vbsv_r[5]),
	.d(n249733));
   ao22f01 U268581 (.o(n249608),
	.a(n249811),
	.b(g_mbc_r[5]),
	.c(regtop_g_nfst_r[5]),
	.d(n249713));
   na02f01 U268582 (.o(n249607),
	.a(regtop_g_udb_cpu_r[5]),
	.b(n249729));
   na02f01 U268583 (.o(n249613),
	.a(regtop_g_pali_r[5]),
	.b(n249739));
   ao22f02 U268584 (.o(n249612),
	.a(g_field_offset_r[5]),
	.b(n249731),
	.c(g_cbcr_offset_r[5]),
	.d(n249732));
   ao22f01 U268585 (.o(n249610),
	.a(FE_OFN552_n245462),
	.b(regtop_g_vd_r[5]),
	.c(n249823),
	.d(regtop_g_vsv_r[5]));
   in01s01 U268586 (.o(n249616),
	.a(regtop_g_embv_adr_r[5]));
   ao22f02 U268587 (.o(n249614),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[5]),
	.c(n249825),
	.d(regtop_g_vldstatus_r[1]));
   oa12s01 U268588 (.o(n249621),
	.a(n249614),
	.b(n249616),
	.c(n249615));
   ao22s01 U268589 (.o(n249619),
	.a(n249813),
	.b(regtop_g_mc_r[5]),
	.c(n249824),
	.d(regtop_g_dvs_r[5]));
   ao22s01 U268590 (.o(n249617),
	.a(FE_OFN527_n249828),
	.b(regtop_g_fcvo2_r[5]),
	.c(n249838),
	.d(regtop_g_fcvo1_r[5]));
   in01s01 U268591 (.o(n253001),
	.a(g_field_offset_r[3]));
   no02f01 U268592 (.o(n249660),
	.a(n249627),
	.b(n253001));
   ao22s01 U268593 (.o(n249633),
	.a(n253014),
	.b(g_cbcr_offset_r[3]),
	.c(n249628),
	.d(regtop_g_vsv_r[3]));
   na02s01 U268594 (.o(n249632),
	.a(n249629),
	.b(regtop_g_brv_r[3]));
   ao22m01 U268595 (.o(n249631),
	.a(n249630),
	.b(regtop_g_vbsv_r[3]),
	.c(n249769),
	.d(regtop_g_pali_r[3]));
   na03f04 U268596 (.o(n249659),
	.a(n249633),
	.b(n249632),
	.c(n249631));
   ao22f02 U268597 (.o(n249644),
	.a(FE_OFN392_n249635),
	.b(regtop_g_dvs_r[3]),
	.c(n249634),
	.d(regtop_g_tmc_r[3]));
   ao22s01 U268598 (.o(n249643),
	.a(n249787),
	.b(regtop_g_scp_r[3]),
	.c(FE_OFN264_n249636),
	.d(regtop_g_vd_r[3]));
   ao22s01 U268599 (.o(n249642),
	.a(n249638),
	.b(regtop_g_mc_r[3]),
	.c(n249637),
	.d(regtop_g_fcvo1_r[3]));
   ao22s01 U268600 (.o(n249641),
	.a(n249640),
	.b(regtop_g_fcvo0_r[3]),
	.c(n249639),
	.d(regtop_g_fcvo2_r[3]));
   ao22s01 U268601 (.o(n249656),
	.a(g_vs60p_r[3]),
	.b(FE_OFN398_n249646),
	.c(n249645),
	.d(regtop_g_adb_cpu_r[3]));
   ao22m02 U268602 (.o(n249655),
	.a(n249647),
	.b(regtop_g_fpst_r[3]),
	.c(n252874),
	.d(g_mbc_r[3]));
   na02s01 U268603 (.o(n249654),
	.a(regtop_g_udb_cpu_r[3]),
	.b(n249648));
   in01s01 U268604 (.o(n252936),
	.a(g_fcyc_r[3]));
   in01s01 U268605 (.o(n252293),
	.a(regtop_g_fbst_r[3]));
   oa22f01 U268606 (.o(n249651),
	.a(n252936),
	.b(FE_OFN544_n252912),
	.c(n249649),
	.d(n252293));
   ao12f01 U268607 (.o(n249653),
	.a(n249651),
	.b(n249652),
	.c(regtop_g_embv_adr_r[3]));
   na02f40 U268608 (.o(n249661),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[3]));
   ao22s01 U268609 (.o(n249684),
	.a(n249811),
	.b(g_mbc_r[2]),
	.c(n249746),
	.d(regtop_g_embv_adr_r[2]));
   na02s01 U268610 (.o(n249686),
	.a(n249663),
	.b(FE_OFN4_n245443));
   in01s01 U268611 (.o(n249738),
	.a(n249686));
   no02f01 U268612 (.o(n249730),
	.a(n245444),
	.b(n252958));
   ao22f01 U268613 (.o(n249667),
	.a(n249728),
	.b(regtop_g_adb_cpu_r[2]),
	.c(regtop_g_icpi_r),
	.d(n249730));
   ao22f01 U268614 (.o(n249666),
	.a(n249729),
	.b(regtop_g_udb_cpu_r[2]),
	.c(n249739),
	.d(regtop_g_pali_r[2]));
   na02f06 U268615 (.o(n249665),
	.a(n249733),
	.b(regtop_g_vbsv_r[2]));
   ao22f02 U268616 (.o(n249670),
	.a(FE_OFN552_n245462),
	.b(regtop_g_vd_r[2]),
	.c(n249823),
	.d(regtop_g_vsv_r[2]));
   ao22f01 U268617 (.o(n249669),
	.a(n249813),
	.b(regtop_g_mc_r[2]),
	.c(n249824),
	.d(regtop_g_dvs_r[2]));
   na02f01 U268618 (.o(n249673),
	.a(g_vs60p_r[2]),
	.b(n249786));
   in01f01 U268619 (.o(n249679),
	.a(n249673));
   ao22f02 U268620 (.o(n249677),
	.a(n249838),
	.b(regtop_g_fcvo1_r[2]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcvo0_r[2]));
   ao22f01 U268621 (.o(n249676),
	.a(FE_OFN527_n249828),
	.b(regtop_g_fcvo2_r[2]),
	.c(FE_OFN545_n245460),
	.d(regtop_g_brv_r[2]));
   na02f01 U268622 (.o(n249675),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[2]));
   na02s01 U268623 (.o(n249674),
	.a(n249712),
	.b(regtop_g_fpst_r[2]));
   in01s01 U268624 (.o(n252266),
	.a(regtop_g_isph_r));
   oa12s01 U268625 (.o(n249687),
	.a(n249685),
	.b(n252266),
	.c(n249686));
   ao22f04 U268626 (.o(n249710),
	.a(n249811),
	.b(g_mbc_r[1]),
	.c(n249744),
	.d(regtop_g_fbst_r[1]));
   ao22s01 U268627 (.o(n249691),
	.a(n249728),
	.b(regtop_g_adb_cpu_r[1]),
	.c(n249730),
	.d(regtop_g_icph_r));
   ao22s01 U268628 (.o(n249690),
	.a(n249729),
	.b(regtop_g_udb_cpu_r[1]),
	.c(n249739),
	.d(regtop_g_pali_r[1]));
   ao22s01 U268629 (.o(n249688),
	.a(n249731),
	.b(g_field_offset_r[1]),
	.c(n249732),
	.d(g_cbcr_offset_r[1]));
   ao22f01 U268630 (.o(n249694),
	.a(n249824),
	.b(regtop_g_dvs_r[1]),
	.c(n249823),
	.d(regtop_g_vsv_r[1]));
   ao22s01 U268631 (.o(n249693),
	.a(n249813),
	.b(regtop_g_mc_r[1]),
	.c(FE_OFN552_n245462),
	.d(regtop_g_vd_r[1]));
   ao22f02 U268632 (.o(n249692),
	.a(FE_OFN527_n249828),
	.b(regtop_g_fcvo2_r[1]),
	.c(FE_OFN545_n245460),
	.d(regtop_g_brv_r[1]));
   in01s01 U268633 (.o(n252841),
	.a(g_vs60p_r[1]));
   in01s01 U268634 (.o(n252751),
	.a(regtop_g_fpst_r[1]));
   oa22s01 U268635 (.o(n249706),
	.a(n252841),
	.b(n249829),
	.c(n249696),
	.d(n252751));
   ao22f01 U268636 (.o(n249704),
	.a(n249838),
	.b(regtop_g_fcvo1_r[1]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcvo0_r[1]));
   ao22s01 U268637 (.o(n249703),
	.a(n249841),
	.b(g_fcyc_r[1]),
	.c(n249713),
	.d(regtop_g_nfst_r[1]));
   no03f03 U268638 (.o(n249745),
	.a(n249698),
	.b(n245444),
	.c(n249697));
   ao22s01 U268639 (.o(n249702),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[1]),
	.c(regtop_g_nfco_r[1]),
	.d(n249745));
   na02s01 U268640 (.o(n249699),
	.a(FE_OFN4_n245443),
	.b(n252944));
   in01s01 U268641 (.o(n249700),
	.a(n249699));
   na02s01 U268642 (.o(n249701),
	.a(g_bmod_r),
	.b(n249700));
   ao22s01 U268643 (.o(n249756),
	.a(FE_OFN545_n245460),
	.b(regtop_g_brv_r[0]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcvo0_r[0]));
   ao22f01 U268644 (.o(n249755),
	.a(n249712),
	.b(regtop_g_fpst_r[0]),
	.c(n249841),
	.d(g_fcyc_r[0]));
   ao22f01 U268645 (.o(n249715),
	.a(g_vs60p_r[0]),
	.b(n249786),
	.c(n249713),
	.d(regtop_g_nfst_r[0]));
   na02s01 U268646 (.o(n249714),
	.a(FE_OFN527_n249828),
	.b(regtop_g_fcvo2_r[0]));
   na02s01 U268647 (.o(n249716),
	.a(n249715),
	.b(n249714));
   ao12f02 U268648 (.o(n249754),
	.a(n249716),
	.b(regtop_g_mem_rd2_r[0]),
	.c(regtop_g_memr_ok_r));
   ao22s01 U268649 (.o(n249727),
	.a(n249768),
	.b(regtop_g_pf_r),
	.c(n249717),
	.d(g_line_offset_r));
   oa12s01 U268650 (.o(n249724),
	.a(n249719),
	.b(n245083),
	.c(n249720));
   ao12s01 U268651 (.o(n249722),
	.a(n249721),
	.b(regtop_g_imod_r),
	.c(n252944));
   oa12f02 U268652 (.o(n249723),
	.a(n249722),
	.b(g_swrst_r_n),
	.c(n249771));
   ao22s01 U268653 (.o(n249737),
	.a(n249729),
	.b(regtop_g_udb_cpu_r[0]),
	.c(n249728),
	.d(regtop_g_adb_cpu_r[0]));
   na02s01 U268654 (.o(n249735),
	.a(n249732),
	.b(g_cbcr_offset_r[0]));
   ao22s01 U268655 (.o(n249734),
	.a(n249838),
	.b(regtop_g_fcvo1_r[0]),
	.c(n249733),
	.d(regtop_g_vbsv_r[0]));
   ao22s01 U268656 (.o(n249742),
	.a(n249757),
	.b(regtop_g_scp_r[0]),
	.c(n249738),
	.d(regtop_g_issh_r));
   ao22s01 U268657 (.o(n249741),
	.a(FE_OFN552_n245462),
	.b(regtop_g_vd_r[0]),
	.c(n249739),
	.d(regtop_g_pali_r[0]));
   ao22s01 U268658 (.o(n249747),
	.a(n249746),
	.b(regtop_g_embv_adr_r[0]),
	.c(n249745),
	.d(regtop_g_nfco_r[0]));
   ao22s01 U268659 (.o(n249767),
	.a(g_hsdc_r[4]),
	.b(n249786),
	.c(n249757),
	.d(regtop_g_cdf_r));
   ao22f01 U268660 (.o(n249761),
	.a(n249824),
	.b(regtop_g_dhs_r[12]),
	.c(FE_OFN400_n249836),
	.d(g_field_start_add_r[28]));
   ao22s01 U268661 (.o(n249760),
	.a(FE_OFN552_n245462),
	.b(regtop_g_pct_r[0]),
	.c(n249812),
	.d(regtop_g_cg_r));
   ao22s01 U268662 (.o(n249759),
	.a(n249813),
	.b(regtop_g_vf_r[0]),
	.c(FE_OFN546_n245460),
	.d(regtop_g_ari_r[0]));
   ao22f01 U268663 (.o(n249758),
	.a(FE_OFN527_n249828),
	.b(regtop_g_fcho2_r[12]),
	.c(n249838),
	.d(regtop_g_fcho1_r[12]));
   in01s01 U268664 (.o(n252417),
	.a(regtop_g_fcho0_r[12]));
   ao12f01 U268665 (.o(n249762),
	.a(n249825),
	.b(regtop_g_mem_rd2_r[28]),
	.c(regtop_g_memr_ok_r));
   oa12s01 U268666 (.o(n249764),
	.a(n249762),
	.b(n249763),
	.c(n252417));
   na02f01 U268667 (.o(n244221),
	.a(n249767),
	.b(n249766));
   ao12s01 U268668 (.o(n249785),
	.a(n249825),
	.b(regtop_g_fcho0_r[8]),
	.c(FE_OFN489_n249763));
   ao22s01 U268669 (.o(n249780),
	.a(n252944),
	.b(g_vldmode_r[1]),
	.c(n249768),
	.d(regtop_g_pis_r[0]));
   ao22s01 U268670 (.o(n249779),
	.a(FE_OFN266_n249787),
	.b(regtop_g_va_r),
	.c(n252972),
	.d(g_field_start_add_r[24]));
   in01s01 U268671 (.o(n252828),
	.a(g_vden_r));
   na02s01 U268672 (.o(n249774),
	.a(n249838),
	.b(regtop_g_fcho1_r[8]));
   ao12s01 U268673 (.o(n249783),
	.a(n249664),
	.b(n249812),
	.c(regtop_g_bl_r));
   na02f01 U268674 (.o(n249782),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[24]));
   ao22f01 U268675 (.o(n249800),
	.a(g_vsdc_r[4]),
	.b(n249786),
	.c(n249811),
	.d(g_pcut_r[4]));
   ao22s01 U268676 (.o(n249799),
	.a(n249813),
	.b(regtop_g_cp_r[4]),
	.c(n249838),
	.d(regtop_g_fcho1_r[4]));
   ao12s01 U268677 (.o(n249798),
	.a(n249664),
	.b(FE_OFN527_n249828),
	.c(regtop_g_fcho2_r[4]));
   ao22s01 U268678 (.o(n249795),
	.a(FE_OFN552_n245462),
	.b(regtop_g_tr_r[4]),
	.c(n249812),
	.d(regtop_g_tmc_r[20]));
   ao22s01 U268679 (.o(n249794),
	.a(n249824),
	.b(regtop_g_dhs_r[4]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcho0_r[4]));
   in01s01 U268680 (.o(n252982),
	.a(g_field_start_add_r[20]));
   na02s01 U268681 (.o(n249788),
	.a(n249787),
	.b(regtop_g_fs_r[0]));
   oa12s01 U268682 (.o(n249791),
	.a(n249788),
	.b(n249789),
	.c(n252982));
   ao12s01 U268683 (.o(n249793),
	.a(n249825),
	.b(n249791),
	.c(FE_OFN4_n245443));
   ao22s01 U268684 (.o(n249792),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[20]),
	.c(n249823),
	.d(regtop_g_hsv_r[4]));
   ao12s01 U268685 (.o(n249810),
	.a(n249825),
	.b(regtop_g_mem_rd2_r[19]),
	.c(regtop_g_memr_ok_r));
   ao22s01 U268686 (.o(n249809),
	.a(FE_OFN527_n249828),
	.b(regtop_g_fcho2_r[3]),
	.c(n249813),
	.d(regtop_g_cp_r[3]));
   no02s01 U268687 (.o(n249806),
	.a(n252854),
	.b(n249829));
   ao22s01 U268688 (.o(n249804),
	.a(FE_OFN552_n245462),
	.b(regtop_g_tr_r[3]),
	.c(n249812),
	.d(regtop_g_tmc_r[19]));
   ao12s01 U268689 (.o(n249803),
	.a(n249664),
	.b(g_field_start_add_r[19]),
	.c(FE_OFN400_n249836));
   ao22s01 U268690 (.o(n249802),
	.a(n249838),
	.b(regtop_g_fcho1_r[3]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcho0_r[3]));
   ao22s01 U268691 (.o(n249801),
	.a(n249824),
	.b(regtop_g_dhs_r[3]),
	.c(n249823),
	.d(regtop_g_hsv_r[3]));
   na02s01 U268692 (.o(n249807),
	.a(n249811),
	.b(g_pcut_r[3]));
   na02s01 U268693 (.o(n249822),
	.a(n249823),
	.b(regtop_g_hsv_r[7]));
   ao22f01 U268694 (.o(n249821),
	.a(regtop_g_memr_ok_r),
	.b(regtop_g_mem_rd2_r[23]),
	.c(n249811),
	.d(g_pcut_r[7]));
   ao22s01 U268695 (.o(n249818),
	.a(n249812),
	.b(regtop_g_tmc_r[23]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcho0_r[7]));
   ao22s01 U268696 (.o(n249817),
	.a(n249813),
	.b(regtop_g_cp_r[7]),
	.c(n249838),
	.d(regtop_g_fcho1_r[7]));
   ao22s01 U268697 (.o(n249816),
	.a(FE_OFN527_n249828),
	.b(regtop_g_fcho2_r[7]),
	.c(FE_OFN552_n245462),
	.d(regtop_g_tr_r[7]));
   ao22s01 U268698 (.o(n249815),
	.a(n249824),
	.b(regtop_g_dhs_r[7]),
	.c(n249836),
	.d(g_field_start_add_r[23]));
   ao22s01 U268699 (.o(n249835),
	.a(n249824),
	.b(regtop_g_dhs_r[11]),
	.c(n249823),
	.d(regtop_g_hsv_r[11]));
   ao22f01 U268700 (.o(n249834),
	.a(FE_OFN547_n245460),
	.b(regtop_g_frc_r[3]),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcho0_r[11]));
   ao22f01 U268701 (.o(n249833),
	.a(n249838),
	.b(regtop_g_fcho1_r[11]),
	.c(FE_OFN400_n249836),
	.d(g_field_start_add_r[27]));
   ao12s01 U268702 (.o(n249826),
	.a(n249825),
	.b(regtop_g_mem_rd2_r[27]),
	.c(regtop_g_memr_ok_r));
   oa12f01 U268703 (.o(n249831),
	.a(n249826),
	.b(n249827),
	.c(n252908));
   in01s01 U268704 (.o(n252859),
	.a(g_hsdc_r[3]));
   in01s01 U268705 (.o(n252395),
	.a(regtop_g_fcho2_r[11]));
   oa22s01 U268706 (.o(n249830),
	.a(n252859),
	.b(n249829),
	.c(n249828),
	.d(n252395));
   ao12f02 U268707 (.o(n249845),
	.a(n249664),
	.b(regtop_g_memr_ok_r),
	.c(regtop_g_mem_rd2_r[31]));
   ao22f01 U268708 (.o(n249844),
	.a(FE_OFN546_n245460),
	.b(regtop_g_ari_r[3]),
	.c(FE_OFN400_n249836),
	.d(g_field_start_add_r[31]));
   ao22s01 U268709 (.o(n249843),
	.a(FE_OFN527_n249828),
	.b(regtop_g_fcho2_r[15]),
	.c(n249838),
	.d(regtop_g_fcho1_r[15]));
   ao22s01 U268710 (.o(n249842),
	.a(g_fcyc_en_r),
	.b(n249841),
	.c(FE_OFN489_n249763),
	.d(regtop_g_fcho0_r[15]));
   in01s01 U268711 (.o(n243097),
	.a(wbb_we_i));
   in01s01 U268712 (.o(n243096),
	.a(wbb_stb_i));
   in01s01 U268713 (.o(n252880),
	.a(regtop_g_wd_r[10]));
   ao12s01 U268714 (.o(n249846),
	.a(n252269),
	.b(n252270),
	.c(regtop_g_wd_r[10]));
   na02s01 U268715 (.o(n249847),
	.a(regtop_g_isuc_r),
	.b(n249846));
   oa12s01 U268716 (.o(n157815),
	.a(n249847),
	.b(n252273),
	.c(n252880));
   na02s01 U268717 (.o(n249854),
	.a(n253125),
	.b(vh_1_ph_add[9]));
   in01s01 U268718 (.o(n249903),
	.a(vh_1_ph_add[2]));
   in01s01 U268719 (.o(n249886),
	.a(vh_1_ph_add[4]));
   in01s01 U268720 (.o(n249850),
	.a(busrtop_b_rreq_vrh_add1_r[9]));
   no02s01 U268721 (.o(n249851),
	.a(n249913),
	.b(n249850));
   in01s01 U268722 (.o(n249852),
	.a(n249851));
   na02s01 U268723 (.o(n249862),
	.a(n253125),
	.b(vh_1_ph_add[8]));
   in01s01 U268724 (.o(n249858),
	.a(busrtop_b_rreq_vrh_add1_r[8]));
   no02s01 U268725 (.o(n249859),
	.a(n249913),
	.b(n249858));
   in01s01 U268726 (.o(n249860),
	.a(n249859));
   in01s01 U268727 (.o(n249867),
	.a(n249864));
   in01s01 U268728 (.o(n249865),
	.a(busrtop_b_rreq_vrh_add1_r[7]));
   no02s01 U268729 (.o(n249866),
	.a(n249913),
	.b(n249865));
   na02s01 U268730 (.o(n249877),
	.a(n253125),
	.b(vh_1_ph_add[6]));
   no02s01 U268731 (.o(n249874),
	.a(n249913),
	.b(n249873));
   in01s01 U268732 (.o(n249875),
	.a(n249874));
   na02s01 U268733 (.o(n249884),
	.a(n253125),
	.b(vh_1_ph_add[5]));
   oa12s01 U268734 (.o(n249879),
	.a(n249878),
	.b(n249885),
	.c(vh_1_ph_add[5]));
   in01s01 U268735 (.o(n249882),
	.a(n249879));
   in01s01 U268736 (.o(n249880),
	.a(busrtop_b_rreq_vrh_add1_r[5]));
   no02s01 U268737 (.o(n249881),
	.a(n249913),
	.b(n249880));
   na02s01 U268738 (.o(n157835),
	.a(n249884),
	.b(n249883));
   na02s01 U268739 (.o(n249892),
	.a(n253125),
	.b(vh_1_ph_add[4]));
   na02s01 U268740 (.o(n249891),
	.a(n249916),
	.b(n249887));
   no02s01 U268741 (.o(n249889),
	.a(n249913),
	.b(n249888));
   in01s01 U268742 (.o(n249890),
	.a(n249889));
   na02s01 U268743 (.o(n249901),
	.a(n253125),
	.b(vh_1_ph_add[3]));
   oa12s01 U268744 (.o(n249894),
	.a(n249893),
	.b(n249902),
	.c(vh_1_ph_add[3]));
   in01s01 U268745 (.o(n249895),
	.a(n249894));
   na02s01 U268746 (.o(n249896),
	.a(n249916),
	.b(n249895));
   in01s01 U268747 (.o(n249899),
	.a(n249896));
   in01s01 U268748 (.o(n249897),
	.a(busrtop_b_rreq_vrh_add1_r[3]));
   no02s01 U268749 (.o(n249898),
	.a(n249897),
	.b(n249913));
   no02s01 U268750 (.o(n249900),
	.a(n249899),
	.b(n249898));
   na02s01 U268751 (.o(n157837),
	.a(n249901),
	.b(n249900));
   na02s01 U268752 (.o(n249909),
	.a(n253125),
	.b(vh_1_ph_add[2]));
   ao12s01 U268753 (.o(n249904),
	.a(n249902),
	.b(n249910),
	.c(n249903));
   na02s01 U268754 (.o(n249908),
	.a(n249916),
	.b(n249904));
   in01s01 U268755 (.o(n249905),
	.a(busrtop_b_rreq_vrh_add1_r[2]));
   no02s01 U268756 (.o(n249906),
	.a(n249913),
	.b(n249905));
   in01s01 U268757 (.o(n249907),
	.a(n249906));
   na03s01 U268758 (.o(n157838),
	.a(n249909),
	.b(n249908),
	.c(n249907));
   oa12s01 U268759 (.o(n249911),
	.a(n249910),
	.b(vh_1_ph_add[0]),
	.c(vh_1_ph_add[1]));
   in01s01 U268760 (.o(n249915),
	.a(n249911));
   no02s01 U268761 (.o(n249914),
	.a(n249913),
	.b(n249912));
   ao12s01 U268762 (.o(n249917),
	.a(n249914),
	.b(n249916),
	.c(n249915));
   na02s01 U268763 (.o(n157839),
	.a(n249918),
	.b(n249917));
   in01f01 U268764 (.o(n252878),
	.a(regtop_g_wd_r[11]));
   ao12s01 U268765 (.o(n249919),
	.a(n252269),
	.b(n252270),
	.c(regtop_g_wd_r[11]));
   na02s01 U268766 (.o(n249920),
	.a(regtop_g_isdc_r),
	.b(n249919));
   oa12s01 U268767 (.o(n162088),
	.a(n249920),
	.b(n252273),
	.c(n252878));
   in01s01 U268768 (.o(n249921),
	.a(busrtop_b_rreq_vrh_cnt_18byte_r[1]));
   in01s01 U268769 (.o(n249922),
	.a(busrtop_b_rreq_vrh_cnt_18byte_r[0]));
   na02s01 U268770 (.o(n249923),
	.a(busiftop_status_b_current_0_),
	.b(n249921));
   oa22s01 U268771 (.o(n170932),
	.a(busiftop_status_b_current_0_),
	.b(n249921),
	.c(n249922),
	.d(n249923));
   ao22s01 U268772 (.o(n170937),
	.a(busrtop_b_rreq_vrh_cnt_18byte_r[0]),
	.b(busiftop_status_b_current_0_),
	.c(n249923),
	.d(n249922));
   ao12m01 U268773 (.o(n249931),
	.a(n249944),
	.b(regtop_g_embv_adr_r[6]),
	.c(n249945));
   ao12m01 U268774 (.o(n249932),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embv_adr_r[5]));
   ao12m01 U268775 (.o(n249933),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embv_adr_r[4]));
   ao12m01 U268776 (.o(n249934),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embv_adr_r[3]));
   ao12m01 U268777 (.o(n249935),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embv_adr_r[2]));
   ao12m01 U268778 (.o(n249936),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embv_adr_r[1]));
   ao12m01 U268779 (.o(n249937),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embv_adr_r[0]));
   ao12f01 U268780 (.o(n249938),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embh_adr_r[6]));
   ao12m01 U268781 (.o(n249939),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embh_adr_r[5]));
   ao12m01 U268782 (.o(n249940),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embh_adr_r[4]));
   ao12m01 U268783 (.o(n249941),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embh_adr_r[3]));
   ao12m01 U268784 (.o(n249942),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embh_adr_r[2]));
   ao12m01 U268785 (.o(n249943),
	.a(n249944),
	.b(n249945),
	.c(regtop_g_embh_adr_r[1]));
   in01s01 U268786 (.o(n184630),
	.a(n249949));
   in01s01 U268787 (.o(n184631),
	.a(n249950));
   in01s01 U268788 (.o(n184632),
	.a(n249951));
   in01s01 U268789 (.o(n184633),
	.a(n249952));
   in01s01 U268790 (.o(n184634),
	.a(n249953));
   oa22s01 U268791 (.o(n249954),
	.a(n249982),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[506]),
	.d(FE_OFN268_n249964));
   in01s01 U268792 (.o(n184636),
	.a(n249955));
   in01s01 U268793 (.o(n184637),
	.a(n249956));
   in01s01 U268794 (.o(n184638),
	.a(n249957));
   in01s01 U268795 (.o(n184639),
	.a(n249958));
   in01s01 U268796 (.o(n184640),
	.a(n249959));
   in01s01 U268797 (.o(n184641),
	.a(n249960));
   in01s01 U268798 (.o(n184642),
	.a(n249961));
   in01s01 U268799 (.o(n184643),
	.a(n249962));
   in01s01 U268800 (.o(n184644),
	.a(n249963));
   in01s01 U268801 (.o(n184645),
	.a(n249965));
   in01s01 U268802 (.o(n184646),
	.a(n249966));
   in01s01 U268803 (.o(n184647),
	.a(n249967));
   in01s01 U268804 (.o(n184648),
	.a(n249968));
   in01s01 U268805 (.o(n184649),
	.a(n249969));
   oa22s01 U268806 (.o(n249970),
	.a(n249982),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[491]),
	.d(FE_OFN268_n249964));
   in01s01 U268807 (.o(n184651),
	.a(n249971));
   in01s01 U268808 (.o(n184652),
	.a(n249972));
   in01s01 U268809 (.o(n184653),
	.a(n249973));
   in01s01 U268810 (.o(n184654),
	.a(n249974));
   in01s01 U268811 (.o(n184655),
	.a(n249976));
   oa22s01 U268812 (.o(n249977),
	.a(n249982),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[485]),
	.d(FE_OFN268_n249964));
   in01s01 U268813 (.o(n184656),
	.a(n249977));
   oa22s01 U268814 (.o(n249978),
	.a(n249982),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[484]),
	.d(FE_OFN268_n249964));
   in01s01 U268815 (.o(n184657),
	.a(n249978));
   oa22s01 U268816 (.o(n249979),
	.a(n249982),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[483]),
	.d(FE_OFN268_n249964));
   in01s01 U268817 (.o(n184658),
	.a(n249979));
   oa22s01 U268818 (.o(n249980),
	.a(n249982),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[482]),
	.d(FE_OFN268_n249964));
   in01s01 U268819 (.o(n184659),
	.a(n249980));
   oa22s01 U268820 (.o(n249981),
	.a(n249982),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[481]),
	.d(FE_OFN268_n249964));
   in01s01 U268821 (.o(n184660),
	.a(n249981));
   oa22s01 U268822 (.o(n249983),
	.a(n249982),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[480]),
	.d(FE_OFN268_n249964));
   in01s01 U268823 (.o(n184661),
	.a(n249983));
   in01s01 U268824 (.o(n184662),
	.a(n249984));
   in01s01 U268825 (.o(n184663),
	.a(n249985));
   in01s01 U268826 (.o(n184664),
	.a(n249986));
   oa22s01 U268827 (.o(n249987),
	.a(n250018),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[476]),
	.d(FE_OFN402_n249999));
   in01s01 U268828 (.o(n184666),
	.a(n249988));
   in01s01 U268829 (.o(n184667),
	.a(n249989));
   in01s01 U268830 (.o(n184668),
	.a(n249990));
   in01s01 U268831 (.o(n184669),
	.a(n249991));
   in01s01 U268832 (.o(n184670),
	.a(n249992));
   in01s01 U268833 (.o(n184671),
	.a(n249993));
   in01s01 U268834 (.o(n184672),
	.a(n249994));
   in01s01 U268835 (.o(n184673),
	.a(n249995));
   in01s01 U268836 (.o(n184674),
	.a(n249996));
   in01s01 U268837 (.o(n184675),
	.a(n249997));
   in01s01 U268838 (.o(n184676),
	.a(n249998));
   in01s01 U268839 (.o(n184677),
	.a(n250000));
   in01s01 U268840 (.o(n184678),
	.a(n250001));
   in01s01 U268841 (.o(n184679),
	.a(n250002));
   oa22s01 U268842 (.o(n250003),
	.a(n250018),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[461]),
	.d(n249999));
   in01s01 U268843 (.o(n184681),
	.a(n250004));
   in01s01 U268844 (.o(n184682),
	.a(n250005));
   in01s01 U268845 (.o(n184683),
	.a(n250006));
   in01s01 U268846 (.o(n184684),
	.a(n250007));
   in01s01 U268847 (.o(n184685),
	.a(n250008));
   in01s01 U268848 (.o(n184686),
	.a(n250009));
   in01s01 U268849 (.o(n184687),
	.a(n250011));
   oa22s01 U268850 (.o(n250012),
	.a(n250018),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[453]),
	.d(FE_OFN402_n249999));
   in01s01 U268851 (.o(n184688),
	.a(n250012));
   oa22s01 U268852 (.o(n250013),
	.a(n250018),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[452]),
	.d(FE_OFN402_n249999));
   in01s01 U268853 (.o(n184689),
	.a(n250013));
   oa22s01 U268854 (.o(n250014),
	.a(n250018),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[451]),
	.d(FE_OFN402_n249999));
   in01s01 U268855 (.o(n184690),
	.a(n250014));
   oa22s01 U268856 (.o(n250015),
	.a(n250018),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[450]),
	.d(FE_OFN402_n249999));
   in01s01 U268857 (.o(n184691),
	.a(n250015));
   oa22s01 U268858 (.o(n250016),
	.a(n250018),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[449]),
	.d(FE_OFN402_n249999));
   in01s01 U268859 (.o(n184692),
	.a(n250016));
   oa22s01 U268860 (.o(n250019),
	.a(n250018),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[448]),
	.d(FE_OFN402_n249999));
   in01s01 U268861 (.o(n184693),
	.a(n250019));
   in01s01 U268862 (.o(n184694),
	.a(n250020));
   oa22s01 U268863 (.o(n250021),
	.a(n250053),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[446]),
	.d(FE_OFN270_n250035));
   in01s01 U268864 (.o(n184696),
	.a(n250022));
   in01s01 U268865 (.o(n184697),
	.a(n250023));
   in01s01 U268866 (.o(n184698),
	.a(n250024));
   in01s01 U268867 (.o(n184699),
	.a(n250025));
   in01s01 U268868 (.o(n184700),
	.a(n250026));
   in01s01 U268869 (.o(n184701),
	.a(n250027));
   in01s01 U268870 (.o(n184702),
	.a(n250028));
   in01s01 U268871 (.o(n184703),
	.a(n250029));
   in01s01 U268872 (.o(n184704),
	.a(n250030));
   in01s01 U268873 (.o(n184705),
	.a(n250031));
   in01s01 U268874 (.o(n184706),
	.a(n250032));
   in01s01 U268875 (.o(n184707),
	.a(n250033));
   in01s01 U268876 (.o(n184708),
	.a(n250034));
   in01s01 U268877 (.o(n184709),
	.a(n250036));
   oa22s01 U268878 (.o(n250037),
	.a(n250053),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[431]),
	.d(FE_OFN270_n250035));
   in01s01 U268879 (.o(n184711),
	.a(n250038));
   in01s01 U268880 (.o(n184712),
	.a(n250039));
   in01s01 U268881 (.o(n184713),
	.a(n250040));
   in01s01 U268882 (.o(n184714),
	.a(n250041));
   in01s01 U268883 (.o(n184715),
	.a(n250042));
   in01s01 U268884 (.o(n184716),
	.a(n250043));
   in01s01 U268885 (.o(n184717),
	.a(n250044));
   in01s01 U268886 (.o(n184718),
	.a(n250045));
   in01s01 U268887 (.o(n184719),
	.a(n250047));
   oa22s01 U268888 (.o(n250048),
	.a(n250053),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[421]),
	.d(FE_OFN270_n250035));
   in01s01 U268889 (.o(n184720),
	.a(n250048));
   oa22s01 U268890 (.o(n250049),
	.a(n250053),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[420]),
	.d(FE_OFN270_n250035));
   in01s01 U268891 (.o(n184721),
	.a(n250049));
   oa22s01 U268892 (.o(n250050),
	.a(n250053),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[419]),
	.d(FE_OFN270_n250035));
   in01s01 U268893 (.o(n184722),
	.a(n250050));
   oa22s01 U268894 (.o(n250051),
	.a(n250053),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[418]),
	.d(FE_OFN270_n250035));
   in01s01 U268895 (.o(n184723),
	.a(n250051));
   oa22s01 U268896 (.o(n250052),
	.a(n250053),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[417]),
	.d(FE_OFN270_n250035));
   in01s01 U268897 (.o(n184724),
	.a(n250052));
   oa22s01 U268898 (.o(n250054),
	.a(n250053),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[416]),
	.d(FE_OFN270_n250035));
   in01s01 U268899 (.o(n184726),
	.a(n250056));
   in01s01 U268900 (.o(n184727),
	.a(n250057));
   in01s01 U268901 (.o(n184728),
	.a(n250058));
   in01s01 U268902 (.o(n184729),
	.a(n250059));
   in01s01 U268903 (.o(n184730),
	.a(n250060));
   in01s01 U268904 (.o(n184731),
	.a(n250061));
   in01s01 U268905 (.o(n184732),
	.a(n250062));
   in01s01 U268906 (.o(n184733),
	.a(n250063));
   in01s01 U268907 (.o(n184734),
	.a(n250064));
   in01s01 U268908 (.o(n184735),
	.a(n250065));
   in01s01 U268909 (.o(n184736),
	.a(n250066));
   in01s01 U268910 (.o(n184737),
	.a(n250067));
   in01s01 U268911 (.o(n184738),
	.a(n250068));
   in01s01 U268912 (.o(n184739),
	.a(n250069));
   oa22s01 U268913 (.o(n250070),
	.a(n250089),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[401]),
	.d(FE_OFN404_n250071));
   in01s01 U268914 (.o(n184741),
	.a(n250072));
   in01s01 U268915 (.o(n184742),
	.a(n250073));
   in01s01 U268916 (.o(n184743),
	.a(n250074));
   in01s01 U268917 (.o(n184744),
	.a(n250075));
   in01s01 U268918 (.o(n184745),
	.a(n250076));
   in01s01 U268919 (.o(n184746),
	.a(n250077));
   in01s01 U268920 (.o(n184747),
	.a(n250078));
   in01s01 U268921 (.o(n184748),
	.a(n250079));
   in01s01 U268922 (.o(n184749),
	.a(n250080));
   in01s01 U268923 (.o(n184750),
	.a(n250081));
   in01s01 U268924 (.o(n184751),
	.a(n250083));
   oa22s01 U268925 (.o(n250084),
	.a(n250089),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[389]),
	.d(FE_OFN404_n250071));
   in01s01 U268926 (.o(n184752),
	.a(n250084));
   oa22s01 U268927 (.o(n250085),
	.a(n250089),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[388]),
	.d(FE_OFN404_n250071));
   in01s01 U268928 (.o(n184753),
	.a(n250085));
   oa22s01 U268929 (.o(n250086),
	.a(n250089),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[387]),
	.d(FE_OFN404_n250071));
   in01s01 U268930 (.o(n184754),
	.a(n250086));
   oa22s01 U268931 (.o(n250087),
	.a(n250089),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[386]),
	.d(FE_OFN404_n250071));
   oa22s01 U268932 (.o(n250088),
	.a(n250089),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[385]),
	.d(FE_OFN404_n250071));
   in01s01 U268933 (.o(n184756),
	.a(n250088));
   oa22s01 U268934 (.o(n250090),
	.a(n250089),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[384]),
	.d(FE_OFN404_n250071));
   in01s01 U268935 (.o(n184757),
	.a(n250090));
   in01s01 U268936 (.o(n184758),
	.a(n250092));
   in01s01 U268937 (.o(n184759),
	.a(n250093));
   in01s01 U268938 (.o(n184760),
	.a(n250094));
   in01s01 U268939 (.o(n184761),
	.a(n250095));
   in01s01 U268940 (.o(n184762),
	.a(n250096));
   in01s01 U268941 (.o(n184763),
	.a(n250097));
   in01s01 U268942 (.o(n184764),
	.a(n250098));
   in01s01 U268943 (.o(n184765),
	.a(n250099));
   in01s01 U268944 (.o(n184766),
	.a(n250100));
   in01s01 U268945 (.o(n184767),
	.a(n250101));
   in01s01 U268946 (.o(n184768),
	.a(n250102));
   in01s01 U268947 (.o(n184769),
	.a(n250103));
   oa22s01 U268948 (.o(n250104),
	.a(n250126),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[371]),
	.d(FE_OFN193_n250107));
   in01s01 U268949 (.o(n184771),
	.a(n250105));
   in01s01 U268950 (.o(n184772),
	.a(n250106));
   in01s01 U268951 (.o(n184773),
	.a(n250108));
   in01s01 U268952 (.o(n184774),
	.a(n250109));
   in01s01 U268953 (.o(n184775),
	.a(n250110));
   in01s01 U268954 (.o(n184776),
	.a(n250111));
   in01s01 U268955 (.o(n184777),
	.a(n250112));
   in01s01 U268956 (.o(n184778),
	.a(n250113));
   in01s01 U268957 (.o(n184779),
	.a(n250114));
   in01s01 U268958 (.o(n184780),
	.a(n250115));
   in01s01 U268959 (.o(n184781),
	.a(n250116));
   in01s01 U268960 (.o(n184782),
	.a(n250117));
   in01s01 U268961 (.o(n184783),
	.a(n250119));
   oa22s01 U268962 (.o(n250120),
	.a(n250126),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[357]),
	.d(FE_OFN193_n250107));
   in01s01 U268963 (.o(n184784),
	.a(n250120));
   oa22s01 U268964 (.o(n250121),
	.a(n250126),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[356]),
	.d(FE_OFN193_n250107));
   oa22s01 U268965 (.o(n250122),
	.a(n250126),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[355]),
	.d(FE_OFN193_n250107));
   in01s01 U268966 (.o(n184786),
	.a(n250122));
   oa22s01 U268967 (.o(n250123),
	.a(n250126),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[354]),
	.d(FE_OFN193_n250107));
   in01s01 U268968 (.o(n184787),
	.a(n250123));
   oa22s01 U268969 (.o(n250124),
	.a(n250126),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[353]),
	.d(FE_OFN193_n250107));
   in01s01 U268970 (.o(n184788),
	.a(n250124));
   oa22s01 U268971 (.o(n250127),
	.a(n250126),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[352]),
	.d(FE_OFN192_n250107));
   in01s01 U268972 (.o(n184789),
	.a(n250127));
   oa22s01 U268973 (.o(n250129),
	.a(FE_OFN406_n250162),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[351]),
	.d(FE_OFN272_n250144));
   in01s01 U268974 (.o(n184790),
	.a(n250129));
   oa22s01 U268975 (.o(n250130),
	.a(n250162),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[350]),
	.d(FE_OFN272_n250144));
   in01s01 U268976 (.o(n184791),
	.a(n250130));
   oa22s01 U268977 (.o(n250131),
	.a(n250162),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[349]),
	.d(n250144));
   in01s01 U268978 (.o(n184792),
	.a(n250131));
   oa22s01 U268979 (.o(n250132),
	.a(n250162),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[348]),
	.d(n250144));
   in01s01 U268980 (.o(n184793),
	.a(n250132));
   oa22s01 U268981 (.o(n250133),
	.a(n250162),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[347]),
	.d(n250144));
   in01s01 U268982 (.o(n184794),
	.a(n250133));
   in01s01 U268983 (.o(n184795),
	.a(n250134));
   oa22s01 U268984 (.o(n250135),
	.a(n250162),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[345]),
	.d(FE_OFN272_n250144));
   in01s01 U268985 (.o(n184796),
	.a(n250135));
   in01s01 U268986 (.o(n184797),
	.a(n250136));
   oa22s01 U268987 (.o(n250137),
	.a(n250162),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[343]),
	.d(FE_OFN272_n250144));
   in01s01 U268988 (.o(n184798),
	.a(n250137));
   in01s01 U268989 (.o(n184799),
	.a(n250138));
   oa22s01 U268990 (.o(n250139),
	.a(n250162),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[341]),
	.d(FE_OFN272_n250144));
   in01s01 U268991 (.o(n184801),
	.a(n250140));
   oa22s01 U268992 (.o(n250141),
	.a(n250162),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[339]),
	.d(FE_OFN272_n250144));
   in01s01 U268993 (.o(n184802),
	.a(n250141));
   in01s01 U268994 (.o(n184803),
	.a(n250142));
   oa22s01 U268995 (.o(n250143),
	.a(FE_OFN406_n250162),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[337]),
	.d(FE_OFN272_n250144));
   in01s01 U268996 (.o(n184804),
	.a(n250143));
   oa22s01 U268997 (.o(n250145),
	.a(FE_OFN406_n250162),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[336]),
	.d(FE_OFN272_n250144));
   in01s01 U268998 (.o(n184805),
	.a(n250145));
   in01s01 U268999 (.o(n184806),
	.a(n250146));
   in01s01 U269000 (.o(n184807),
	.a(n250147));
   oa22s01 U269001 (.o(n250148),
	.a(n250162),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[333]),
	.d(n250144));
   in01s01 U269002 (.o(n184808),
	.a(n250148));
   oa22s01 U269003 (.o(n250149),
	.a(FE_OFN406_n250162),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[332]),
	.d(FE_OFN272_n250144));
   in01s01 U269004 (.o(n184809),
	.a(n250149));
   oa22s01 U269005 (.o(n250150),
	.a(FE_OFN406_n250162),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[331]),
	.d(FE_OFN272_n250144));
   in01s01 U269006 (.o(n184810),
	.a(n250150));
   oa22s01 U269007 (.o(n250151),
	.a(n250162),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[330]),
	.d(n250144));
   in01s01 U269008 (.o(n184811),
	.a(n250151));
   oa22s01 U269009 (.o(n250152),
	.a(n250162),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[329]),
	.d(FE_OFN272_n250144));
   in01s01 U269010 (.o(n184812),
	.a(n250152));
   in01s01 U269011 (.o(n184813),
	.a(n250153));
   in01s01 U269012 (.o(n184814),
	.a(n250154));
   oa22s01 U269013 (.o(n250156),
	.a(n250162),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[326]),
	.d(n250144));
   oa22s01 U269014 (.o(n250157),
	.a(FE_OFN406_n250162),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[325]),
	.d(FE_OFN272_n250144));
   in01s01 U269015 (.o(n184816),
	.a(n250157));
   oa22s01 U269016 (.o(n250158),
	.a(FE_OFN406_n250162),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[324]),
	.d(FE_OFN272_n250144));
   in01s01 U269017 (.o(n184817),
	.a(n250158));
   oa22s01 U269018 (.o(n250159),
	.a(FE_OFN406_n250162),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[323]),
	.d(FE_OFN272_n250144));
   in01s01 U269019 (.o(n184818),
	.a(n250159));
   oa22s01 U269020 (.o(n250160),
	.a(n250162),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[322]),
	.d(FE_OFN272_n250144));
   in01s01 U269021 (.o(n184819),
	.a(n250160));
   oa22s01 U269022 (.o(n250161),
	.a(FE_OFN406_n250162),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[321]),
	.d(FE_OFN272_n250144));
   in01s01 U269023 (.o(n184820),
	.a(n250161));
   oa22s01 U269024 (.o(n250163),
	.a(n250162),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[320]),
	.d(FE_OFN272_n250144));
   in01s01 U269025 (.o(n184821),
	.a(n250163));
   in01s01 U269026 (.o(n184822),
	.a(n250165));
   in01s01 U269027 (.o(n184823),
	.a(n250166));
   in01s01 U269028 (.o(n184824),
	.a(n250167));
   in01s01 U269029 (.o(n184825),
	.a(n250168));
   in01s01 U269030 (.o(n184826),
	.a(n250169));
   in01s01 U269031 (.o(n184827),
	.a(n250170));
   in01s01 U269032 (.o(n184828),
	.a(n250171));
   in01s01 U269033 (.o(n184829),
	.a(n250172));
   oa22s01 U269034 (.o(n250173),
	.a(n250198),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[311]),
	.d(FE_OFN274_n250180));
   in01s01 U269035 (.o(n184831),
	.a(n250174));
   in01s01 U269036 (.o(n184832),
	.a(n250175));
   in01s01 U269037 (.o(n184833),
	.a(n250176));
   in01s01 U269038 (.o(n184834),
	.a(n250177));
   in01s01 U269039 (.o(n184835),
	.a(n250178));
   in01s01 U269040 (.o(n184836),
	.a(n250179));
   in01s01 U269041 (.o(n184837),
	.a(n250181));
   in01s01 U269042 (.o(n184838),
	.a(n250182));
   in01s01 U269043 (.o(n184839),
	.a(n250183));
   in01s01 U269044 (.o(n184840),
	.a(n250184));
   in01s01 U269045 (.o(n184841),
	.a(n250185));
   in01s01 U269046 (.o(n184842),
	.a(n250186));
   in01s01 U269047 (.o(n184843),
	.a(n250187));
   in01s01 U269048 (.o(n184844),
	.a(n250188));
   oa22s01 U269049 (.o(n250189),
	.a(n250198),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[296]),
	.d(FE_OFN274_n250180));
   in01s01 U269050 (.o(n184846),
	.a(n250190));
   in01s01 U269051 (.o(n184847),
	.a(n250192));
   oa22s01 U269052 (.o(n250193),
	.a(n250198),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[293]),
	.d(FE_OFN274_n250180));
   in01s01 U269053 (.o(n184848),
	.a(n250193));
   oa22s01 U269054 (.o(n250194),
	.a(n250198),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[292]),
	.d(FE_OFN274_n250180));
   in01s01 U269055 (.o(n184849),
	.a(n250194));
   oa22s01 U269056 (.o(n250195),
	.a(n250198),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[291]),
	.d(FE_OFN274_n250180));
   in01s01 U269057 (.o(n184850),
	.a(n250195));
   oa22s01 U269058 (.o(n250196),
	.a(n250198),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[290]),
	.d(FE_OFN274_n250180));
   in01s01 U269059 (.o(n184851),
	.a(n250196));
   oa22s01 U269060 (.o(n250197),
	.a(n250198),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[289]),
	.d(FE_OFN274_n250180));
   in01s01 U269061 (.o(n184852),
	.a(n250197));
   oa22s01 U269062 (.o(n250199),
	.a(n250198),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[288]),
	.d(FE_OFN274_n250180));
   in01s01 U269063 (.o(n184853),
	.a(n250199));
   oa22s01 U269064 (.o(n250203),
	.a(n250237),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[287]),
	.d(FE_OFN276_n250218));
   in01s01 U269065 (.o(n184854),
	.a(n250203));
   oa22s01 U269066 (.o(n250204),
	.a(n250237),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[286]),
	.d(FE_OFN276_n250218));
   in01s01 U269067 (.o(n184855),
	.a(n250204));
   oa22s01 U269068 (.o(n250205),
	.a(n250237),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[285]),
	.d(FE_OFN276_n250218));
   in01s01 U269069 (.o(n184856),
	.a(n250205));
   oa22s01 U269070 (.o(n250206),
	.a(n250237),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[284]),
	.d(FE_OFN276_n250218));
   in01s01 U269071 (.o(n184857),
	.a(n250206));
   oa22s01 U269072 (.o(n250207),
	.a(n250237),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[283]),
	.d(FE_OFN276_n250218));
   in01s01 U269073 (.o(n184858),
	.a(n250207));
   oa22s01 U269074 (.o(n250208),
	.a(n250237),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[282]),
	.d(FE_OFN276_n250218));
   in01s01 U269075 (.o(n184859),
	.a(n250208));
   oa22s01 U269076 (.o(n250209),
	.a(n250237),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[281]),
	.d(FE_OFN276_n250218));
   oa22s01 U269077 (.o(n250210),
	.a(n250237),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[280]),
	.d(FE_OFN276_n250218));
   in01s01 U269078 (.o(n184861),
	.a(n250210));
   oa22s01 U269079 (.o(n250211),
	.a(n250237),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[279]),
	.d(FE_OFN276_n250218));
   in01s01 U269080 (.o(n184862),
	.a(n250211));
   oa22s01 U269081 (.o(n250212),
	.a(n250237),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[278]),
	.d(FE_OFN276_n250218));
   in01s01 U269082 (.o(n184863),
	.a(n250212));
   oa22s01 U269083 (.o(n250213),
	.a(n250237),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[277]),
	.d(FE_OFN276_n250218));
   in01s01 U269084 (.o(n184864),
	.a(n250213));
   oa22s01 U269085 (.o(n250214),
	.a(n250237),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[276]),
	.d(FE_OFN276_n250218));
   in01s01 U269086 (.o(n184865),
	.a(n250214));
   oa22s01 U269087 (.o(n250215),
	.a(n250237),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[275]),
	.d(FE_OFN276_n250218));
   in01s01 U269088 (.o(n184866),
	.a(n250215));
   oa22s01 U269089 (.o(n250216),
	.a(n250237),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[274]),
	.d(FE_OFN276_n250218));
   in01s01 U269090 (.o(n184867),
	.a(n250216));
   oa22s01 U269091 (.o(n250217),
	.a(n250237),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[273]),
	.d(FE_OFN276_n250218));
   in01s01 U269092 (.o(n184868),
	.a(n250217));
   oa22s01 U269093 (.o(n250219),
	.a(n250237),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[272]),
	.d(FE_OFN276_n250218));
   in01s01 U269094 (.o(n184869),
	.a(n250219));
   oa22s01 U269095 (.o(n250220),
	.a(n250237),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[271]),
	.d(FE_OFN276_n250218));
   in01s01 U269096 (.o(n184870),
	.a(n250220));
   oa22s01 U269097 (.o(n250221),
	.a(n250237),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[270]),
	.d(FE_OFN276_n250218));
   in01s01 U269098 (.o(n184871),
	.a(n250221));
   oa22s01 U269099 (.o(n250222),
	.a(n250237),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[269]),
	.d(FE_OFN276_n250218));
   in01s01 U269100 (.o(n184872),
	.a(n250222));
   oa22s01 U269101 (.o(n250223),
	.a(n250237),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[268]),
	.d(FE_OFN276_n250218));
   in01s01 U269102 (.o(n184873),
	.a(n250223));
   oa22s01 U269103 (.o(n250224),
	.a(n250237),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[267]),
	.d(FE_OFN276_n250218));
   in01s01 U269104 (.o(n184874),
	.a(n250224));
   oa22s01 U269105 (.o(n250225),
	.a(n250237),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[266]),
	.d(FE_OFN276_n250218));
   oa22s01 U269106 (.o(n250226),
	.a(n250237),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[265]),
	.d(FE_OFN276_n250218));
   in01s01 U269107 (.o(n184876),
	.a(n250226));
   oa22s01 U269108 (.o(n250227),
	.a(n250237),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[264]),
	.d(FE_OFN276_n250218));
   in01s01 U269109 (.o(n184877),
	.a(n250227));
   oa22s01 U269110 (.o(n250228),
	.a(n250237),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[263]),
	.d(FE_OFN276_n250218));
   in01s01 U269111 (.o(n184878),
	.a(n250228));
   oa22s01 U269112 (.o(n250230),
	.a(n250237),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[262]),
	.d(FE_OFN276_n250218));
   in01s01 U269113 (.o(n184879),
	.a(n250230));
   oa22s01 U269114 (.o(n250231),
	.a(n250237),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[261]),
	.d(FE_OFN276_n250218));
   in01s01 U269115 (.o(n184880),
	.a(n250231));
   oa22s01 U269116 (.o(n250232),
	.a(n250237),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[260]),
	.d(FE_OFN276_n250218));
   in01s01 U269117 (.o(n184881),
	.a(n250232));
   oa22s01 U269118 (.o(n250233),
	.a(n250237),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[259]),
	.d(FE_OFN276_n250218));
   in01s01 U269119 (.o(n184882),
	.a(n250233));
   oa22s01 U269120 (.o(n250234),
	.a(n250237),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[258]),
	.d(FE_OFN276_n250218));
   in01s01 U269121 (.o(n184883),
	.a(n250234));
   oa22s01 U269122 (.o(n250235),
	.a(n250237),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[257]),
	.d(FE_OFN276_n250218));
   in01s01 U269123 (.o(n184884),
	.a(n250235));
   oa22s01 U269124 (.o(n250238),
	.a(n250237),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[256]),
	.d(FE_OFN276_n250218));
   in01s01 U269125 (.o(n184885),
	.a(n250238));
   in01s01 U269126 (.o(n184886),
	.a(n250239));
   in01s01 U269127 (.o(n184887),
	.a(n250240));
   in01s01 U269128 (.o(n184888),
	.a(n250241));
   in01s01 U269129 (.o(n184889),
	.a(n250242));
   oa22s01 U269130 (.o(n250243),
	.a(n250272),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[251]),
	.d(FE_OFN278_n250254));
   in01s01 U269131 (.o(n184891),
	.a(n250244));
   in01s01 U269132 (.o(n184892),
	.a(n250245));
   in01s01 U269133 (.o(n184893),
	.a(n250246));
   in01s01 U269134 (.o(n184894),
	.a(n250247));
   in01s01 U269135 (.o(n184895),
	.a(n250248));
   in01s01 U269136 (.o(n184896),
	.a(n250249));
   in01s01 U269137 (.o(n184897),
	.a(n250250));
   in01s01 U269138 (.o(n184898),
	.a(n250251));
   in01s01 U269139 (.o(n184899),
	.a(n250252));
   in01s01 U269140 (.o(n184900),
	.a(n250253));
   in01s01 U269141 (.o(n184901),
	.a(n250255));
   in01s01 U269142 (.o(n184902),
	.a(n250256));
   in01s01 U269143 (.o(n184903),
	.a(n250257));
   in01s01 U269144 (.o(n184904),
	.a(n250258));
   oa22s01 U269145 (.o(n250259),
	.a(n250272),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[236]),
	.d(FE_OFN278_n250254));
   in01s01 U269146 (.o(n184906),
	.a(n250260));
   in01s01 U269147 (.o(n184907),
	.a(n250261));
   in01s01 U269148 (.o(n184908),
	.a(n250262));
   in01s01 U269149 (.o(n184909),
	.a(n250263));
   in01s01 U269150 (.o(n184910),
	.a(n250264));
   in01s01 U269151 (.o(n184911),
	.a(n250266));
   oa22s01 U269152 (.o(n250267),
	.a(n250272),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[229]),
	.d(FE_OFN278_n250254));
   in01s01 U269153 (.o(n184912),
	.a(n250267));
   oa22s01 U269154 (.o(n250268),
	.a(n250272),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[228]),
	.d(FE_OFN278_n250254));
   in01s01 U269155 (.o(n184913),
	.a(n250268));
   oa22s01 U269156 (.o(n250269),
	.a(n250272),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[227]),
	.d(FE_OFN278_n250254));
   in01s01 U269157 (.o(n184914),
	.a(n250269));
   oa22s01 U269158 (.o(n250270),
	.a(n250272),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[226]),
	.d(FE_OFN278_n250254));
   in01s01 U269159 (.o(n184915),
	.a(n250270));
   oa22s01 U269160 (.o(n250271),
	.a(n250272),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[225]),
	.d(FE_OFN278_n250254));
   in01s01 U269161 (.o(n184916),
	.a(n250271));
   oa22s01 U269162 (.o(n250273),
	.a(n250272),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[224]),
	.d(FE_OFN278_n250254));
   in01s01 U269163 (.o(n184917),
	.a(n250273));
   in01s01 U269164 (.o(n184918),
	.a(n250274));
   in01s01 U269165 (.o(n184919),
	.a(n250275));
   oa22s01 U269166 (.o(n250276),
	.a(n250307),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[221]),
	.d(FE_OFN408_n250289));
   in01s01 U269167 (.o(n184921),
	.a(n250277));
   in01s01 U269168 (.o(n184922),
	.a(n250278));
   in01s01 U269169 (.o(n184923),
	.a(n250279));
   in01s01 U269170 (.o(n184924),
	.a(n250280));
   in01s01 U269171 (.o(n184925),
	.a(n250281));
   in01s01 U269172 (.o(n184926),
	.a(n250282));
   in01s01 U269173 (.o(n184927),
	.a(n250283));
   in01s01 U269174 (.o(n184928),
	.a(n250284));
   in01s01 U269175 (.o(n184929),
	.a(n250285));
   in01s01 U269176 (.o(n184930),
	.a(n250286));
   in01s01 U269177 (.o(n184931),
	.a(n250287));
   in01s01 U269178 (.o(n184932),
	.a(n250288));
   in01s01 U269179 (.o(n184933),
	.a(n250290));
   in01s01 U269180 (.o(n184934),
	.a(n250291));
   oa22s01 U269181 (.o(n250292),
	.a(n250307),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[206]),
	.d(FE_OFN408_n250289));
   in01s01 U269182 (.o(n184936),
	.a(n250293));
   in01s01 U269183 (.o(n184937),
	.a(n250294));
   in01s01 U269184 (.o(n184938),
	.a(n250295));
   in01s01 U269185 (.o(n184939),
	.a(n250296));
   in01s01 U269186 (.o(n184940),
	.a(n250297));
   in01s01 U269187 (.o(n184941),
	.a(n250298));
   in01s01 U269188 (.o(n184942),
	.a(n250299));
   in01s01 U269189 (.o(n184943),
	.a(n250301));
   oa22s01 U269190 (.o(n250302),
	.a(n250307),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[197]),
	.d(FE_OFN408_n250289));
   in01s01 U269191 (.o(n184944),
	.a(n250302));
   oa22s01 U269192 (.o(n250303),
	.a(n250307),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[196]),
	.d(FE_OFN408_n250289));
   in01s01 U269193 (.o(n184945),
	.a(n250303));
   oa22s01 U269194 (.o(n250304),
	.a(n250307),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[195]),
	.d(FE_OFN408_n250289));
   in01s01 U269195 (.o(n184946),
	.a(n250304));
   oa22s01 U269196 (.o(n250305),
	.a(n250307),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[194]),
	.d(FE_OFN408_n250289));
   in01s01 U269197 (.o(n184947),
	.a(n250305));
   oa22s01 U269198 (.o(n250306),
	.a(n250307),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[193]),
	.d(FE_OFN408_n250289));
   in01s01 U269199 (.o(n184948),
	.a(n250306));
   oa22s01 U269200 (.o(n250308),
	.a(n250307),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[192]),
	.d(FE_OFN408_n250289));
   in01s01 U269201 (.o(n184949),
	.a(n250308));
   oa22s01 U269202 (.o(n250309),
	.a(n250343),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[191]),
	.d(FE_OFN280_n250324));
   in01s01 U269203 (.o(n184951),
	.a(n250310));
   in01s01 U269204 (.o(n184952),
	.a(n250311));
   in01s01 U269205 (.o(n184953),
	.a(n250312));
   in01s01 U269206 (.o(n184954),
	.a(n250313));
   in01s01 U269207 (.o(n184955),
	.a(n250314));
   in01s01 U269208 (.o(n184956),
	.a(n250315));
   in01s01 U269209 (.o(n184957),
	.a(n250316));
   in01s01 U269210 (.o(n184958),
	.a(n250317));
   in01s01 U269211 (.o(n184959),
	.a(n250318));
   in01s01 U269212 (.o(n184960),
	.a(n250319));
   in01s01 U269213 (.o(n184961),
	.a(n250320));
   in01s01 U269214 (.o(n184962),
	.a(n250321));
   in01s01 U269215 (.o(n184963),
	.a(n250322));
   in01s01 U269216 (.o(n184964),
	.a(n250323));
   oa22s01 U269217 (.o(n250325),
	.a(n250343),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[176]),
	.d(FE_OFN280_n250324));
   in01s01 U269218 (.o(n184966),
	.a(n250326));
   in01s01 U269219 (.o(n184967),
	.a(n250327));
   in01s01 U269220 (.o(n184968),
	.a(n250328));
   in01s01 U269221 (.o(n184969),
	.a(n250329));
   in01s01 U269222 (.o(n184970),
	.a(n250330));
   in01s01 U269223 (.o(n184971),
	.a(n250331));
   in01s01 U269224 (.o(n184972),
	.a(n250332));
   in01s01 U269225 (.o(n184973),
	.a(n250333));
   in01s01 U269226 (.o(n184974),
	.a(n250334));
   in01s01 U269227 (.o(n184975),
	.a(n250336));
   oa22s01 U269228 (.o(n250337),
	.a(n250343),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[165]),
	.d(FE_OFN280_n250324));
   in01s01 U269229 (.o(n184976),
	.a(n250337));
   oa22s01 U269230 (.o(n250338),
	.a(n250343),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[164]),
	.d(FE_OFN280_n250324));
   in01s01 U269231 (.o(n184977),
	.a(n250338));
   oa22s01 U269232 (.o(n250339),
	.a(n250343),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[163]),
	.d(FE_OFN280_n250324));
   in01s01 U269233 (.o(n184978),
	.a(n250339));
   oa22s01 U269234 (.o(n250340),
	.a(n250343),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[162]),
	.d(FE_OFN280_n250324));
   in01s01 U269235 (.o(n184979),
	.a(n250340));
   oa22s01 U269236 (.o(n250341),
	.a(n250343),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[161]),
	.d(FE_OFN280_n250324));
   oa22s01 U269237 (.o(n250344),
	.a(n250343),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[160]),
	.d(FE_OFN280_n250324));
   in01s01 U269238 (.o(n184981),
	.a(n250344));
   in01s01 U269239 (.o(n184982),
	.a(n250345));
   in01s01 U269240 (.o(n184983),
	.a(n250346));
   in01s01 U269241 (.o(n184984),
	.a(n250347));
   in01s01 U269242 (.o(n184985),
	.a(n250348));
   in01s01 U269243 (.o(n184986),
	.a(n250349));
   in01s01 U269244 (.o(n184987),
	.a(n250350));
   in01s01 U269245 (.o(n184988),
	.a(n250351));
   in01s01 U269246 (.o(n184989),
	.a(n250352));
   in01s01 U269247 (.o(n184990),
	.a(n250353));
   in01s01 U269248 (.o(n184991),
	.a(n250354));
   in01s01 U269249 (.o(n184992),
	.a(n250355));
   in01s01 U269250 (.o(n184993),
	.a(n250356));
   in01s01 U269251 (.o(n184994),
	.a(n250357));
   oa22s01 U269252 (.o(n250358),
	.a(n250378),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[146]),
	.d(FE_OFN410_n250360));
   in01s01 U269253 (.o(n184996),
	.a(n250359));
   in01s01 U269254 (.o(n184997),
	.a(n250361));
   in01s01 U269255 (.o(n184998),
	.a(n250362));
   in01s01 U269256 (.o(n184999),
	.a(n250363));
   in01s01 U269257 (.o(n185000),
	.a(n250364));
   in01s01 U269258 (.o(n185001),
	.a(n250365));
   in01s01 U269259 (.o(n185002),
	.a(n250366));
   in01s01 U269260 (.o(n185003),
	.a(n250367));
   in01s01 U269261 (.o(n185004),
	.a(n250368));
   in01s01 U269262 (.o(n185005),
	.a(n250369));
   in01s01 U269263 (.o(n185006),
	.a(n250370));
   in01s01 U269264 (.o(n185007),
	.a(n250372));
   oa22s01 U269265 (.o(n250373),
	.a(n250378),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[133]),
	.d(FE_OFN410_n250360));
   in01s01 U269266 (.o(n185008),
	.a(n250373));
   oa22s01 U269267 (.o(n250374),
	.a(n250378),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[132]),
	.d(FE_OFN410_n250360));
   in01s01 U269268 (.o(n185009),
	.a(n250374));
   oa22s01 U269269 (.o(n250375),
	.a(n250378),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[131]),
	.d(FE_OFN410_n250360));
   oa22s01 U269270 (.o(n250376),
	.a(n250378),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[130]),
	.d(FE_OFN410_n250360));
   in01s01 U269271 (.o(n185011),
	.a(n250376));
   oa22s01 U269272 (.o(n250377),
	.a(n250378),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[129]),
	.d(FE_OFN410_n250360));
   in01s01 U269273 (.o(n185012),
	.a(n250377));
   oa22s01 U269274 (.o(n250379),
	.a(n250378),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[128]),
	.d(FE_OFN410_n250360));
   in01s01 U269275 (.o(n185013),
	.a(n250379));
   in01s01 U269276 (.o(n185014),
	.a(n250380));
   in01s01 U269277 (.o(n185015),
	.a(n250381));
   in01s01 U269278 (.o(n185016),
	.a(n250382));
   in01s01 U269279 (.o(n185017),
	.a(n250383));
   in01s01 U269280 (.o(n185018),
	.a(n250384));
   in01s01 U269281 (.o(n185019),
	.a(n250385));
   in01s01 U269282 (.o(n185020),
	.a(n250386));
   in01s01 U269283 (.o(n185021),
	.a(n250387));
   in01s01 U269284 (.o(n185022),
	.a(n250388));
   in01s01 U269285 (.o(n185023),
	.a(n250389));
   in01s01 U269286 (.o(n185024),
	.a(n250390));
   oa22s01 U269287 (.o(n250391),
	.a(n250413),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[116]),
	.d(FE_OFN195_n250395));
   in01s01 U269288 (.o(n185026),
	.a(n250392));
   in01s01 U269289 (.o(n185027),
	.a(n250393));
   in01s01 U269290 (.o(n185028),
	.a(n250394));
   in01s01 U269291 (.o(n185029),
	.a(n250396));
   in01s01 U269292 (.o(n185030),
	.a(n250397));
   in01s01 U269293 (.o(n185031),
	.a(n250398));
   in01s01 U269294 (.o(n185032),
	.a(n250399));
   in01s01 U269295 (.o(n185033),
	.a(n250400));
   in01s01 U269296 (.o(n185034),
	.a(n250401));
   in01s01 U269297 (.o(n185035),
	.a(n250402));
   in01s01 U269298 (.o(n185036),
	.a(n250403));
   in01s01 U269299 (.o(n185037),
	.a(n250404));
   in01s01 U269300 (.o(n185038),
	.a(n250405));
   in01s01 U269301 (.o(n185039),
	.a(n250407));
   oa22s01 U269302 (.o(n250408),
	.a(n250413),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[101]),
	.d(FE_OFN195_n250395));
   oa22s01 U269303 (.o(n250409),
	.a(n250413),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[100]),
	.d(FE_OFN195_n250395));
   in01s01 U269304 (.o(n185041),
	.a(n250409));
   oa22s01 U269305 (.o(n250410),
	.a(n250413),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[99]),
	.d(FE_OFN195_n250395));
   in01s01 U269306 (.o(n185042),
	.a(n250410));
   oa22s01 U269307 (.o(n250411),
	.a(n250413),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[98]),
	.d(FE_OFN195_n250395));
   in01s01 U269308 (.o(n185043),
	.a(n250411));
   oa22s01 U269309 (.o(n250412),
	.a(n250413),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[97]),
	.d(FE_OFN195_n250395));
   in01s01 U269310 (.o(n185044),
	.a(n250412));
   oa22s01 U269311 (.o(n250414),
	.a(n250413),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[96]),
	.d(FE_OFN195_n250395));
   in01s01 U269312 (.o(n185045),
	.a(n250414));
   oa22s01 U269313 (.o(n250415),
	.a(n250449),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[95]),
	.d(FE_OFN282_n250430));
   in01s01 U269314 (.o(n185046),
	.a(n250415));
   oa22s01 U269315 (.o(n250416),
	.a(n250449),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[94]),
	.d(FE_OFN282_n250430));
   in01s01 U269316 (.o(n185047),
	.a(n250416));
   oa22s01 U269317 (.o(n250417),
	.a(n250449),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[93]),
	.d(FE_OFN282_n250430));
   in01s01 U269318 (.o(n185048),
	.a(n250417));
   oa22s01 U269319 (.o(n250418),
	.a(n250449),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[92]),
	.d(FE_OFN282_n250430));
   in01s01 U269320 (.o(n185049),
	.a(n250418));
   oa22s01 U269321 (.o(n250419),
	.a(n250449),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[91]),
	.d(FE_OFN282_n250430));
   in01s01 U269322 (.o(n185050),
	.a(n250419));
   oa22s01 U269323 (.o(n250420),
	.a(n250449),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[90]),
	.d(FE_OFN282_n250430));
   in01s01 U269324 (.o(n185051),
	.a(n250420));
   oa22s01 U269325 (.o(n250421),
	.a(n250449),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[89]),
	.d(FE_OFN282_n250430));
   in01s01 U269326 (.o(n185052),
	.a(n250421));
   oa22s01 U269327 (.o(n250422),
	.a(n250449),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[88]),
	.d(FE_OFN282_n250430));
   in01s01 U269328 (.o(n185053),
	.a(n250422));
   oa22s01 U269329 (.o(n250423),
	.a(n250449),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[87]),
	.d(FE_OFN282_n250430));
   in01s01 U269330 (.o(n185054),
	.a(n250423));
   oa22s01 U269331 (.o(n250424),
	.a(n250449),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[86]),
	.d(FE_OFN282_n250430));
   oa22s01 U269332 (.o(n250425),
	.a(n250449),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[85]),
	.d(FE_OFN282_n250430));
   in01s01 U269333 (.o(n185056),
	.a(n250425));
   oa22s01 U269334 (.o(n250426),
	.a(n250449),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[84]),
	.d(FE_OFN282_n250430));
   in01s01 U269335 (.o(n185057),
	.a(n250426));
   oa22s01 U269336 (.o(n250427),
	.a(n250449),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[83]),
	.d(FE_OFN282_n250430));
   in01s01 U269337 (.o(n185058),
	.a(n250427));
   oa22s01 U269338 (.o(n250428),
	.a(n250449),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[82]),
	.d(FE_OFN282_n250430));
   in01s01 U269339 (.o(n185059),
	.a(n250428));
   oa22s01 U269340 (.o(n250429),
	.a(n250449),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[81]),
	.d(FE_OFN282_n250430));
   in01s01 U269341 (.o(n185060),
	.a(n250429));
   oa22s01 U269342 (.o(n250431),
	.a(n250449),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[80]),
	.d(FE_OFN282_n250430));
   in01s01 U269343 (.o(n185061),
	.a(n250431));
   oa22s01 U269344 (.o(n250432),
	.a(n250449),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[79]),
	.d(FE_OFN282_n250430));
   in01s01 U269345 (.o(n185062),
	.a(n250432));
   oa22s01 U269346 (.o(n250433),
	.a(n250449),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[78]),
	.d(FE_OFN282_n250430));
   in01s01 U269347 (.o(n185063),
	.a(n250433));
   oa22s01 U269348 (.o(n250434),
	.a(n250449),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[77]),
	.d(FE_OFN282_n250430));
   in01s01 U269349 (.o(n185064),
	.a(n250434));
   oa22s01 U269350 (.o(n250435),
	.a(n250449),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[76]),
	.d(FE_OFN282_n250430));
   in01s01 U269351 (.o(n185065),
	.a(n250435));
   oa22s01 U269352 (.o(n250436),
	.a(n250449),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[75]),
	.d(FE_OFN282_n250430));
   in01s01 U269353 (.o(n185066),
	.a(n250436));
   oa22s01 U269354 (.o(n250437),
	.a(n250449),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[74]),
	.d(FE_OFN282_n250430));
   in01s01 U269355 (.o(n185067),
	.a(n250437));
   oa22s01 U269356 (.o(n250438),
	.a(n250449),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[73]),
	.d(FE_OFN282_n250430));
   in01s01 U269357 (.o(n185068),
	.a(n250438));
   oa22s01 U269358 (.o(n250439),
	.a(n250449),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[72]),
	.d(FE_OFN282_n250430));
   in01s01 U269359 (.o(n185069),
	.a(n250439));
   oa22s01 U269360 (.o(n250440),
	.a(n250449),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[71]),
	.d(FE_OFN282_n250430));
   oa22s01 U269361 (.o(n250442),
	.a(n250449),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[70]),
	.d(FE_OFN282_n250430));
   in01s01 U269362 (.o(n185071),
	.a(n250442));
   oa22s01 U269363 (.o(n250443),
	.a(n250449),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[69]),
	.d(FE_OFN282_n250430));
   in01s01 U269364 (.o(n185072),
	.a(n250443));
   oa22s01 U269365 (.o(n250444),
	.a(n250449),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[68]),
	.d(FE_OFN282_n250430));
   in01s01 U269366 (.o(n185073),
	.a(n250444));
   oa22s01 U269367 (.o(n250445),
	.a(n250449),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[67]),
	.d(FE_OFN282_n250430));
   in01s01 U269368 (.o(n185074),
	.a(n250445));
   oa22s01 U269369 (.o(n250446),
	.a(n250449),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[66]),
	.d(FE_OFN282_n250430));
   in01s01 U269370 (.o(n185075),
	.a(n250446));
   oa22s01 U269371 (.o(n250447),
	.a(n250449),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[65]),
	.d(FE_OFN282_n250430));
   in01s01 U269372 (.o(n185076),
	.a(n250447));
   oa22s01 U269373 (.o(n250450),
	.a(n250449),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[64]),
	.d(FE_OFN282_n250430));
   in01s01 U269374 (.o(n185077),
	.a(n250450));
   in01s01 U269375 (.o(n185078),
	.a(n250451));
   in01s01 U269376 (.o(n185079),
	.a(n250452));
   in01s01 U269377 (.o(n185080),
	.a(n250453));
   in01s01 U269378 (.o(n185081),
	.a(n250454));
   in01s01 U269379 (.o(n185082),
	.a(n250455));
   in01s01 U269380 (.o(n185083),
	.a(n250456));
   in01s01 U269381 (.o(n185084),
	.a(n250457));
   oa22s01 U269382 (.o(n250458),
	.a(n250484),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[56]),
	.d(FE_OFN284_n250466));
   in01s01 U269383 (.o(n185086),
	.a(n250459));
   in01s01 U269384 (.o(n185087),
	.a(n250460));
   in01s01 U269385 (.o(n185088),
	.a(n250461));
   in01s01 U269386 (.o(n185089),
	.a(n250462));
   in01s01 U269387 (.o(n185090),
	.a(n250463));
   in01s01 U269388 (.o(n185091),
	.a(n250464));
   in01s01 U269389 (.o(n185092),
	.a(n250465));
   in01s01 U269390 (.o(n185093),
	.a(n250467));
   in01s01 U269391 (.o(n185094),
	.a(n250468));
   in01s01 U269392 (.o(n185095),
	.a(n250469));
   in01s01 U269393 (.o(n185096),
	.a(n250470));
   in01s01 U269394 (.o(n185097),
	.a(n250471));
   in01s01 U269395 (.o(n185098),
	.a(n250472));
   in01s01 U269396 (.o(n185099),
	.a(n250473));
   oa22s01 U269397 (.o(n250474),
	.a(n250484),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[41]),
	.d(n250466));
   in01s01 U269398 (.o(n185101),
	.a(n250475));
   in01s01 U269399 (.o(n185102),
	.a(n250476));
   in01s01 U269400 (.o(n185103),
	.a(n250478));
   oa22s01 U269401 (.o(n250479),
	.a(n250484),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[37]),
	.d(FE_OFN284_n250466));
   in01s01 U269402 (.o(n185104),
	.a(n250479));
   oa22s01 U269403 (.o(n250480),
	.a(n250484),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[36]),
	.d(FE_OFN284_n250466));
   in01s01 U269404 (.o(n185105),
	.a(n250480));
   oa22s01 U269405 (.o(n250481),
	.a(n250484),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[35]),
	.d(FE_OFN284_n250466));
   in01s01 U269406 (.o(n185106),
	.a(n250481));
   oa22s01 U269407 (.o(n250482),
	.a(n250484),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[34]),
	.d(FE_OFN284_n250466));
   in01s01 U269408 (.o(n185107),
	.a(n250482));
   oa22s01 U269409 (.o(n250483),
	.a(n250484),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[33]),
	.d(FE_OFN284_n250466));
   in01s01 U269410 (.o(n185108),
	.a(n250483));
   oa22s01 U269411 (.o(n250485),
	.a(n250484),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[32]),
	.d(n250466));
   in01s01 U269412 (.o(n185109),
	.a(n250485));
   in01s01 U269413 (.o(n185110),
	.a(n250487));
   in01s01 U269414 (.o(n185111),
	.a(n250488));
   in01s01 U269415 (.o(n185112),
	.a(n250489));
   in01s01 U269416 (.o(n185113),
	.a(n250490));
   in01s01 U269417 (.o(n185114),
	.a(n250491));
   oa22s01 U269418 (.o(n250492),
	.a(n250520),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[26]),
	.d(FE_OFN286_n250502));
   in01s01 U269419 (.o(n185116),
	.a(n250493));
   in01s01 U269420 (.o(n185117),
	.a(n250494));
   in01s01 U269421 (.o(n185118),
	.a(n250495));
   in01s01 U269422 (.o(n185119),
	.a(n250496));
   in01s01 U269423 (.o(n185120),
	.a(n250497));
   in01s01 U269424 (.o(n185121),
	.a(n250498));
   in01s01 U269425 (.o(n185122),
	.a(n250499));
   in01s01 U269426 (.o(n185123),
	.a(n250500));
   in01s01 U269427 (.o(n185124),
	.a(n250501));
   in01s01 U269428 (.o(n185125),
	.a(n250503));
   in01s01 U269429 (.o(n185126),
	.a(n250504));
   in01s01 U269430 (.o(n185127),
	.a(n250505));
   in01s01 U269431 (.o(n185128),
	.a(n250506));
   in01s01 U269432 (.o(n185129),
	.a(n250507));
   oa22s01 U269433 (.o(n250508),
	.a(n250520),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[11]),
	.d(FE_OFN286_n250502));
   in01s01 U269434 (.o(n185131),
	.a(n250509));
   in01s01 U269435 (.o(n185132),
	.a(n250510));
   in01s01 U269436 (.o(n185133),
	.a(n250511));
   in01s01 U269437 (.o(n185134),
	.a(n250512));
   in01s01 U269438 (.o(n185135),
	.a(n250514));
   oa22s01 U269439 (.o(n250515),
	.a(n250520),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[5]),
	.d(FE_OFN286_n250502));
   in01s01 U269440 (.o(n185136),
	.a(n250515));
   oa22s01 U269441 (.o(n250516),
	.a(n250520),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[4]),
	.d(FE_OFN286_n250502));
   in01s01 U269442 (.o(n185137),
	.a(n250516));
   oa22s01 U269443 (.o(n250517),
	.a(n250520),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[3]),
	.d(FE_OFN286_n250502));
   in01s01 U269444 (.o(n185138),
	.a(n250517));
   oa22s01 U269445 (.o(n250518),
	.a(n250520),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[2]),
	.d(FE_OFN286_n250502));
   in01s01 U269446 (.o(n185139),
	.a(n250518));
   oa22s01 U269447 (.o(n250519),
	.a(n250520),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1]),
	.d(FE_OFN286_n250502));
   in01s01 U269448 (.o(n185140),
	.a(n250519));
   oa22s01 U269449 (.o(n250521),
	.a(n250520),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[0]),
	.d(n250502));
   in01s01 U269450 (.o(n185141),
	.a(n250521));
   in01s01 U269451 (.o(n185142),
	.a(n250522));
   in01s01 U269452 (.o(n185143),
	.a(n250523));
   in01s01 U269453 (.o(n185144),
	.a(n250524));
   oa22s01 U269454 (.o(n250525),
	.a(n250556),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1020]),
	.d(FE_OFN288_n250540));
   in01s01 U269455 (.o(n185146),
	.a(n250526));
   in01s01 U269456 (.o(n185147),
	.a(n250527));
   in01s01 U269457 (.o(n185148),
	.a(n250528));
   in01s01 U269458 (.o(n185149),
	.a(n250529));
   in01s01 U269459 (.o(n185150),
	.a(n250530));
   in01s01 U269460 (.o(n185151),
	.a(n250531));
   in01s01 U269461 (.o(n185152),
	.a(n250532));
   in01s01 U269462 (.o(n185153),
	.a(n250533));
   in01s01 U269463 (.o(n185154),
	.a(n250534));
   in01s01 U269464 (.o(n185155),
	.a(n250535));
   in01s01 U269465 (.o(n185156),
	.a(n250536));
   in01s01 U269466 (.o(n185157),
	.a(n250537));
   in01s01 U269467 (.o(n185158),
	.a(n250538));
   in01s01 U269468 (.o(n185159),
	.a(n250539));
   oa22s01 U269469 (.o(n250541),
	.a(n250556),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1005]),
	.d(FE_OFN288_n250540));
   in01s01 U269470 (.o(n185161),
	.a(n250542));
   in01s01 U269471 (.o(n185162),
	.a(n250543));
   in01s01 U269472 (.o(n185163),
	.a(n250544));
   in01s01 U269473 (.o(n185164),
	.a(n250545));
   in01s01 U269474 (.o(n185165),
	.a(n250546));
   in01s01 U269475 (.o(n185166),
	.a(n250547));
   in01s01 U269476 (.o(n185167),
	.a(n250549));
   oa22s01 U269477 (.o(n250550),
	.a(n250556),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[997]),
	.d(FE_OFN288_n250540));
   in01s01 U269478 (.o(n185168),
	.a(n250550));
   oa22s01 U269479 (.o(n250551),
	.a(n250556),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[996]),
	.d(FE_OFN288_n250540));
   in01s01 U269480 (.o(n185169),
	.a(n250551));
   oa22s01 U269481 (.o(n250552),
	.a(n250556),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[995]),
	.d(FE_OFN288_n250540));
   in01s01 U269482 (.o(n185170),
	.a(n250552));
   oa22s01 U269483 (.o(n250553),
	.a(n250556),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[994]),
	.d(FE_OFN288_n250540));
   in01s01 U269484 (.o(n185171),
	.a(n250553));
   oa22s01 U269485 (.o(n250554),
	.a(n250556),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[993]),
	.d(FE_OFN288_n250540));
   in01s01 U269486 (.o(n185172),
	.a(n250554));
   oa22s01 U269487 (.o(n250557),
	.a(n250556),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[992]),
	.d(FE_OFN288_n250540));
   in01s01 U269488 (.o(n185173),
	.a(n250557));
   in01s01 U269489 (.o(n185174),
	.a(n250558));
   oa22s01 U269490 (.o(n250559),
	.a(n250591),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[990]),
	.d(FE_OFN412_n250576));
   in01s01 U269491 (.o(n185176),
	.a(n250560));
   in01s01 U269492 (.o(n185177),
	.a(n250561));
   in01s01 U269493 (.o(n185178),
	.a(n250562));
   in01s01 U269494 (.o(n185179),
	.a(n250563));
   in01s01 U269495 (.o(n185180),
	.a(n250564));
   in01s01 U269496 (.o(n185181),
	.a(n250565));
   in01s01 U269497 (.o(n185182),
	.a(n250566));
   in01s01 U269498 (.o(n185183),
	.a(n250567));
   in01s01 U269499 (.o(n185184),
	.a(n250568));
   in01s01 U269500 (.o(n185185),
	.a(n250569));
   in01s01 U269501 (.o(n185186),
	.a(n250570));
   in01s01 U269502 (.o(n185187),
	.a(n250571));
   in01s01 U269503 (.o(n185188),
	.a(n250572));
   in01s01 U269504 (.o(n185189),
	.a(n250573));
   oa22s01 U269505 (.o(n250574),
	.a(n250591),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[975]),
	.d(FE_OFN412_n250576));
   in01s01 U269506 (.o(n185191),
	.a(n250575));
   in01s01 U269507 (.o(n185192),
	.a(n250577));
   in01s01 U269508 (.o(n185193),
	.a(n250578));
   in01s01 U269509 (.o(n185194),
	.a(n250579));
   in01s01 U269510 (.o(n185195),
	.a(n250580));
   in01s01 U269511 (.o(n185196),
	.a(n250581));
   in01s01 U269512 (.o(n185197),
	.a(n250582));
   in01s01 U269513 (.o(n185198),
	.a(n250583));
   in01s01 U269514 (.o(n185199),
	.a(n250585));
   oa22s01 U269515 (.o(n250586),
	.a(n250591),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[965]),
	.d(FE_OFN412_n250576));
   in01s01 U269516 (.o(n185200),
	.a(n250586));
   oa22s01 U269517 (.o(n250587),
	.a(n250591),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[964]),
	.d(FE_OFN412_n250576));
   in01s01 U269518 (.o(n185201),
	.a(n250587));
   oa22s01 U269519 (.o(n250588),
	.a(n250591),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[963]),
	.d(FE_OFN412_n250576));
   in01s01 U269520 (.o(n185202),
	.a(n250588));
   oa22s01 U269521 (.o(n250589),
	.a(n250591),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[962]),
	.d(FE_OFN412_n250576));
   in01s01 U269522 (.o(n185203),
	.a(n250589));
   oa22s01 U269523 (.o(n250590),
	.a(n250591),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[961]),
	.d(FE_OFN412_n250576));
   in01s01 U269524 (.o(n185204),
	.a(n250590));
   oa22s01 U269525 (.o(n250592),
	.a(n250591),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[960]),
	.d(FE_OFN412_n250576));
   in01s01 U269526 (.o(n185206),
	.a(n250593));
   in01s01 U269527 (.o(n185207),
	.a(n250594));
   in01s01 U269528 (.o(n185208),
	.a(n250595));
   in01s01 U269529 (.o(n185209),
	.a(n250596));
   in01s01 U269530 (.o(n185210),
	.a(n250597));
   in01s01 U269531 (.o(n185211),
	.a(n250598));
   in01s01 U269532 (.o(n185212),
	.a(n250599));
   in01s01 U269533 (.o(n185213),
	.a(n250600));
   in01s01 U269534 (.o(n185214),
	.a(n250601));
   in01s01 U269535 (.o(n185215),
	.a(n250602));
   in01s01 U269536 (.o(n185216),
	.a(n250603));
   in01s01 U269537 (.o(n185217),
	.a(n250604));
   in01s01 U269538 (.o(n185218),
	.a(n250605));
   in01s01 U269539 (.o(n185219),
	.a(n250606));
   oa22s01 U269540 (.o(n250607),
	.a(n250626),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[945]),
	.d(FE_OFN290_n250611));
   in01s01 U269541 (.o(n185221),
	.a(n250608));
   in01s01 U269542 (.o(n185222),
	.a(n250609));
   in01s01 U269543 (.o(n185223),
	.a(n250610));
   in01s01 U269544 (.o(n185224),
	.a(n250612));
   in01s01 U269545 (.o(n185225),
	.a(n250613));
   in01s01 U269546 (.o(n185226),
	.a(n250614));
   in01s01 U269547 (.o(n185227),
	.a(n250615));
   in01s01 U269548 (.o(n185228),
	.a(n250616));
   in01s01 U269549 (.o(n185229),
	.a(n250617));
   in01s01 U269550 (.o(n185230),
	.a(n250618));
   in01s01 U269551 (.o(n185231),
	.a(n250620));
   oa22s01 U269552 (.o(n250621),
	.a(n250626),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[933]),
	.d(FE_OFN290_n250611));
   in01s01 U269553 (.o(n185232),
	.a(n250621));
   oa22s01 U269554 (.o(n250622),
	.a(n250626),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[932]),
	.d(FE_OFN290_n250611));
   in01s01 U269555 (.o(n185233),
	.a(n250622));
   oa22s01 U269556 (.o(n250623),
	.a(n250626),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[931]),
	.d(FE_OFN290_n250611));
   in01s01 U269557 (.o(n185234),
	.a(n250623));
   oa22s01 U269558 (.o(n250624),
	.a(n250626),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[930]),
	.d(FE_OFN290_n250611));
   oa22s01 U269559 (.o(n250625),
	.a(n250626),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[929]),
	.d(FE_OFN290_n250611));
   in01s01 U269560 (.o(n185236),
	.a(n250625));
   oa22s01 U269561 (.o(n250627),
	.a(n250626),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[928]),
	.d(FE_OFN290_n250611));
   in01s01 U269562 (.o(n185237),
	.a(n250627));
   in01s01 U269563 (.o(n185238),
	.a(n250628));
   in01s01 U269564 (.o(n185239),
	.a(n250629));
   in01s01 U269565 (.o(n185240),
	.a(n250630));
   in01s01 U269566 (.o(n185241),
	.a(n250631));
   in01s01 U269567 (.o(n185242),
	.a(n250632));
   in01s01 U269568 (.o(n185243),
	.a(n250633));
   in01s01 U269569 (.o(n185244),
	.a(n250634));
   in01s01 U269570 (.o(n185245),
	.a(n250635));
   in01s01 U269571 (.o(n185246),
	.a(n250636));
   in01s01 U269572 (.o(n185247),
	.a(n250637));
   in01s01 U269573 (.o(n185248),
	.a(n250638));
   in01s01 U269574 (.o(n185249),
	.a(n250639));
   oa22s01 U269575 (.o(n250640),
	.a(n250662),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[915]),
	.d(FE_OFN414_n250646));
   in01s01 U269576 (.o(n185251),
	.a(n250641));
   in01s01 U269577 (.o(n185252),
	.a(n250642));
   in01s01 U269578 (.o(n185253),
	.a(n250643));
   in01s01 U269579 (.o(n185254),
	.a(n250644));
   in01s01 U269580 (.o(n185255),
	.a(n250645));
   in01s01 U269581 (.o(n185256),
	.a(n250647));
   in01s01 U269582 (.o(n185257),
	.a(n250648));
   in01s01 U269583 (.o(n185258),
	.a(n250649));
   in01s01 U269584 (.o(n185259),
	.a(n250650));
   in01s01 U269585 (.o(n185260),
	.a(n250651));
   in01s01 U269586 (.o(n185261),
	.a(n250652));
   in01s01 U269587 (.o(n185262),
	.a(n250653));
   in01s01 U269588 (.o(n185263),
	.a(n250655));
   oa22s01 U269589 (.o(n250656),
	.a(n250662),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[901]),
	.d(FE_OFN414_n250646));
   in01s01 U269590 (.o(n185264),
	.a(n250656));
   oa22s01 U269591 (.o(n250657),
	.a(n250662),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[900]),
	.d(FE_OFN414_n250646));
   oa22s01 U269592 (.o(n250658),
	.a(n250662),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[899]),
	.d(FE_OFN414_n250646));
   in01s01 U269593 (.o(n185266),
	.a(n250658));
   oa22s01 U269594 (.o(n250659),
	.a(n250662),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[898]),
	.d(FE_OFN414_n250646));
   in01s01 U269595 (.o(n185267),
	.a(n250659));
   oa22s01 U269596 (.o(n250660),
	.a(n250662),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[897]),
	.d(FE_OFN414_n250646));
   in01s01 U269597 (.o(n185268),
	.a(n250660));
   oa22s01 U269598 (.o(n250663),
	.a(n250662),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[896]),
	.d(FE_OFN414_n250646));
   in01s01 U269599 (.o(n185269),
	.a(n250663));
   in01s01 U269600 (.o(n185270),
	.a(n250664));
   in01s01 U269601 (.o(n185271),
	.a(n250665));
   in01s01 U269602 (.o(n185272),
	.a(n250666));
   in01s01 U269603 (.o(n185273),
	.a(n250667));
   in01s01 U269604 (.o(n185274),
	.a(n250668));
   in01s01 U269605 (.o(n185275),
	.a(n250669));
   in01s01 U269606 (.o(n185276),
	.a(n250670));
   in01s01 U269607 (.o(n185277),
	.a(n250671));
   in01s01 U269608 (.o(n185278),
	.a(n250672));
   in01s01 U269609 (.o(n185279),
	.a(n250673));
   oa22s01 U269610 (.o(n250674),
	.a(n250697),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[885]),
	.d(FE_OFN198_n250682));
   in01s01 U269611 (.o(n185281),
	.a(n250675));
   in01s01 U269612 (.o(n185282),
	.a(n250676));
   in01s01 U269613 (.o(n185283),
	.a(n250677));
   in01s01 U269614 (.o(n185284),
	.a(n250678));
   in01s01 U269615 (.o(n185285),
	.a(n250679));
   in01s01 U269616 (.o(n185286),
	.a(n250680));
   in01s01 U269617 (.o(n185287),
	.a(n250681));
   in01s01 U269618 (.o(n185288),
	.a(n250683));
   in01s01 U269619 (.o(n185289),
	.a(n250684));
   in01s01 U269620 (.o(n185290),
	.a(n250685));
   in01s01 U269621 (.o(n185291),
	.a(n250686));
   in01s01 U269622 (.o(n185292),
	.a(n250687));
   in01s01 U269623 (.o(n185293),
	.a(n250688));
   in01s01 U269624 (.o(n185294),
	.a(n250689));
   oa22s01 U269625 (.o(n250691),
	.a(n250697),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[870]),
	.d(n250682));
   oa22s01 U269626 (.o(n250692),
	.a(n250697),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[869]),
	.d(FE_OFN198_n250682));
   in01s01 U269627 (.o(n185296),
	.a(n250692));
   oa22s01 U269628 (.o(n250693),
	.a(n250697),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[868]),
	.d(FE_OFN198_n250682));
   in01s01 U269629 (.o(n185297),
	.a(n250693));
   oa22s01 U269630 (.o(n250694),
	.a(n250697),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[867]),
	.d(FE_OFN198_n250682));
   in01s01 U269631 (.o(n185298),
	.a(n250694));
   oa22s01 U269632 (.o(n250695),
	.a(n250697),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[866]),
	.d(FE_OFN198_n250682));
   in01s01 U269633 (.o(n185299),
	.a(n250695));
   oa22s01 U269634 (.o(n250696),
	.a(n250697),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[865]),
	.d(FE_OFN198_n250682));
   in01s01 U269635 (.o(n185300),
	.a(n250696));
   oa22s01 U269636 (.o(n250698),
	.a(n250697),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[864]),
	.d(n250682));
   in01s01 U269637 (.o(n185301),
	.a(n250698));
   in01s01 U269638 (.o(n185302),
	.a(n250699));
   in01s01 U269639 (.o(n185303),
	.a(n250700));
   in01s01 U269640 (.o(n185304),
	.a(n250701));
   in01s01 U269641 (.o(n185305),
	.a(n250702));
   in01s01 U269642 (.o(n185306),
	.a(n250703));
   in01s01 U269643 (.o(n185307),
	.a(n250704));
   oa22s01 U269644 (.o(n250705),
	.a(n250732),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[857]),
	.d(FE_OFN292_n250717));
   in01s01 U269645 (.o(n185308),
	.a(n250705));
   in01s01 U269646 (.o(n185309),
	.a(n250706));
   oa22s01 U269647 (.o(n250707),
	.a(n250732),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[855]),
	.d(FE_OFN292_n250717));
   in01s01 U269648 (.o(n185311),
	.a(n250708));
   oa22s01 U269649 (.o(n250709),
	.a(n250732),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[853]),
	.d(FE_OFN292_n250717));
   in01s01 U269650 (.o(n185312),
	.a(n250709));
   in01s01 U269651 (.o(n185313),
	.a(n250710));
   oa22s01 U269652 (.o(n250711),
	.a(n250732),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[851]),
	.d(FE_OFN292_n250717));
   in01s01 U269653 (.o(n185314),
	.a(n250711));
   in01s01 U269654 (.o(n185315),
	.a(n250712));
   oa22s01 U269655 (.o(n250713),
	.a(n250732),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[849]),
	.d(FE_OFN563_n250717));
   in01s01 U269656 (.o(n185316),
	.a(n250713));
   oa22s01 U269657 (.o(n250714),
	.a(n250732),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[848]),
	.d(FE_OFN563_n250717));
   in01s01 U269658 (.o(n185317),
	.a(n250714));
   in01s01 U269659 (.o(n185318),
	.a(n250715));
   in01s01 U269660 (.o(n185319),
	.a(n250716));
   oa22s01 U269661 (.o(n250718),
	.a(n250732),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[845]),
	.d(FE_OFN292_n250717));
   in01s01 U269662 (.o(n185320),
	.a(n250718));
   in01s01 U269663 (.o(n185321),
	.a(n250719));
   in01s01 U269664 (.o(n185322),
	.a(n250720));
   in01s01 U269665 (.o(n185323),
	.a(n250721));
   in01s01 U269666 (.o(n185324),
	.a(n250722));
   oa22s01 U269667 (.o(n250723),
	.a(n250732),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[840]),
	.d(FE_OFN563_n250717));
   in01s01 U269668 (.o(n185326),
	.a(n250724));
   in01s01 U269669 (.o(n185327),
	.a(n250726));
   oa22s01 U269670 (.o(n250727),
	.a(n250732),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[837]),
	.d(FE_OFN563_n250717));
   in01s01 U269671 (.o(n185328),
	.a(n250727));
   oa22s01 U269672 (.o(n250728),
	.a(n250732),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[836]),
	.d(FE_OFN563_n250717));
   in01s01 U269673 (.o(n185329),
	.a(n250728));
   oa22s01 U269674 (.o(n250729),
	.a(n250732),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[835]),
	.d(FE_OFN563_n250717));
   in01s01 U269675 (.o(n185330),
	.a(n250729));
   oa22s01 U269676 (.o(n250730),
	.a(n250732),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[834]),
	.d(FE_OFN563_n250717));
   in01s01 U269677 (.o(n185331),
	.a(n250730));
   oa22s01 U269678 (.o(n250731),
	.a(n250732),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[833]),
	.d(FE_OFN563_n250717));
   in01s01 U269679 (.o(n185332),
	.a(n250731));
   oa22s01 U269680 (.o(n250733),
	.a(n250732),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[832]),
	.d(FE_OFN292_n250717));
   in01s01 U269681 (.o(n185333),
	.a(n250733));
   in01s01 U269682 (.o(n185334),
	.a(n250734));
   in01s01 U269683 (.o(n185335),
	.a(n250735));
   in01s01 U269684 (.o(n185336),
	.a(n250736));
   in01s01 U269685 (.o(n185337),
	.a(n250737));
   in01s01 U269686 (.o(n185338),
	.a(n250738));
   in01s01 U269687 (.o(n185339),
	.a(n250739));
   oa22s01 U269688 (.o(n250740),
	.a(n250768),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[825]),
	.d(FE_OFN294_n250752));
   in01s01 U269689 (.o(n185341),
	.a(n250741));
   in01s01 U269690 (.o(n185342),
	.a(n250742));
   in01s01 U269691 (.o(n185343),
	.a(n250743));
   in01s01 U269692 (.o(n185344),
	.a(n250744));
   in01s01 U269693 (.o(n185345),
	.a(n250745));
   in01s01 U269694 (.o(n185346),
	.a(n250746));
   in01s01 U269695 (.o(n185347),
	.a(n250747));
   in01s01 U269696 (.o(n185348),
	.a(n250748));
   in01s01 U269697 (.o(n185349),
	.a(n250749));
   in01s01 U269698 (.o(n185350),
	.a(n250750));
   in01s01 U269699 (.o(n185351),
	.a(n250751));
   in01s01 U269700 (.o(n185352),
	.a(n250753));
   in01s01 U269701 (.o(n185353),
	.a(n250754));
   in01s01 U269702 (.o(n185354),
	.a(n250755));
   oa22s01 U269703 (.o(n250756),
	.a(n250768),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[810]),
	.d(FE_OFN294_n250752));
   in01s01 U269704 (.o(n185356),
	.a(n250757));
   in01s01 U269705 (.o(n185357),
	.a(n250758));
   in01s01 U269706 (.o(n185358),
	.a(n250759));
   in01s01 U269707 (.o(n185359),
	.a(n250761));
   oa22s01 U269708 (.o(n250762),
	.a(n250768),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[805]),
	.d(FE_OFN294_n250752));
   in01s01 U269709 (.o(n185360),
	.a(n250762));
   oa22s01 U269710 (.o(n250763),
	.a(n250768),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[804]),
	.d(FE_OFN294_n250752));
   in01s01 U269711 (.o(n185361),
	.a(n250763));
   oa22s01 U269712 (.o(n250764),
	.a(n250768),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[803]),
	.d(FE_OFN294_n250752));
   in01s01 U269713 (.o(n185362),
	.a(n250764));
   oa22s01 U269714 (.o(n250765),
	.a(n250768),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[802]),
	.d(FE_OFN294_n250752));
   in01s01 U269715 (.o(n185363),
	.a(n250765));
   oa22s01 U269716 (.o(n250766),
	.a(n250768),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[801]),
	.d(FE_OFN294_n250752));
   in01s01 U269717 (.o(n185364),
	.a(n250766));
   oa22s01 U269718 (.o(n250769),
	.a(n250768),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[800]),
	.d(FE_OFN294_n250752));
   in01s01 U269719 (.o(n185365),
	.a(n250769));
   in01s01 U269720 (.o(n185366),
	.a(n250771));
   in01s01 U269721 (.o(n185367),
	.a(n250772));
   in01s01 U269722 (.o(n185368),
	.a(n250773));
   in01s01 U269723 (.o(n185369),
	.a(n250774));
   oa22s01 U269724 (.o(n250775),
	.a(n250804),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[795]),
	.d(FE_OFN296_n250789));
   in01s01 U269725 (.o(n185371),
	.a(n250776));
   in01s01 U269726 (.o(n185372),
	.a(n250777));
   in01s01 U269727 (.o(n185373),
	.a(n250778));
   in01s01 U269728 (.o(n185374),
	.a(n250779));
   in01s01 U269729 (.o(n185375),
	.a(n250780));
   in01s01 U269730 (.o(n185376),
	.a(n250781));
   in01s01 U269731 (.o(n185377),
	.a(n250782));
   in01s01 U269732 (.o(n185378),
	.a(n250783));
   in01s01 U269733 (.o(n185379),
	.a(n250784));
   in01s01 U269734 (.o(n185380),
	.a(n250785));
   in01s01 U269735 (.o(n185381),
	.a(n250786));
   in01s01 U269736 (.o(n185382),
	.a(n250787));
   in01s01 U269737 (.o(n185383),
	.a(n250788));
   in01s01 U269738 (.o(n185384),
	.a(n250790));
   oa22s01 U269739 (.o(n250791),
	.a(n250804),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[780]),
	.d(FE_OFN296_n250789));
   in01s01 U269740 (.o(n185386),
	.a(n250792));
   in01s01 U269741 (.o(n185387),
	.a(n250793));
   in01s01 U269742 (.o(n185388),
	.a(n250794));
   in01s01 U269743 (.o(n185389),
	.a(n250795));
   in01s01 U269744 (.o(n185390),
	.a(n250796));
   in01s01 U269745 (.o(n185391),
	.a(n250798));
   oa22s01 U269746 (.o(n250799),
	.a(n250804),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[773]),
	.d(FE_OFN296_n250789));
   in01s01 U269747 (.o(n185392),
	.a(n250799));
   oa22s01 U269748 (.o(n250800),
	.a(n250804),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[772]),
	.d(FE_OFN296_n250789));
   in01s01 U269749 (.o(n185393),
	.a(n250800));
   oa22s01 U269750 (.o(n250801),
	.a(n250804),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[771]),
	.d(FE_OFN296_n250789));
   in01s01 U269751 (.o(n185394),
	.a(n250801));
   oa22s01 U269752 (.o(n250802),
	.a(n250804),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[770]),
	.d(FE_OFN296_n250789));
   in01s01 U269753 (.o(n185395),
	.a(n250802));
   oa22s01 U269754 (.o(n250803),
	.a(n250804),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[769]),
	.d(FE_OFN296_n250789));
   in01s01 U269755 (.o(n185396),
	.a(n250803));
   oa22s01 U269756 (.o(n250805),
	.a(n250804),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[768]),
	.d(FE_OFN296_n250789));
   in01s01 U269757 (.o(n185397),
	.a(n250805));
   in01s01 U269758 (.o(n185398),
	.a(n250806));
   in01s01 U269759 (.o(n185399),
	.a(n250807));
   oa22s01 U269760 (.o(n250808),
	.a(n250839),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[765]),
	.d(FE_OFN298_n250824));
   in01s01 U269761 (.o(n185401),
	.a(n250809));
   in01s01 U269762 (.o(n185402),
	.a(n250810));
   in01s01 U269763 (.o(n185403),
	.a(n250811));
   in01s01 U269764 (.o(n185404),
	.a(n250812));
   in01s01 U269765 (.o(n185405),
	.a(n250813));
   in01s01 U269766 (.o(n185406),
	.a(n250814));
   in01s01 U269767 (.o(n185407),
	.a(n250815));
   in01s01 U269768 (.o(n185408),
	.a(n250816));
   in01s01 U269769 (.o(n185409),
	.a(n250817));
   in01s01 U269770 (.o(n185410),
	.a(n250818));
   in01s01 U269771 (.o(n185411),
	.a(n250819));
   in01s01 U269772 (.o(n185412),
	.a(n250820));
   in01s01 U269773 (.o(n185413),
	.a(n250821));
   in01s01 U269774 (.o(n185414),
	.a(n250822));
   oa22s01 U269775 (.o(n250823),
	.a(n250839),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[750]),
	.d(FE_OFN298_n250824));
   in01s01 U269776 (.o(n185416),
	.a(n250825));
   in01s01 U269777 (.o(n185417),
	.a(n250826));
   in01s01 U269778 (.o(n185418),
	.a(n250827));
   in01s01 U269779 (.o(n185419),
	.a(n250828));
   in01s01 U269780 (.o(n185420),
	.a(n250829));
   in01s01 U269781 (.o(n185421),
	.a(n250830));
   in01s01 U269782 (.o(n185422),
	.a(n250831));
   in01s01 U269783 (.o(n185423),
	.a(n250833));
   oa22s01 U269784 (.o(n250834),
	.a(n250839),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[741]),
	.d(FE_OFN298_n250824));
   in01s01 U269785 (.o(n185424),
	.a(n250834));
   oa22s01 U269786 (.o(n250835),
	.a(n250839),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[740]),
	.d(FE_OFN298_n250824));
   in01s01 U269787 (.o(n185425),
	.a(n250835));
   oa22s01 U269788 (.o(n250836),
	.a(n250839),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[739]),
	.d(n250824));
   in01s01 U269789 (.o(n185426),
	.a(n250836));
   oa22s01 U269790 (.o(n250837),
	.a(n250839),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[738]),
	.d(FE_OFN298_n250824));
   in01s01 U269791 (.o(n185427),
	.a(n250837));
   oa22s01 U269792 (.o(n250838),
	.a(n250839),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[737]),
	.d(FE_OFN298_n250824));
   in01s01 U269793 (.o(n185428),
	.a(n250838));
   oa22s01 U269794 (.o(n250840),
	.a(n250839),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[736]),
	.d(FE_OFN298_n250824));
   in01s01 U269795 (.o(n185429),
	.a(n250840));
   oa22s01 U269796 (.o(n250841),
	.a(n250875),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[735]),
	.d(FE_OFN416_n250859));
   in01s01 U269797 (.o(n185431),
	.a(n250842));
   in01s01 U269798 (.o(n185432),
	.a(n250843));
   in01s01 U269799 (.o(n185433),
	.a(n250844));
   in01s01 U269800 (.o(n185434),
	.a(n250845));
   in01s01 U269801 (.o(n185435),
	.a(n250846));
   in01s01 U269802 (.o(n185436),
	.a(n250847));
   in01s01 U269803 (.o(n185437),
	.a(n250848));
   in01s01 U269804 (.o(n185438),
	.a(n250849));
   in01s01 U269805 (.o(n185439),
	.a(n250850));
   in01s01 U269806 (.o(n185440),
	.a(n250851));
   in01s01 U269807 (.o(n185441),
	.a(n250852));
   in01s01 U269808 (.o(n185442),
	.a(n250853));
   in01s01 U269809 (.o(n185443),
	.a(n250854));
   in01s01 U269810 (.o(n185444),
	.a(n250855));
   oa22s01 U269811 (.o(n250856),
	.a(n250875),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[720]),
	.d(FE_OFN416_n250859));
   in01s01 U269812 (.o(n185446),
	.a(n250857));
   in01s01 U269813 (.o(n185447),
	.a(n250858));
   in01s01 U269814 (.o(n185448),
	.a(n250860));
   in01s01 U269815 (.o(n185449),
	.a(n250861));
   in01s01 U269816 (.o(n185450),
	.a(n250862));
   in01s01 U269817 (.o(n185451),
	.a(n250863));
   in01s01 U269818 (.o(n185452),
	.a(n250864));
   in01s01 U269819 (.o(n185453),
	.a(n250865));
   in01s01 U269820 (.o(n185454),
	.a(n250866));
   in01s01 U269821 (.o(n185455),
	.a(n250868));
   oa22s01 U269822 (.o(n250869),
	.a(n250875),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[709]),
	.d(FE_OFN416_n250859));
   in01s01 U269823 (.o(n185456),
	.a(n250869));
   oa22s01 U269824 (.o(n250870),
	.a(n250875),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[708]),
	.d(FE_OFN416_n250859));
   in01s01 U269825 (.o(n185457),
	.a(n250870));
   oa22s01 U269826 (.o(n250871),
	.a(n250875),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[707]),
	.d(FE_OFN416_n250859));
   in01s01 U269827 (.o(n185458),
	.a(n250871));
   oa22s01 U269828 (.o(n250872),
	.a(n250875),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[706]),
	.d(FE_OFN416_n250859));
   in01s01 U269829 (.o(n185459),
	.a(n250872));
   oa22s01 U269830 (.o(n250873),
	.a(n250875),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[705]),
	.d(FE_OFN416_n250859));
   oa22s01 U269831 (.o(n250876),
	.a(n250875),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[704]),
	.d(FE_OFN416_n250859));
   in01s01 U269832 (.o(n185461),
	.a(n250876));
   in01s01 U269833 (.o(n185462),
	.a(n250877));
   in01s01 U269834 (.o(n185463),
	.a(n250878));
   in01s01 U269835 (.o(n185464),
	.a(n250879));
   in01s01 U269836 (.o(n185465),
	.a(n250880));
   in01s01 U269837 (.o(n185466),
	.a(n250881));
   in01s01 U269838 (.o(n185467),
	.a(n250882));
   in01s01 U269839 (.o(n185468),
	.a(n250883));
   in01s01 U269840 (.o(n185469),
	.a(n250884));
   in01s01 U269841 (.o(n185470),
	.a(n250885));
   in01s01 U269842 (.o(n185471),
	.a(n250886));
   in01s01 U269843 (.o(n185472),
	.a(n250887));
   in01s01 U269844 (.o(n185473),
	.a(n250888));
   in01s01 U269845 (.o(n185474),
	.a(n250889));
   oa22s01 U269846 (.o(n250890),
	.a(n250910),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[690]),
	.d(FE_OFN300_n250895));
   in01s01 U269847 (.o(n185476),
	.a(n250891));
   in01s01 U269848 (.o(n185477),
	.a(n250892));
   in01s01 U269849 (.o(n185478),
	.a(n250893));
   in01s01 U269850 (.o(n185479),
	.a(n250894));
   in01s01 U269851 (.o(n185480),
	.a(n250896));
   in01s01 U269852 (.o(n185481),
	.a(n250897));
   in01s01 U269853 (.o(n185482),
	.a(n250898));
   in01s01 U269854 (.o(n185483),
	.a(n250899));
   in01s01 U269855 (.o(n185484),
	.a(n250900));
   in01s01 U269856 (.o(n185485),
	.a(n250901));
   in01s01 U269857 (.o(n185486),
	.a(n250902));
   in01s01 U269858 (.o(n185487),
	.a(n250904));
   oa22s01 U269859 (.o(n250905),
	.a(n250910),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[677]),
	.d(FE_OFN300_n250895));
   in01s01 U269860 (.o(n185488),
	.a(n250905));
   oa22s01 U269861 (.o(n250906),
	.a(n250910),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[676]),
	.d(FE_OFN300_n250895));
   in01s01 U269862 (.o(n185489),
	.a(n250906));
   oa22s01 U269863 (.o(n250907),
	.a(n250910),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[675]),
	.d(FE_OFN300_n250895));
   oa22s01 U269864 (.o(n250908),
	.a(n250910),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[674]),
	.d(FE_OFN300_n250895));
   in01s01 U269865 (.o(n185491),
	.a(n250908));
   oa22s01 U269866 (.o(n250909),
	.a(n250910),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[673]),
	.d(FE_OFN300_n250895));
   in01s01 U269867 (.o(n185492),
	.a(n250909));
   oa22s01 U269868 (.o(n250911),
	.a(n250910),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[672]),
	.d(FE_OFN300_n250895));
   in01s01 U269869 (.o(n185493),
	.a(n250911));
   in01s01 U269870 (.o(n185494),
	.a(n250912));
   in01s01 U269871 (.o(n185495),
	.a(n250913));
   in01s01 U269872 (.o(n185496),
	.a(n250914));
   in01s01 U269873 (.o(n185497),
	.a(n250915));
   in01s01 U269874 (.o(n185498),
	.a(n250916));
   in01s01 U269875 (.o(n185499),
	.a(n250917));
   in01s01 U269876 (.o(n185500),
	.a(n250918));
   in01s01 U269877 (.o(n185501),
	.a(n250919));
   in01s01 U269878 (.o(n185502),
	.a(n250920));
   in01s01 U269879 (.o(n185503),
	.a(n250921));
   in01s01 U269880 (.o(n185504),
	.a(n250922));
   oa22s01 U269881 (.o(n250923),
	.a(n250945),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[660]),
	.d(FE_OFN418_n250930));
   in01s01 U269882 (.o(n185506),
	.a(n250924));
   in01s01 U269883 (.o(n185507),
	.a(n250925));
   in01s01 U269884 (.o(n185508),
	.a(n250926));
   in01s01 U269885 (.o(n185509),
	.a(n250927));
   in01s01 U269886 (.o(n185510),
	.a(n250928));
   in01s01 U269887 (.o(n185511),
	.a(n250929));
   in01s01 U269888 (.o(n185512),
	.a(n250931));
   in01s01 U269889 (.o(n185513),
	.a(n250932));
   in01s01 U269890 (.o(n185514),
	.a(n250933));
   in01s01 U269891 (.o(n185515),
	.a(n250934));
   in01s01 U269892 (.o(n185516),
	.a(n250935));
   in01s01 U269893 (.o(n185517),
	.a(n250936));
   in01s01 U269894 (.o(n185518),
	.a(n250937));
   in01s01 U269895 (.o(n185519),
	.a(n250939));
   oa22s01 U269896 (.o(n250940),
	.a(n250945),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[645]),
	.d(FE_OFN418_n250930));
   oa22s01 U269897 (.o(n250941),
	.a(n250945),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[644]),
	.d(FE_OFN418_n250930));
   in01s01 U269898 (.o(n185521),
	.a(n250941));
   oa22s01 U269899 (.o(n250942),
	.a(n250945),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[643]),
	.d(FE_OFN418_n250930));
   in01s01 U269900 (.o(n185522),
	.a(n250942));
   oa22s01 U269901 (.o(n250943),
	.a(n250945),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[642]),
	.d(FE_OFN418_n250930));
   in01s01 U269902 (.o(n185523),
	.a(n250943));
   oa22s01 U269903 (.o(n250944),
	.a(n250945),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[641]),
	.d(FE_OFN418_n250930));
   in01s01 U269904 (.o(n185524),
	.a(n250944));
   oa22s01 U269905 (.o(n250946),
	.a(n250945),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[640]),
	.d(FE_OFN418_n250930));
   in01s01 U269906 (.o(n185525),
	.a(n250946));
   in01s01 U269907 (.o(n185526),
	.a(n250947));
   in01s01 U269908 (.o(n185527),
	.a(n250948));
   in01s01 U269909 (.o(n185528),
	.a(n250949));
   in01s01 U269910 (.o(n185529),
	.a(n250950));
   in01s01 U269911 (.o(n185530),
	.a(n250951));
   in01s01 U269912 (.o(n185531),
	.a(n250952));
   in01s01 U269913 (.o(n185532),
	.a(n250953));
   in01s01 U269914 (.o(n185533),
	.a(n250954));
   in01s01 U269915 (.o(n185534),
	.a(n250955));
   oa22s01 U269916 (.o(n250956),
	.a(n250981),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[630]),
	.d(FE_OFN200_n250965));
   in01s01 U269917 (.o(n185536),
	.a(n250957));
   in01s01 U269918 (.o(n185537),
	.a(n250958));
   in01s01 U269919 (.o(n185538),
	.a(n250959));
   in01s01 U269920 (.o(n185539),
	.a(n250960));
   in01s01 U269921 (.o(n185540),
	.a(n250961));
   in01s01 U269922 (.o(n185541),
	.a(n250962));
   in01s01 U269923 (.o(n185542),
	.a(n250963));
   in01s01 U269924 (.o(n185543),
	.a(n250964));
   in01s01 U269925 (.o(n185544),
	.a(n250966));
   in01s01 U269926 (.o(n185545),
	.a(n250967));
   in01s01 U269927 (.o(n185546),
	.a(n250968));
   in01s01 U269928 (.o(n185547),
	.a(n250969));
   in01s01 U269929 (.o(n185548),
	.a(n250970));
   in01s01 U269930 (.o(n185549),
	.a(n250971));
   oa22s01 U269931 (.o(n250972),
	.a(n250981),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[615]),
	.d(FE_OFN200_n250965));
   in01s01 U269932 (.o(n185551),
	.a(n250974));
   oa22s01 U269933 (.o(n250975),
	.a(n250981),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[613]),
	.d(FE_OFN200_n250965));
   in01s01 U269934 (.o(n185552),
	.a(n250975));
   oa22s01 U269935 (.o(n250976),
	.a(n250981),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[612]),
	.d(FE_OFN200_n250965));
   in01s01 U269936 (.o(n185553),
	.a(n250976));
   oa22s01 U269937 (.o(n250977),
	.a(n250981),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[611]),
	.d(FE_OFN200_n250965));
   in01s01 U269938 (.o(n185554),
	.a(n250977));
   oa22s01 U269939 (.o(n250978),
	.a(n250981),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[610]),
	.d(FE_OFN200_n250965));
   in01s01 U269940 (.o(n185555),
	.a(n250978));
   oa22s01 U269941 (.o(n250979),
	.a(n250981),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[609]),
	.d(FE_OFN200_n250965));
   in01s01 U269942 (.o(n185556),
	.a(n250979));
   oa22s01 U269943 (.o(n250982),
	.a(n250981),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[608]),
	.d(FE_OFN200_n250965));
   in01s01 U269944 (.o(n185557),
	.a(n250982));
   oa22s01 U269945 (.o(n250983),
	.a(n251016),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[607]),
	.d(FE_OFN302_n251001));
   in01s01 U269946 (.o(n185558),
	.a(n250983));
   oa22s01 U269947 (.o(n250984),
	.a(n251016),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[606]),
	.d(FE_OFN302_n251001));
   in01s01 U269948 (.o(n185559),
	.a(n250984));
   oa22s01 U269949 (.o(n250985),
	.a(n251016),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[605]),
	.d(FE_OFN302_n251001));
   in01s01 U269950 (.o(n185560),
	.a(n250985));
   oa22s01 U269951 (.o(n250986),
	.a(n251016),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[604]),
	.d(FE_OFN302_n251001));
   in01s01 U269952 (.o(n185561),
	.a(n250986));
   oa22s01 U269953 (.o(n250987),
	.a(n251016),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[603]),
	.d(FE_OFN302_n251001));
   in01s01 U269954 (.o(n185562),
	.a(n250987));
   in01s01 U269955 (.o(n185563),
	.a(n250988));
   oa22s01 U269956 (.o(n250989),
	.a(n251016),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[601]),
	.d(FE_OFN302_n251001));
   in01s01 U269957 (.o(n185564),
	.a(n250989));
   oa22s01 U269958 (.o(n250990),
	.a(n251016),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[600]),
	.d(FE_OFN302_n251001));
   oa22s01 U269959 (.o(n250991),
	.a(n251016),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[599]),
	.d(FE_OFN302_n251001));
   in01s01 U269960 (.o(n185566),
	.a(n250991));
   in01s01 U269961 (.o(n185567),
	.a(n250992));
   oa22s01 U269962 (.o(n250993),
	.a(n251016),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[597]),
	.d(FE_OFN302_n251001));
   in01s01 U269963 (.o(n185568),
	.a(n250993));
   in01s01 U269964 (.o(n185569),
	.a(n250994));
   oa22s01 U269965 (.o(n250995),
	.a(n251016),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[595]),
	.d(FE_OFN302_n251001));
   in01s01 U269966 (.o(n185570),
	.a(n250995));
   in01s01 U269967 (.o(n185571),
	.a(n250996));
   oa22s01 U269968 (.o(n250997),
	.a(n251016),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[593]),
	.d(FE_OFN302_n251001));
   in01s01 U269969 (.o(n185572),
	.a(n250997));
   oa22s01 U269970 (.o(n250998),
	.a(n251016),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[592]),
	.d(FE_OFN302_n251001));
   in01s01 U269971 (.o(n185573),
	.a(n250998));
   in01s01 U269972 (.o(n185574),
	.a(n250999));
   in01s01 U269973 (.o(n185575),
	.a(n251000));
   oa22s01 U269974 (.o(n251002),
	.a(n251016),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[589]),
	.d(FE_OFN302_n251001));
   in01s01 U269975 (.o(n185576),
	.a(n251002));
   oa22s01 U269976 (.o(n251003),
	.a(n251016),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[588]),
	.d(FE_OFN302_n251001));
   in01s01 U269977 (.o(n185577),
	.a(n251003));
   oa22s01 U269978 (.o(n251004),
	.a(n251016),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[587]),
	.d(FE_OFN302_n251001));
   in01s01 U269979 (.o(n185578),
	.a(n251004));
   oa22s01 U269980 (.o(n251005),
	.a(n251016),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[586]),
	.d(FE_OFN302_n251001));
   in01s01 U269981 (.o(n185579),
	.a(n251005));
   oa22s01 U269982 (.o(n251006),
	.a(n251016),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[585]),
	.d(FE_OFN302_n251001));
   in01s01 U269983 (.o(n185581),
	.a(n251007));
   in01s01 U269984 (.o(n185582),
	.a(n251008));
   in01s01 U269985 (.o(n185583),
	.a(n251010));
   oa22s01 U269986 (.o(n251011),
	.a(n251016),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[581]),
	.d(FE_OFN302_n251001));
   in01s01 U269987 (.o(n185584),
	.a(n251011));
   oa22s01 U269988 (.o(n251012),
	.a(n251016),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[580]),
	.d(FE_OFN302_n251001));
   in01s01 U269989 (.o(n185585),
	.a(n251012));
   oa22s01 U269990 (.o(n251013),
	.a(n251016),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[579]),
	.d(FE_OFN302_n251001));
   in01s01 U269991 (.o(n185586),
	.a(n251013));
   oa22s01 U269992 (.o(n251014),
	.a(n251016),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[578]),
	.d(FE_OFN302_n251001));
   in01s01 U269993 (.o(n185587),
	.a(n251014));
   oa22s01 U269994 (.o(n251015),
	.a(n251016),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[577]),
	.d(FE_OFN302_n251001));
   in01s01 U269995 (.o(n185588),
	.a(n251015));
   oa22s01 U269996 (.o(n251017),
	.a(n251016),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[576]),
	.d(FE_OFN302_n251001));
   in01s01 U269997 (.o(n185589),
	.a(n251017));
   in01s01 U269998 (.o(n185590),
	.a(n251018));
   in01s01 U269999 (.o(n185591),
	.a(n251019));
   in01s01 U270000 (.o(n185592),
	.a(n251020));
   in01s01 U270001 (.o(n185593),
	.a(n251021));
   in01s01 U270002 (.o(n185594),
	.a(n251022));
   oa22s01 U270003 (.o(n251023),
	.a(n251051),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[570]),
	.d(FE_OFN304_n251036));
   in01s01 U270004 (.o(n185596),
	.a(n251024));
   in01s01 U270005 (.o(n185597),
	.a(n251025));
   in01s01 U270006 (.o(n185598),
	.a(n251026));
   in01s01 U270007 (.o(n185599),
	.a(n251027));
   in01s01 U270008 (.o(n185600),
	.a(n251028));
   in01s01 U270009 (.o(n185601),
	.a(n251029));
   in01s01 U270010 (.o(n185602),
	.a(n251030));
   in01s01 U270011 (.o(n185603),
	.a(n251031));
   in01s01 U270012 (.o(n185604),
	.a(n251032));
   in01s01 U270013 (.o(n185605),
	.a(n251033));
   in01s01 U270014 (.o(n185606),
	.a(n251034));
   in01s01 U270015 (.o(n185607),
	.a(n251035));
   in01s01 U270016 (.o(n185608),
	.a(n251037));
   in01s01 U270017 (.o(n185609),
	.a(n251038));
   oa22s01 U270018 (.o(n251039),
	.a(n251051),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[555]),
	.d(FE_OFN304_n251036));
   in01s01 U270019 (.o(n185611),
	.a(n251040));
   in01s01 U270020 (.o(n185612),
	.a(n251041));
   in01s01 U270021 (.o(n185613),
	.a(n251042));
   in01s01 U270022 (.o(n185614),
	.a(n251043));
   in01s01 U270023 (.o(n185615),
	.a(n251045));
   oa22s01 U270024 (.o(n251046),
	.a(n251051),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[549]),
	.d(FE_OFN304_n251036));
   in01s01 U270025 (.o(n185616),
	.a(n251046));
   oa22s01 U270026 (.o(n251047),
	.a(n251051),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[548]),
	.d(FE_OFN304_n251036));
   in01s01 U270027 (.o(n185617),
	.a(n251047));
   oa22s01 U270028 (.o(n251048),
	.a(n251051),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[547]),
	.d(FE_OFN304_n251036));
   in01s01 U270029 (.o(n185618),
	.a(n251048));
   oa22s01 U270030 (.o(n251049),
	.a(n251051),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[546]),
	.d(FE_OFN304_n251036));
   in01s01 U270031 (.o(n185619),
	.a(n251049));
   oa22s01 U270032 (.o(n251050),
	.a(n251051),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[545]),
	.d(FE_OFN304_n251036));
   in01s01 U270033 (.o(n185620),
	.a(n251050));
   oa22s01 U270034 (.o(n251052),
	.a(n251051),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[544]),
	.d(FE_OFN304_n251036));
   in01s01 U270035 (.o(n185621),
	.a(n251052));
   in01s01 U270036 (.o(n185622),
	.a(n251054));
   in01s01 U270037 (.o(n185623),
	.a(n251055));
   in01s01 U270038 (.o(n185624),
	.a(n251056));
   oa22s01 U270039 (.o(n251057),
	.a(n251088),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[540]),
	.d(FE_OFN306_n251072));
   in01s01 U270040 (.o(n185626),
	.a(n251058));
   in01s01 U270041 (.o(n185627),
	.a(n251059));
   in01s01 U270042 (.o(n185628),
	.a(n251060));
   in01s01 U270043 (.o(n185629),
	.a(n251061));
   in01s01 U270044 (.o(n185630),
	.a(n251062));
   in01s01 U270045 (.o(n185631),
	.a(n251063));
   in01s01 U270046 (.o(n185632),
	.a(n251064));
   in01s01 U270047 (.o(n185633),
	.a(n251065));
   in01s01 U270048 (.o(n185634),
	.a(n251066));
   in01s01 U270049 (.o(n185635),
	.a(n251067));
   in01s01 U270050 (.o(n185636),
	.a(n251068));
   in01s01 U270051 (.o(n185637),
	.a(n251069));
   in01s01 U270052 (.o(n185638),
	.a(n251070));
   in01s01 U270053 (.o(n185639),
	.a(n251071));
   oa22s01 U270054 (.o(n251073),
	.a(n251088),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[525]),
	.d(FE_OFN306_n251072));
   in01s01 U270055 (.o(n185641),
	.a(n251074));
   in01s01 U270056 (.o(n185642),
	.a(n251075));
   in01s01 U270057 (.o(n185643),
	.a(n251076));
   in01s01 U270058 (.o(n185644),
	.a(n251077));
   in01s01 U270059 (.o(n185645),
	.a(n251078));
   in01s01 U270060 (.o(n185646),
	.a(n251079));
   in01s01 U270061 (.o(n185647),
	.a(n251081));
   oa22s01 U270062 (.o(n251082),
	.a(n251088),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[517]),
	.d(FE_OFN307_n251072));
   in01s01 U270063 (.o(n185648),
	.a(n251082));
   oa22s01 U270064 (.o(n251083),
	.a(n251088),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[516]),
	.d(FE_OFN307_n251072));
   in01s01 U270065 (.o(n185649),
	.a(n251083));
   oa22s01 U270066 (.o(n251084),
	.a(n251088),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[515]),
	.d(FE_OFN307_n251072));
   in01s01 U270067 (.o(n185650),
	.a(n251084));
   oa22s01 U270068 (.o(n251085),
	.a(n251088),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[514]),
	.d(FE_OFN307_n251072));
   in01s01 U270069 (.o(n185651),
	.a(n251085));
   oa22s01 U270070 (.o(n251086),
	.a(n251088),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[513]),
	.d(FE_OFN307_n251072));
   in01s01 U270071 (.o(n185652),
	.a(n251086));
   oa22s01 U270072 (.o(n251089),
	.a(n251088),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[512]),
	.d(FE_OFN306_n251072));
   in01s01 U270073 (.o(n185653),
	.a(n251089));
   in01s01 U270074 (.o(n185654),
	.a(n251090));
   oa22s01 U270075 (.o(n251091),
	.a(n251123),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1534]),
	.d(FE_OFN309_n251105));
   in01s01 U270076 (.o(n185656),
	.a(n251092));
   in01s01 U270077 (.o(n185657),
	.a(n251093));
   in01s01 U270078 (.o(n185658),
	.a(n251094));
   in01s01 U270079 (.o(n185659),
	.a(n251095));
   in01s01 U270080 (.o(n185660),
	.a(n251096));
   in01s01 U270081 (.o(n185661),
	.a(n251097));
   in01s01 U270082 (.o(n185662),
	.a(n251098));
   in01s01 U270083 (.o(n185663),
	.a(n251099));
   in01s01 U270084 (.o(n185664),
	.a(n251100));
   in01s01 U270085 (.o(n185665),
	.a(n251101));
   in01s01 U270086 (.o(n185666),
	.a(n251102));
   in01s01 U270087 (.o(n185667),
	.a(n251103));
   in01s01 U270088 (.o(n185668),
	.a(n251104));
   in01s01 U270089 (.o(n185669),
	.a(n251106));
   oa22s01 U270090 (.o(n251107),
	.a(n251123),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1519]),
	.d(FE_OFN309_n251105));
   in01s01 U270091 (.o(n185671),
	.a(n251108));
   in01s01 U270092 (.o(n185672),
	.a(n251109));
   in01s01 U270093 (.o(n185673),
	.a(n251110));
   in01s01 U270094 (.o(n185674),
	.a(n251111));
   in01s01 U270095 (.o(n185675),
	.a(n251112));
   in01s01 U270096 (.o(n185676),
	.a(n251113));
   in01s01 U270097 (.o(n185677),
	.a(n251114));
   in01s01 U270098 (.o(n185678),
	.a(n251115));
   in01s01 U270099 (.o(n185679),
	.a(n251117));
   oa22s01 U270100 (.o(n251118),
	.a(n251123),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1509]),
	.d(n251105));
   in01s01 U270101 (.o(n185680),
	.a(n251118));
   oa22s01 U270102 (.o(n251119),
	.a(n251123),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1508]),
	.d(FE_OFN309_n251105));
   in01s01 U270103 (.o(n185681),
	.a(n251119));
   oa22s01 U270104 (.o(n251120),
	.a(n251123),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1507]),
	.d(FE_OFN309_n251105));
   in01s01 U270105 (.o(n185682),
	.a(n251120));
   oa22s01 U270106 (.o(n251121),
	.a(n251123),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1506]),
	.d(FE_OFN309_n251105));
   in01s01 U270107 (.o(n185683),
	.a(n251121));
   oa22s01 U270108 (.o(n251122),
	.a(n251123),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1505]),
	.d(FE_OFN309_n251105));
   in01s01 U270109 (.o(n185684),
	.a(n251122));
   oa22s01 U270110 (.o(n251124),
	.a(n251123),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1504]),
	.d(FE_OFN309_n251105));
   in01s01 U270111 (.o(n185686),
	.a(n251125));
   in01s01 U270112 (.o(n185687),
	.a(n251126));
   in01s01 U270113 (.o(n185688),
	.a(n251127));
   in01s01 U270114 (.o(n185689),
	.a(n251128));
   in01s01 U270115 (.o(n185690),
	.a(n251129));
   in01s01 U270116 (.o(n185691),
	.a(n251130));
   in01s01 U270117 (.o(n185692),
	.a(n251131));
   in01s01 U270118 (.o(n185693),
	.a(n251132));
   in01s01 U270119 (.o(n185694),
	.a(n251133));
   in01s01 U270120 (.o(n185695),
	.a(n251134));
   in01s01 U270121 (.o(n185696),
	.a(n251135));
   in01s01 U270122 (.o(n185697),
	.a(n251136));
   in01s01 U270123 (.o(n185698),
	.a(n251137));
   in01s01 U270124 (.o(n185699),
	.a(n251138));
   oa22s01 U270125 (.o(n251139),
	.a(n251158),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1489]),
	.d(FE_OFN420_n251140));
   in01s01 U270126 (.o(n185701),
	.a(n251141));
   in01s01 U270127 (.o(n185702),
	.a(n251142));
   in01s01 U270128 (.o(n185703),
	.a(n251143));
   in01s01 U270129 (.o(n185704),
	.a(n251144));
   in01s01 U270130 (.o(n185705),
	.a(n251145));
   in01s01 U270131 (.o(n185706),
	.a(n251146));
   in01s01 U270132 (.o(n185707),
	.a(n251147));
   in01s01 U270133 (.o(n185708),
	.a(n251148));
   in01s01 U270134 (.o(n185709),
	.a(n251149));
   in01s01 U270135 (.o(n185710),
	.a(n251150));
   in01s01 U270136 (.o(n185711),
	.a(n251152));
   oa22s01 U270137 (.o(n251153),
	.a(n251158),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1477]),
	.d(FE_OFN420_n251140));
   in01s01 U270138 (.o(n185712),
	.a(n251153));
   oa22s01 U270139 (.o(n251154),
	.a(n251158),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1476]),
	.d(FE_OFN420_n251140));
   in01s01 U270140 (.o(n185713),
	.a(n251154));
   oa22s01 U270141 (.o(n251155),
	.a(n251158),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1475]),
	.d(FE_OFN420_n251140));
   in01s01 U270142 (.o(n185714),
	.a(n251155));
   oa22s01 U270143 (.o(n251156),
	.a(n251158),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1474]),
	.d(FE_OFN420_n251140));
   oa22s01 U270144 (.o(n251157),
	.a(n251158),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1473]),
	.d(FE_OFN420_n251140));
   in01s01 U270145 (.o(n185716),
	.a(n251157));
   oa22s01 U270146 (.o(n251159),
	.a(n251158),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1472]),
	.d(FE_OFN420_n251140));
   in01s01 U270147 (.o(n185717),
	.a(n251159));
   in01s01 U270148 (.o(n185718),
	.a(n251160));
   in01s01 U270149 (.o(n185719),
	.a(n251161));
   in01s01 U270150 (.o(n185720),
	.a(n251162));
   in01s01 U270151 (.o(n185721),
	.a(n251163));
   in01s01 U270152 (.o(n185722),
	.a(n251164));
   in01s01 U270153 (.o(n185723),
	.a(n251165));
   in01s01 U270154 (.o(n185724),
	.a(n251166));
   in01s01 U270155 (.o(n185725),
	.a(n251167));
   in01s01 U270156 (.o(n185726),
	.a(n251168));
   in01s01 U270157 (.o(n185727),
	.a(n251169));
   in01s01 U270158 (.o(n185728),
	.a(n251170));
   in01s01 U270159 (.o(n185729),
	.a(n251171));
   oa22s01 U270160 (.o(n251172),
	.a(n251194),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1459]),
	.d(FE_OFN311_n251175));
   in01s01 U270161 (.o(n185731),
	.a(n251173));
   in01s01 U270162 (.o(n185732),
	.a(n251174));
   in01s01 U270163 (.o(n185733),
	.a(n251176));
   in01s01 U270164 (.o(n185734),
	.a(n251177));
   in01s01 U270165 (.o(n185735),
	.a(n251178));
   in01s01 U270166 (.o(n185736),
	.a(n251179));
   in01s01 U270167 (.o(n185737),
	.a(n251180));
   in01s01 U270168 (.o(n185738),
	.a(n251181));
   in01s01 U270169 (.o(n185739),
	.a(n251182));
   in01s01 U270170 (.o(n185740),
	.a(n251183));
   in01s01 U270171 (.o(n185741),
	.a(n251184));
   in01s01 U270172 (.o(n185742),
	.a(n251185));
   in01s01 U270173 (.o(n185743),
	.a(n251187));
   oa22s01 U270174 (.o(n251188),
	.a(n251194),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1445]),
	.d(FE_OFN311_n251175));
   in01s01 U270175 (.o(n185744),
	.a(n251188));
   oa22s01 U270176 (.o(n251189),
	.a(n251194),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1444]),
	.d(FE_OFN311_n251175));
   oa22s01 U270177 (.o(n251190),
	.a(n251194),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1443]),
	.d(FE_OFN311_n251175));
   in01s01 U270178 (.o(n185746),
	.a(n251190));
   oa22s01 U270179 (.o(n251191),
	.a(n251194),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1442]),
	.d(FE_OFN311_n251175));
   in01s01 U270180 (.o(n185747),
	.a(n251191));
   oa22s01 U270181 (.o(n251192),
	.a(n251194),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1441]),
	.d(FE_OFN311_n251175));
   in01s01 U270182 (.o(n185748),
	.a(n251192));
   oa22s01 U270183 (.o(n251195),
	.a(n251194),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1440]),
	.d(FE_OFN311_n251175));
   in01s01 U270184 (.o(n185749),
	.a(n251195));
   oa22s01 U270185 (.o(n251196),
	.a(n251229),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1439]),
	.d(FE_OFN422_n251211));
   in01s01 U270186 (.o(n185750),
	.a(n251196));
   oa22s01 U270187 (.o(n251197),
	.a(n251229),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1438]),
	.d(FE_OFN422_n251211));
   in01s01 U270188 (.o(n185751),
	.a(n251197));
   oa22s01 U270189 (.o(n251198),
	.a(n251229),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1437]),
	.d(FE_OFN422_n251211));
   in01s01 U270190 (.o(n185752),
	.a(n251198));
   oa22s01 U270191 (.o(n251199),
	.a(n251229),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1436]),
	.d(FE_OFN422_n251211));
   in01s01 U270192 (.o(n185753),
	.a(n251199));
   oa22s01 U270193 (.o(n251200),
	.a(n251229),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1435]),
	.d(FE_OFN422_n251211));
   in01s01 U270194 (.o(n185754),
	.a(n251200));
   oa22s01 U270195 (.o(n251201),
	.a(n251229),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1434]),
	.d(FE_OFN422_n251211));
   in01s01 U270196 (.o(n185755),
	.a(n251201));
   oa22s01 U270197 (.o(n251202),
	.a(n251229),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1433]),
	.d(FE_OFN422_n251211));
   in01s01 U270198 (.o(n185756),
	.a(n251202));
   oa22s01 U270199 (.o(n251203),
	.a(n251229),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1432]),
	.d(FE_OFN422_n251211));
   in01s01 U270200 (.o(n185757),
	.a(n251203));
   oa22s01 U270201 (.o(n251204),
	.a(n251229),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1431]),
	.d(FE_OFN422_n251211));
   in01s01 U270202 (.o(n185758),
	.a(n251204));
   oa22s01 U270203 (.o(n251205),
	.a(n251229),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1430]),
	.d(FE_OFN422_n251211));
   in01s01 U270204 (.o(n185759),
	.a(n251205));
   oa22s01 U270205 (.o(n251206),
	.a(n251229),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1429]),
	.d(FE_OFN422_n251211));
   oa22s01 U270206 (.o(n251207),
	.a(n251229),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1428]),
	.d(FE_OFN422_n251211));
   in01s01 U270207 (.o(n185761),
	.a(n251207));
   oa22s01 U270208 (.o(n251208),
	.a(n251229),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1427]),
	.d(FE_OFN422_n251211));
   in01s01 U270209 (.o(n185762),
	.a(n251208));
   oa22s01 U270210 (.o(n251209),
	.a(n251229),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1426]),
	.d(FE_OFN422_n251211));
   in01s01 U270211 (.o(n185763),
	.a(n251209));
   oa22s01 U270212 (.o(n251210),
	.a(n251229),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1425]),
	.d(FE_OFN422_n251211));
   in01s01 U270213 (.o(n185764),
	.a(n251210));
   oa22s01 U270214 (.o(n251212),
	.a(n251229),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1424]),
	.d(FE_OFN422_n251211));
   in01s01 U270215 (.o(n185765),
	.a(n251212));
   oa22s01 U270216 (.o(n251213),
	.a(n251229),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1423]),
	.d(FE_OFN422_n251211));
   in01s01 U270217 (.o(n185766),
	.a(n251213));
   oa22s01 U270218 (.o(n251214),
	.a(n251229),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1422]),
	.d(FE_OFN422_n251211));
   in01s01 U270219 (.o(n185767),
	.a(n251214));
   oa22s01 U270220 (.o(n251215),
	.a(n251229),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1421]),
	.d(FE_OFN422_n251211));
   in01s01 U270221 (.o(n185768),
	.a(n251215));
   oa22s01 U270222 (.o(n251216),
	.a(n251229),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1420]),
	.d(FE_OFN422_n251211));
   in01s01 U270223 (.o(n185769),
	.a(n251216));
   oa22s01 U270224 (.o(n251217),
	.a(n251229),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1419]),
	.d(FE_OFN422_n251211));
   in01s01 U270225 (.o(n185770),
	.a(n251217));
   oa22s01 U270226 (.o(n251218),
	.a(n251229),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1418]),
	.d(FE_OFN422_n251211));
   in01s01 U270227 (.o(n185771),
	.a(n251218));
   oa22s01 U270228 (.o(n251219),
	.a(n251229),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1417]),
	.d(FE_OFN422_n251211));
   in01s01 U270229 (.o(n185772),
	.a(n251219));
   oa22s01 U270230 (.o(n251220),
	.a(n251229),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1416]),
	.d(FE_OFN422_n251211));
   in01s01 U270231 (.o(n185773),
	.a(n251220));
   oa22s01 U270232 (.o(n251221),
	.a(n251229),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1415]),
	.d(FE_OFN422_n251211));
   in01s01 U270233 (.o(n185774),
	.a(n251221));
   oa22s01 U270234 (.o(n251223),
	.a(n251229),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1414]),
	.d(FE_OFN422_n251211));
   oa22s01 U270235 (.o(n251224),
	.a(n251229),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1413]),
	.d(FE_OFN422_n251211));
   in01s01 U270236 (.o(n185776),
	.a(n251224));
   oa22s01 U270237 (.o(n251225),
	.a(n251229),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1412]),
	.d(FE_OFN422_n251211));
   in01s01 U270238 (.o(n185777),
	.a(n251225));
   oa22s01 U270239 (.o(n251226),
	.a(n251229),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1411]),
	.d(FE_OFN422_n251211));
   in01s01 U270240 (.o(n185778),
	.a(n251226));
   oa22s01 U270241 (.o(n251227),
	.a(n251229),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1410]),
	.d(FE_OFN422_n251211));
   in01s01 U270242 (.o(n185779),
	.a(n251227));
   oa22s01 U270243 (.o(n251228),
	.a(n251229),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1409]),
	.d(FE_OFN422_n251211));
   in01s01 U270244 (.o(n185780),
	.a(n251228));
   oa22s01 U270245 (.o(n251230),
	.a(n251229),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1408]),
	.d(FE_OFN422_n251211));
   in01s01 U270246 (.o(n185781),
	.a(n251230));
   in01s01 U270247 (.o(n185782),
	.a(n251231));
   in01s01 U270248 (.o(n185783),
	.a(n251232));
   in01s01 U270249 (.o(n185784),
	.a(n251233));
   in01s01 U270250 (.o(n185785),
	.a(n251234));
   in01s01 U270251 (.o(n185786),
	.a(n251235));
   in01s01 U270252 (.o(n185787),
	.a(n251236));
   in01s01 U270253 (.o(n185788),
	.a(n251237));
   in01s01 U270254 (.o(n185789),
	.a(n251238));
   oa22s01 U270255 (.o(n251239),
	.a(n251264),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1399]),
	.d(FE_OFN202_n251246));
   in01s01 U270256 (.o(n185791),
	.a(n251240));
   in01s01 U270257 (.o(n185792),
	.a(n251241));
   in01s01 U270258 (.o(n185793),
	.a(n251242));
   in01s01 U270259 (.o(n185794),
	.a(n251243));
   in01s01 U270260 (.o(n185795),
	.a(n251244));
   in01s01 U270261 (.o(n185796),
	.a(n251245));
   in01s01 U270262 (.o(n185797),
	.a(n251247));
   in01s01 U270263 (.o(n185798),
	.a(n251248));
   in01s01 U270264 (.o(n185799),
	.a(n251249));
   in01s01 U270265 (.o(n185800),
	.a(n251250));
   in01s01 U270266 (.o(n185801),
	.a(n251251));
   in01s01 U270267 (.o(n185802),
	.a(n251252));
   in01s01 U270268 (.o(n185803),
	.a(n251253));
   in01s01 U270269 (.o(n185804),
	.a(n251254));
   oa22s01 U270270 (.o(n251255),
	.a(n251264),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1384]),
	.d(FE_OFN202_n251246));
   in01s01 U270271 (.o(n185806),
	.a(n251256));
   in01s01 U270272 (.o(n185807),
	.a(n251258));
   oa22s01 U270273 (.o(n251259),
	.a(n251264),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1381]),
	.d(FE_OFN202_n251246));
   in01s01 U270274 (.o(n185808),
	.a(n251259));
   oa22s01 U270275 (.o(n251260),
	.a(n251264),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1380]),
	.d(FE_OFN202_n251246));
   in01s01 U270276 (.o(n185809),
	.a(n251260));
   oa22s01 U270277 (.o(n251261),
	.a(n251264),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1379]),
	.d(FE_OFN202_n251246));
   in01s01 U270278 (.o(n185810),
	.a(n251261));
   oa22s01 U270279 (.o(n251262),
	.a(n251264),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1378]),
	.d(FE_OFN202_n251246));
   in01s01 U270280 (.o(n185811),
	.a(n251262));
   oa22s01 U270281 (.o(n251263),
	.a(n251264),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1377]),
	.d(FE_OFN202_n251246));
   in01s01 U270282 (.o(n185812),
	.a(n251263));
   oa22s01 U270283 (.o(n251265),
	.a(n251264),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1376]),
	.d(FE_OFN202_n251246));
   in01s01 U270284 (.o(n185813),
	.a(n251265));
   oa22s01 U270285 (.o(n251266),
	.a(n251300),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1375]),
	.d(FE_OFN314_n251281));
   in01s01 U270286 (.o(n185814),
	.a(n251266));
   oa22s01 U270287 (.o(n251267),
	.a(n251300),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1374]),
	.d(FE_OFN314_n251281));
   in01s01 U270288 (.o(n185815),
	.a(n251267));
   oa22s01 U270289 (.o(n251268),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1373]),
	.d(FE_OFN313_n251281));
   in01s01 U270290 (.o(n185816),
	.a(n251268));
   oa22s01 U270291 (.o(n251269),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1372]),
	.d(FE_OFN313_n251281));
   in01s01 U270292 (.o(n185817),
	.a(n251269));
   oa22s01 U270293 (.o(n251270),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1371]),
	.d(FE_OFN313_n251281));
   in01s01 U270294 (.o(n185818),
	.a(n251270));
   oa22s01 U270295 (.o(n251271),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1370]),
	.d(FE_OFN314_n251281));
   in01s01 U270296 (.o(n185819),
	.a(n251271));
   oa22s01 U270297 (.o(n251272),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1369]),
	.d(FE_OFN314_n251281));
   oa22s01 U270298 (.o(n251273),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1368]),
	.d(FE_OFN313_n251281));
   in01s01 U270299 (.o(n185821),
	.a(n251273));
   oa22s01 U270300 (.o(n251274),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1367]),
	.d(FE_OFN313_n251281));
   in01s01 U270301 (.o(n185822),
	.a(n251274));
   oa22s01 U270302 (.o(n251275),
	.a(n251300),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1366]),
	.d(FE_OFN314_n251281));
   in01s01 U270303 (.o(n185823),
	.a(n251275));
   oa22s01 U270304 (.o(n251276),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1365]),
	.d(FE_OFN314_n251281));
   in01s01 U270305 (.o(n185824),
	.a(n251276));
   oa22s01 U270306 (.o(n251277),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1364]),
	.d(FE_OFN314_n251281));
   in01s01 U270307 (.o(n185825),
	.a(n251277));
   oa22s01 U270308 (.o(n251278),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1363]),
	.d(FE_OFN314_n251281));
   in01s01 U270309 (.o(n185826),
	.a(n251278));
   oa22s01 U270310 (.o(n251279),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1362]),
	.d(FE_OFN314_n251281));
   in01s01 U270311 (.o(n185827),
	.a(n251279));
   oa22s01 U270312 (.o(n251280),
	.a(n251300),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1361]),
	.d(FE_OFN314_n251281));
   in01s01 U270313 (.o(n185828),
	.a(n251280));
   oa22s01 U270314 (.o(n251282),
	.a(n251300),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1360]),
	.d(FE_OFN314_n251281));
   in01s01 U270315 (.o(n185829),
	.a(n251282));
   oa22s01 U270316 (.o(n251283),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1359]),
	.d(FE_OFN313_n251281));
   in01s01 U270317 (.o(n185830),
	.a(n251283));
   oa22s01 U270318 (.o(n251284),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1358]),
	.d(FE_OFN313_n251281));
   in01s01 U270319 (.o(n185831),
	.a(n251284));
   oa22s01 U270320 (.o(n251285),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1357]),
	.d(FE_OFN313_n251281));
   in01s01 U270321 (.o(n185832),
	.a(n251285));
   oa22s01 U270322 (.o(n251286),
	.a(n251300),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1356]),
	.d(FE_OFN314_n251281));
   in01s01 U270323 (.o(n185833),
	.a(n251286));
   oa22s01 U270324 (.o(n251287),
	.a(n251300),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1355]),
	.d(FE_OFN314_n251281));
   in01s01 U270325 (.o(n185834),
	.a(n251287));
   oa22s01 U270326 (.o(n251288),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1354]),
	.d(FE_OFN313_n251281));
   oa22s01 U270327 (.o(n251289),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1353]),
	.d(FE_OFN313_n251281));
   in01s01 U270328 (.o(n185836),
	.a(n251289));
   oa22s01 U270329 (.o(n251290),
	.a(n251300),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1352]),
	.d(FE_OFN314_n251281));
   in01s01 U270330 (.o(n185837),
	.a(n251290));
   oa22s01 U270331 (.o(n251291),
	.a(n251300),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1351]),
	.d(FE_OFN314_n251281));
   in01s01 U270332 (.o(n185838),
	.a(n251291));
   oa22s01 U270333 (.o(n251293),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1350]),
	.d(FE_OFN313_n251281));
   in01s01 U270334 (.o(n185839),
	.a(n251293));
   oa22s01 U270335 (.o(n251294),
	.a(n251300),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1349]),
	.d(FE_OFN314_n251281));
   in01s01 U270336 (.o(n185840),
	.a(n251294));
   oa22s01 U270337 (.o(n251295),
	.a(n251300),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1348]),
	.d(FE_OFN314_n251281));
   in01s01 U270338 (.o(n185841),
	.a(n251295));
   oa22s01 U270339 (.o(n251296),
	.a(n251300),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1347]),
	.d(FE_OFN314_n251281));
   in01s01 U270340 (.o(n185842),
	.a(n251296));
   oa22s01 U270341 (.o(n251297),
	.a(n251300),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1346]),
	.d(FE_OFN314_n251281));
   in01s01 U270342 (.o(n185843),
	.a(n251297));
   oa22s01 U270343 (.o(n251298),
	.a(n251300),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1345]),
	.d(FE_OFN314_n251281));
   in01s01 U270344 (.o(n185844),
	.a(n251298));
   oa22s01 U270345 (.o(n251301),
	.a(FE_OFN424_n251300),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1344]),
	.d(FE_OFN313_n251281));
   in01s01 U270346 (.o(n185845),
	.a(n251301));
   in01s01 U270347 (.o(n185846),
	.a(n251302));
   in01s01 U270348 (.o(n185847),
	.a(n251303));
   in01s01 U270349 (.o(n185848),
	.a(n251304));
   in01s01 U270350 (.o(n185849),
	.a(n251305));
   oa22s01 U270351 (.o(n251306),
	.a(n251335),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1339]),
	.d(FE_OFN316_n251317));
   in01s01 U270352 (.o(n185851),
	.a(n251307));
   in01s01 U270353 (.o(n185852),
	.a(n251308));
   in01s01 U270354 (.o(n185853),
	.a(n251309));
   in01s01 U270355 (.o(n185854),
	.a(n251310));
   in01s01 U270356 (.o(n185855),
	.a(n251311));
   in01s01 U270357 (.o(n185856),
	.a(n251312));
   in01s01 U270358 (.o(n185857),
	.a(n251313));
   in01s01 U270359 (.o(n185858),
	.a(n251314));
   in01s01 U270360 (.o(n185859),
	.a(n251315));
   in01s01 U270361 (.o(n185860),
	.a(n251316));
   in01s01 U270362 (.o(n185861),
	.a(n251318));
   in01s01 U270363 (.o(n185862),
	.a(n251319));
   in01s01 U270364 (.o(n185863),
	.a(n251320));
   in01s01 U270365 (.o(n185864),
	.a(n251321));
   oa22s01 U270366 (.o(n251322),
	.a(n251335),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1324]),
	.d(FE_OFN316_n251317));
   in01s01 U270367 (.o(n185866),
	.a(n251323));
   in01s01 U270368 (.o(n185867),
	.a(n251324));
   in01s01 U270369 (.o(n185868),
	.a(n251325));
   in01s01 U270370 (.o(n185869),
	.a(n251326));
   in01s01 U270371 (.o(n185870),
	.a(n251327));
   in01s01 U270372 (.o(n185871),
	.a(n251329));
   oa22s01 U270373 (.o(n251330),
	.a(n251335),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1317]),
	.d(FE_OFN316_n251317));
   in01s01 U270374 (.o(n185872),
	.a(n251330));
   oa22s01 U270375 (.o(n251331),
	.a(n251335),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1316]),
	.d(FE_OFN316_n251317));
   in01s01 U270376 (.o(n185873),
	.a(n251331));
   oa22s01 U270377 (.o(n251332),
	.a(n251335),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1315]),
	.d(FE_OFN316_n251317));
   in01s01 U270378 (.o(n185874),
	.a(n251332));
   oa22s01 U270379 (.o(n251333),
	.a(n251335),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1314]),
	.d(FE_OFN316_n251317));
   in01s01 U270380 (.o(n185875),
	.a(n251333));
   oa22s01 U270381 (.o(n251334),
	.a(n251335),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1313]),
	.d(FE_OFN316_n251317));
   in01s01 U270382 (.o(n185876),
	.a(n251334));
   oa22s01 U270383 (.o(n251336),
	.a(n251335),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1312]),
	.d(FE_OFN316_n251317));
   in01s01 U270384 (.o(n185877),
	.a(n251336));
   in01s01 U270385 (.o(n185878),
	.a(n251338));
   in01s01 U270386 (.o(n185879),
	.a(n251339));
   oa22s01 U270387 (.o(n251340),
	.a(n251371),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1309]),
	.d(FE_OFN318_n251353));
   in01s01 U270388 (.o(n185881),
	.a(n251341));
   in01s01 U270389 (.o(n185882),
	.a(n251342));
   in01s01 U270390 (.o(n185883),
	.a(n251343));
   in01s01 U270391 (.o(n185884),
	.a(n251344));
   in01s01 U270392 (.o(n185885),
	.a(n251345));
   in01s01 U270393 (.o(n185886),
	.a(n251346));
   in01s01 U270394 (.o(n185887),
	.a(n251347));
   in01s01 U270395 (.o(n185888),
	.a(n251348));
   in01s01 U270396 (.o(n185889),
	.a(n251349));
   in01s01 U270397 (.o(n185890),
	.a(n251350));
   in01s01 U270398 (.o(n185891),
	.a(n251351));
   in01s01 U270399 (.o(n185892),
	.a(n251352));
   in01s01 U270400 (.o(n185893),
	.a(n251354));
   in01s01 U270401 (.o(n185894),
	.a(n251355));
   oa22s01 U270402 (.o(n251356),
	.a(n251371),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1294]),
	.d(FE_OFN318_n251353));
   in01s01 U270403 (.o(n185896),
	.a(n251357));
   in01s01 U270404 (.o(n185897),
	.a(n251358));
   in01s01 U270405 (.o(n185898),
	.a(n251359));
   in01s01 U270406 (.o(n185899),
	.a(n251360));
   in01s01 U270407 (.o(n185900),
	.a(n251361));
   in01s01 U270408 (.o(n185901),
	.a(n251362));
   in01s01 U270409 (.o(n185902),
	.a(n251363));
   in01s01 U270410 (.o(n185903),
	.a(n251365));
   oa22s01 U270411 (.o(n251366),
	.a(n251371),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1285]),
	.d(FE_OFN318_n251353));
   in01s01 U270412 (.o(n185904),
	.a(n251366));
   oa22s01 U270413 (.o(n251367),
	.a(n251371),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1284]),
	.d(FE_OFN318_n251353));
   in01s01 U270414 (.o(n185905),
	.a(n251367));
   oa22s01 U270415 (.o(n251368),
	.a(n251371),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1283]),
	.d(FE_OFN318_n251353));
   in01s01 U270416 (.o(n185906),
	.a(n251368));
   oa22s01 U270417 (.o(n251369),
	.a(n251371),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1282]),
	.d(FE_OFN318_n251353));
   in01s01 U270418 (.o(n185907),
	.a(n251369));
   oa22s01 U270419 (.o(n251370),
	.a(n251371),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1281]),
	.d(FE_OFN318_n251353));
   in01s01 U270420 (.o(n185908),
	.a(n251370));
   oa22s01 U270421 (.o(n251372),
	.a(n251371),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1280]),
	.d(FE_OFN318_n251353));
   in01s01 U270422 (.o(n185909),
	.a(n251372));
   oa22s01 U270423 (.o(n251373),
	.a(n251407),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1279]),
	.d(FE_OFN320_n251388));
   in01s01 U270424 (.o(n185911),
	.a(n251374));
   in01s01 U270425 (.o(n185912),
	.a(n251375));
   in01s01 U270426 (.o(n185913),
	.a(n251376));
   in01s01 U270427 (.o(n185914),
	.a(n251377));
   in01s01 U270428 (.o(n185915),
	.a(n251378));
   in01s01 U270429 (.o(n185916),
	.a(n251379));
   in01s01 U270430 (.o(n185917),
	.a(n251380));
   in01s01 U270431 (.o(n185918),
	.a(n251381));
   in01s01 U270432 (.o(n185919),
	.a(n251382));
   in01s01 U270433 (.o(n185920),
	.a(n251383));
   in01s01 U270434 (.o(n185921),
	.a(n251384));
   in01s01 U270435 (.o(n185922),
	.a(n251385));
   in01s01 U270436 (.o(n185923),
	.a(n251386));
   in01s01 U270437 (.o(n185924),
	.a(n251387));
   oa22s01 U270438 (.o(n251389),
	.a(n251407),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1264]),
	.d(FE_OFN320_n251388));
   in01s01 U270439 (.o(n185926),
	.a(n251390));
   in01s01 U270440 (.o(n185927),
	.a(n251391));
   in01s01 U270441 (.o(n185928),
	.a(n251392));
   in01s01 U270442 (.o(n185929),
	.a(n251393));
   in01s01 U270443 (.o(n185930),
	.a(n251394));
   in01s01 U270444 (.o(n185931),
	.a(n251395));
   in01s01 U270445 (.o(n185932),
	.a(n251396));
   in01s01 U270446 (.o(n185933),
	.a(n251397));
   in01s01 U270447 (.o(n185934),
	.a(n251398));
   in01s01 U270448 (.o(n185935),
	.a(n251400));
   oa22s01 U270449 (.o(n251401),
	.a(n251407),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1253]),
	.d(FE_OFN320_n251388));
   in01s01 U270450 (.o(n185936),
	.a(n251401));
   oa22s01 U270451 (.o(n251402),
	.a(n251407),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1252]),
	.d(FE_OFN320_n251388));
   in01s01 U270452 (.o(n185937),
	.a(n251402));
   oa22s01 U270453 (.o(n251403),
	.a(n251407),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1251]),
	.d(FE_OFN320_n251388));
   in01s01 U270454 (.o(n185938),
	.a(n251403));
   oa22s01 U270455 (.o(n251404),
	.a(n251407),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1250]),
	.d(FE_OFN320_n251388));
   in01s01 U270456 (.o(n185939),
	.a(n251404));
   oa22s01 U270457 (.o(n251405),
	.a(n251407),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1249]),
	.d(FE_OFN320_n251388));
   oa22s01 U270458 (.o(n251408),
	.a(n251407),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1248]),
	.d(FE_OFN320_n251388));
   in01s01 U270459 (.o(n185941),
	.a(n251408));
   in01s01 U270460 (.o(n185942),
	.a(n251409));
   in01s01 U270461 (.o(n185943),
	.a(n251410));
   in01s01 U270462 (.o(n185944),
	.a(n251411));
   in01s01 U270463 (.o(n185945),
	.a(n251412));
   in01s01 U270464 (.o(n185946),
	.a(n251413));
   in01s01 U270465 (.o(n185947),
	.a(n251414));
   in01s01 U270466 (.o(n185948),
	.a(n251415));
   in01s01 U270467 (.o(n185949),
	.a(n251416));
   in01s01 U270468 (.o(n185950),
	.a(n251417));
   in01s01 U270469 (.o(n185951),
	.a(n251418));
   in01s01 U270470 (.o(n185952),
	.a(n251419));
   in01s01 U270471 (.o(n185953),
	.a(n251420));
   in01s01 U270472 (.o(n185954),
	.a(n251421));
   oa22s01 U270473 (.o(n251422),
	.a(n251442),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1234]),
	.d(FE_OFN426_n251424));
   in01s01 U270474 (.o(n185956),
	.a(n251423));
   in01s01 U270475 (.o(n185957),
	.a(n251425));
   in01s01 U270476 (.o(n185958),
	.a(n251426));
   in01s01 U270477 (.o(n185959),
	.a(n251427));
   in01s01 U270478 (.o(n185960),
	.a(n251428));
   in01s01 U270479 (.o(n185961),
	.a(n251429));
   in01s01 U270480 (.o(n185962),
	.a(n251430));
   in01s01 U270481 (.o(n185963),
	.a(n251431));
   in01s01 U270482 (.o(n185964),
	.a(n251432));
   in01s01 U270483 (.o(n185965),
	.a(n251433));
   in01s01 U270484 (.o(n185966),
	.a(n251434));
   in01s01 U270485 (.o(n185967),
	.a(n251436));
   oa22s01 U270486 (.o(n251437),
	.a(n251442),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1221]),
	.d(FE_OFN426_n251424));
   in01s01 U270487 (.o(n185968),
	.a(n251437));
   oa22s01 U270488 (.o(n251438),
	.a(n251442),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1220]),
	.d(FE_OFN426_n251424));
   in01s01 U270489 (.o(n185969),
	.a(n251438));
   oa22s01 U270490 (.o(n251439),
	.a(n251442),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1219]),
	.d(FE_OFN426_n251424));
   oa22s01 U270491 (.o(n251440),
	.a(n251442),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1218]),
	.d(FE_OFN426_n251424));
   in01s01 U270492 (.o(n185971),
	.a(n251440));
   oa22s01 U270493 (.o(n251441),
	.a(n251442),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1217]),
	.d(FE_OFN426_n251424));
   in01s01 U270494 (.o(n185972),
	.a(n251441));
   oa22s01 U270495 (.o(n251443),
	.a(n251442),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1216]),
	.d(FE_OFN426_n251424));
   in01s01 U270496 (.o(n185973),
	.a(n251443));
   in01s01 U270497 (.o(n185974),
	.a(n251444));
   in01s01 U270498 (.o(n185975),
	.a(n251445));
   in01s01 U270499 (.o(n185976),
	.a(n251446));
   in01s01 U270500 (.o(n185977),
	.a(n251447));
   in01s01 U270501 (.o(n185978),
	.a(n251448));
   in01s01 U270502 (.o(n185979),
	.a(n251449));
   in01s01 U270503 (.o(n185980),
	.a(n251450));
   in01s01 U270504 (.o(n185981),
	.a(n251451));
   in01s01 U270505 (.o(n185982),
	.a(n251452));
   in01s01 U270506 (.o(n185983),
	.a(n251453));
   in01s01 U270507 (.o(n185984),
	.a(n251454));
   oa22s01 U270508 (.o(n251455),
	.a(n251477),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1204]),
	.d(FE_OFN322_n251459));
   in01s01 U270509 (.o(n185986),
	.a(n251456));
   in01s01 U270510 (.o(n185987),
	.a(n251457));
   in01s01 U270511 (.o(n185988),
	.a(n251458));
   in01s01 U270512 (.o(n185989),
	.a(n251460));
   in01s01 U270513 (.o(n185990),
	.a(n251461));
   in01s01 U270514 (.o(n185991),
	.a(n251462));
   in01s01 U270515 (.o(n185992),
	.a(n251463));
   in01s01 U270516 (.o(n185993),
	.a(n251464));
   in01s01 U270517 (.o(n185994),
	.a(n251465));
   in01s01 U270518 (.o(n185995),
	.a(n251466));
   in01s01 U270519 (.o(n185996),
	.a(n251467));
   in01s01 U270520 (.o(n185997),
	.a(n251468));
   in01s01 U270521 (.o(n185998),
	.a(n251469));
   in01s01 U270522 (.o(n185999),
	.a(n251471));
   oa22s01 U270523 (.o(n251472),
	.a(n251477),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1189]),
	.d(FE_OFN322_n251459));
   oa22s01 U270524 (.o(n251473),
	.a(n251477),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1188]),
	.d(FE_OFN322_n251459));
   in01s01 U270525 (.o(n186001),
	.a(n251473));
   oa22s01 U270526 (.o(n251474),
	.a(n251477),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1187]),
	.d(FE_OFN322_n251459));
   in01s01 U270527 (.o(n186002),
	.a(n251474));
   oa22s01 U270528 (.o(n251475),
	.a(n251477),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1186]),
	.d(FE_OFN322_n251459));
   in01s01 U270529 (.o(n186003),
	.a(n251475));
   oa22s01 U270530 (.o(n251476),
	.a(n251477),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1185]),
	.d(FE_OFN322_n251459));
   in01s01 U270531 (.o(n186004),
	.a(n251476));
   oa22s01 U270532 (.o(n251478),
	.a(n251477),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1184]),
	.d(FE_OFN322_n251459));
   in01s01 U270533 (.o(n186005),
	.a(n251478));
   oa22s01 U270534 (.o(n251479),
	.a(n251513),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1183]),
	.d(FE_OFN428_n251494));
   in01s01 U270535 (.o(n186006),
	.a(n251479));
   oa22s01 U270536 (.o(n251480),
	.a(n251513),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1182]),
	.d(FE_OFN428_n251494));
   in01s01 U270537 (.o(n186007),
	.a(n251480));
   oa22s01 U270538 (.o(n251481),
	.a(n251513),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1181]),
	.d(FE_OFN428_n251494));
   in01s01 U270539 (.o(n186008),
	.a(n251481));
   oa22s01 U270540 (.o(n251482),
	.a(n251513),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1180]),
	.d(FE_OFN428_n251494));
   in01s01 U270541 (.o(n186009),
	.a(n251482));
   oa22s01 U270542 (.o(n251483),
	.a(n251513),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1179]),
	.d(FE_OFN428_n251494));
   in01s01 U270543 (.o(n186010),
	.a(n251483));
   oa22s01 U270544 (.o(n251484),
	.a(n251513),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1178]),
	.d(FE_OFN428_n251494));
   in01s01 U270545 (.o(n186011),
	.a(n251484));
   oa22s01 U270546 (.o(n251485),
	.a(n251513),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1177]),
	.d(FE_OFN428_n251494));
   in01s01 U270547 (.o(n186012),
	.a(n251485));
   oa22s01 U270548 (.o(n251486),
	.a(n251513),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1176]),
	.d(FE_OFN428_n251494));
   in01s01 U270549 (.o(n186013),
	.a(n251486));
   oa22s01 U270550 (.o(n251487),
	.a(n251513),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1175]),
	.d(FE_OFN428_n251494));
   in01s01 U270551 (.o(n186014),
	.a(n251487));
   oa22s01 U270552 (.o(n251488),
	.a(n251513),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1174]),
	.d(FE_OFN428_n251494));
   oa22s01 U270553 (.o(n251489),
	.a(n251513),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1173]),
	.d(FE_OFN428_n251494));
   in01s01 U270554 (.o(n186016),
	.a(n251489));
   oa22s01 U270555 (.o(n251490),
	.a(n251513),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1172]),
	.d(FE_OFN428_n251494));
   in01s01 U270556 (.o(n186017),
	.a(n251490));
   oa22s01 U270557 (.o(n251491),
	.a(n251513),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1171]),
	.d(FE_OFN428_n251494));
   in01s01 U270558 (.o(n186018),
	.a(n251491));
   oa22s01 U270559 (.o(n251492),
	.a(n251513),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1170]),
	.d(FE_OFN428_n251494));
   in01s01 U270560 (.o(n186019),
	.a(n251492));
   oa22s01 U270561 (.o(n251493),
	.a(n251513),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1169]),
	.d(FE_OFN428_n251494));
   in01s01 U270562 (.o(n186020),
	.a(n251493));
   oa22s01 U270563 (.o(n251495),
	.a(n251513),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1168]),
	.d(FE_OFN428_n251494));
   in01s01 U270564 (.o(n186021),
	.a(n251495));
   oa22s01 U270565 (.o(n251496),
	.a(n251513),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1167]),
	.d(FE_OFN428_n251494));
   in01s01 U270566 (.o(n186022),
	.a(n251496));
   oa22s01 U270567 (.o(n251497),
	.a(n251513),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1166]),
	.d(FE_OFN428_n251494));
   in01s01 U270568 (.o(n186023),
	.a(n251497));
   oa22s01 U270569 (.o(n251498),
	.a(n251513),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1165]),
	.d(FE_OFN428_n251494));
   in01s01 U270570 (.o(n186024),
	.a(n251498));
   oa22s01 U270571 (.o(n251499),
	.a(n251513),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1164]),
	.d(FE_OFN428_n251494));
   in01s01 U270572 (.o(n186025),
	.a(n251499));
   oa22s01 U270573 (.o(n251500),
	.a(n251513),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1163]),
	.d(FE_OFN428_n251494));
   in01s01 U270574 (.o(n186026),
	.a(n251500));
   oa22s01 U270575 (.o(n251501),
	.a(n251513),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1162]),
	.d(FE_OFN428_n251494));
   in01s01 U270576 (.o(n186027),
	.a(n251501));
   oa22s01 U270577 (.o(n251502),
	.a(n251513),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1161]),
	.d(FE_OFN428_n251494));
   in01s01 U270578 (.o(n186028),
	.a(n251502));
   oa22s01 U270579 (.o(n251503),
	.a(n251513),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1160]),
	.d(FE_OFN428_n251494));
   in01s01 U270580 (.o(n186029),
	.a(n251503));
   oa22s01 U270581 (.o(n251504),
	.a(n251513),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1159]),
	.d(FE_OFN428_n251494));
   oa22s01 U270582 (.o(n251506),
	.a(n251513),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1158]),
	.d(FE_OFN428_n251494));
   in01s01 U270583 (.o(n186031),
	.a(n251506));
   oa22s01 U270584 (.o(n251507),
	.a(n251513),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1157]),
	.d(FE_OFN428_n251494));
   in01s01 U270585 (.o(n186032),
	.a(n251507));
   oa22s01 U270586 (.o(n251508),
	.a(n251513),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1156]),
	.d(FE_OFN428_n251494));
   in01s01 U270587 (.o(n186033),
	.a(n251508));
   oa22s01 U270588 (.o(n251509),
	.a(n251513),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1155]),
	.d(FE_OFN428_n251494));
   in01s01 U270589 (.o(n186034),
	.a(n251509));
   oa22s01 U270590 (.o(n251510),
	.a(n251513),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1154]),
	.d(FE_OFN428_n251494));
   in01s01 U270591 (.o(n186035),
	.a(n251510));
   oa22s01 U270592 (.o(n251511),
	.a(n251513),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1153]),
	.d(FE_OFN428_n251494));
   in01s01 U270593 (.o(n186036),
	.a(n251511));
   oa22s01 U270594 (.o(n251514),
	.a(n251513),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1152]),
	.d(FE_OFN428_n251494));
   in01s01 U270595 (.o(n186037),
	.a(n251514));
   in01s01 U270596 (.o(n186038),
	.a(n251515));
   in01s01 U270597 (.o(n186039),
	.a(n251516));
   in01s01 U270598 (.o(n186040),
	.a(n251517));
   in01s01 U270599 (.o(n186041),
	.a(n251518));
   in01s01 U270600 (.o(n186042),
	.a(n251519));
   in01s01 U270601 (.o(n186043),
	.a(n251520));
   in01s01 U270602 (.o(n186044),
	.a(n251521));
   oa22s01 U270603 (.o(n251522),
	.a(n251548),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1144]),
	.d(FE_OFN204_n251530));
   in01s01 U270604 (.o(n186046),
	.a(n251523));
   in01s01 U270605 (.o(n186047),
	.a(n251524));
   in01s01 U270606 (.o(n186048),
	.a(n251525));
   in01s01 U270607 (.o(n186049),
	.a(n251526));
   in01s01 U270608 (.o(n186050),
	.a(n251527));
   in01s01 U270609 (.o(n186051),
	.a(n251528));
   in01s01 U270610 (.o(n186052),
	.a(n251529));
   in01s01 U270611 (.o(n186053),
	.a(n251531));
   in01s01 U270612 (.o(n186054),
	.a(n251532));
   in01s01 U270613 (.o(n186055),
	.a(n251533));
   in01s01 U270614 (.o(n186056),
	.a(n251534));
   in01s01 U270615 (.o(n186057),
	.a(n251535));
   in01s01 U270616 (.o(n186058),
	.a(n251536));
   in01s01 U270617 (.o(n186059),
	.a(n251537));
   oa22s01 U270618 (.o(n251538),
	.a(n251548),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1129]),
	.d(FE_OFN204_n251530));
   in01s01 U270619 (.o(n186061),
	.a(n251539));
   in01s01 U270620 (.o(n186062),
	.a(n251540));
   in01s01 U270621 (.o(n186063),
	.a(n251542));
   oa22s01 U270622 (.o(n251543),
	.a(n251548),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1125]),
	.d(FE_OFN204_n251530));
   in01s01 U270623 (.o(n186064),
	.a(n251543));
   oa22s01 U270624 (.o(n251544),
	.a(n251548),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1124]),
	.d(FE_OFN204_n251530));
   in01s01 U270625 (.o(n186065),
	.a(n251544));
   oa22s01 U270626 (.o(n251545),
	.a(n251548),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1123]),
	.d(FE_OFN204_n251530));
   in01s01 U270627 (.o(n186066),
	.a(n251545));
   oa22s01 U270628 (.o(n251546),
	.a(n251548),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1122]),
	.d(FE_OFN204_n251530));
   in01s01 U270629 (.o(n186067),
	.a(n251546));
   oa22s01 U270630 (.o(n251547),
	.a(n251548),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1121]),
	.d(FE_OFN204_n251530));
   in01s01 U270631 (.o(n186068),
	.a(n251547));
   oa22s01 U270632 (.o(n251549),
	.a(n251548),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1120]),
	.d(FE_OFN204_n251530));
   in01s01 U270633 (.o(n186069),
	.a(n251549));
   oa22s01 U270634 (.o(n251550),
	.a(n251583),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1119]),
	.d(FE_OFN325_n251565));
   in01s01 U270635 (.o(n186070),
	.a(n251550));
   oa22s01 U270636 (.o(n251551),
	.a(n251583),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1118]),
	.d(FE_OFN325_n251565));
   in01s01 U270637 (.o(n186071),
	.a(n251551));
   oa22s01 U270638 (.o(n251552),
	.a(n251583),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1117]),
	.d(FE_OFN324_n251565));
   in01s01 U270639 (.o(n186072),
	.a(n251552));
   oa22s01 U270640 (.o(n251553),
	.a(n251583),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1116]),
	.d(FE_OFN324_n251565));
   in01s01 U270641 (.o(n186073),
	.a(n251553));
   oa22s01 U270642 (.o(n251554),
	.a(n251583),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1115]),
	.d(FE_OFN324_n251565));
   in01s01 U270643 (.o(n186074),
	.a(n251554));
   oa22s01 U270644 (.o(n251555),
	.a(n251583),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1114]),
	.d(FE_OFN325_n251565));
   oa22s01 U270645 (.o(n251556),
	.a(n251583),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1113]),
	.d(FE_OFN325_n251565));
   in01s01 U270646 (.o(n186076),
	.a(n251556));
   in01s01 U270647 (.o(n186077),
	.a(n251557));
   oa22s01 U270648 (.o(n251558),
	.a(n251583),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1111]),
	.d(FE_OFN324_n251565));
   in01s01 U270649 (.o(n186078),
	.a(n251558));
   in01s01 U270650 (.o(n186079),
	.a(n251559));
   oa22s01 U270651 (.o(n251560),
	.a(n251583),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1109]),
	.d(FE_OFN325_n251565));
   in01s01 U270652 (.o(n186080),
	.a(n251560));
   in01s01 U270653 (.o(n186081),
	.a(n251561));
   oa22s01 U270654 (.o(n251562),
	.a(n251583),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1107]),
	.d(FE_OFN325_n251565));
   in01s01 U270655 (.o(n186082),
	.a(n251562));
   in01s01 U270656 (.o(n186083),
	.a(n251563));
   oa22s01 U270657 (.o(n251564),
	.a(n251583),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1105]),
	.d(FE_OFN325_n251565));
   in01s01 U270658 (.o(n186084),
	.a(n251564));
   oa22s01 U270659 (.o(n251566),
	.a(n251583),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1104]),
	.d(FE_OFN325_n251565));
   in01s01 U270660 (.o(n186085),
	.a(n251566));
   in01s01 U270661 (.o(n186086),
	.a(n251567));
   in01s01 U270662 (.o(n186087),
	.a(n251568));
   oa22s01 U270663 (.o(n251569),
	.a(n251583),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1101]),
	.d(FE_OFN324_n251565));
   in01s01 U270664 (.o(n186088),
	.a(n251569));
   oa22s01 U270665 (.o(n251570),
	.a(n251583),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1100]),
	.d(FE_OFN325_n251565));
   in01s01 U270666 (.o(n186089),
	.a(n251570));
   oa22s01 U270667 (.o(n251571),
	.a(n251583),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1099]),
	.d(FE_OFN325_n251565));
   oa22s01 U270668 (.o(n251572),
	.a(n251583),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1098]),
	.d(FE_OFN324_n251565));
   in01s01 U270669 (.o(n186091),
	.a(n251572));
   oa22s01 U270670 (.o(n251573),
	.a(n251583),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1097]),
	.d(FE_OFN324_n251565));
   in01s01 U270671 (.o(n186092),
	.a(n251573));
   in01s01 U270672 (.o(n186093),
	.a(n251574));
   in01s01 U270673 (.o(n186094),
	.a(n251575));
   in01s01 U270674 (.o(n186095),
	.a(n251577));
   oa22s01 U270675 (.o(n251578),
	.a(n251583),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1093]),
	.d(FE_OFN325_n251565));
   in01s01 U270676 (.o(n186096),
	.a(n251578));
   oa22s01 U270677 (.o(n251579),
	.a(n251583),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1092]),
	.d(FE_OFN325_n251565));
   in01s01 U270678 (.o(n186097),
	.a(n251579));
   oa22s01 U270679 (.o(n251580),
	.a(n251583),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1091]),
	.d(FE_OFN325_n251565));
   in01s01 U270680 (.o(n186098),
	.a(n251580));
   oa22s01 U270681 (.o(n251581),
	.a(n251583),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1090]),
	.d(FE_OFN325_n251565));
   in01s01 U270682 (.o(n186099),
	.a(n251581));
   oa22s01 U270683 (.o(n251582),
	.a(n251583),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1089]),
	.d(FE_OFN325_n251565));
   in01s01 U270684 (.o(n186100),
	.a(n251582));
   oa22s01 U270685 (.o(n251584),
	.a(n251583),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1088]),
	.d(FE_OFN324_n251565));
   in01s01 U270686 (.o(n186101),
	.a(n251584));
   in01s01 U270687 (.o(n186102),
	.a(n251585));
   in01s01 U270688 (.o(n186103),
	.a(n251586));
   in01s01 U270689 (.o(n186104),
	.a(n251587));
   oa22s01 U270690 (.o(n251588),
	.a(n251619),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1084]),
	.d(FE_OFN327_n251600));
   in01s01 U270691 (.o(n186106),
	.a(n251589));
   in01s01 U270692 (.o(n186107),
	.a(n251590));
   in01s01 U270693 (.o(n186108),
	.a(n251591));
   in01s01 U270694 (.o(n186109),
	.a(n251592));
   in01s01 U270695 (.o(n186110),
	.a(n251593));
   in01s01 U270696 (.o(n186111),
	.a(n251594));
   in01s01 U270697 (.o(n186112),
	.a(n251595));
   in01s01 U270698 (.o(n186113),
	.a(n251596));
   in01s01 U270699 (.o(n186114),
	.a(n251597));
   in01s01 U270700 (.o(n186115),
	.a(n251598));
   in01s01 U270701 (.o(n186116),
	.a(n251599));
   in01s01 U270702 (.o(n186117),
	.a(n251601));
   in01s01 U270703 (.o(n186118),
	.a(n251602));
   in01s01 U270704 (.o(n186119),
	.a(n251603));
   oa22s01 U270705 (.o(n251604),
	.a(n251619),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1069]),
	.d(FE_OFN327_n251600));
   in01s01 U270706 (.o(n186121),
	.a(n251605));
   in01s01 U270707 (.o(n186122),
	.a(n251606));
   in01s01 U270708 (.o(n186123),
	.a(n251607));
   in01s01 U270709 (.o(n186124),
	.a(n251608));
   in01s01 U270710 (.o(n186125),
	.a(n251609));
   in01s01 U270711 (.o(n186126),
	.a(n251610));
   in01s01 U270712 (.o(n186127),
	.a(n251612));
   oa22s01 U270713 (.o(n251613),
	.a(n251619),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1061]),
	.d(FE_OFN327_n251600));
   in01s01 U270714 (.o(n186128),
	.a(n251613));
   oa22s01 U270715 (.o(n251614),
	.a(n251619),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1060]),
	.d(FE_OFN327_n251600));
   in01s01 U270716 (.o(n186129),
	.a(n251614));
   oa22s01 U270717 (.o(n251615),
	.a(n251619),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1059]),
	.d(FE_OFN327_n251600));
   in01s01 U270718 (.o(n186130),
	.a(n251615));
   oa22s01 U270719 (.o(n251616),
	.a(n251619),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1058]),
	.d(FE_OFN327_n251600));
   in01s01 U270720 (.o(n186131),
	.a(n251616));
   oa22s01 U270721 (.o(n251617),
	.a(n251619),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1057]),
	.d(FE_OFN327_n251600));
   in01s01 U270722 (.o(n186132),
	.a(n251617));
   oa22s01 U270723 (.o(n251620),
	.a(n251619),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1056]),
	.d(FE_OFN327_n251600));
   in01s01 U270724 (.o(n186133),
	.a(n251620));
   in01s01 U270725 (.o(n186134),
	.a(n251622));
   oa22s01 U270726 (.o(n251623),
	.a(n251655),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1054]),
	.d(FE_OFN329_n251637));
   in01s01 U270727 (.o(n186136),
	.a(n251624));
   in01s01 U270728 (.o(n186137),
	.a(n251625));
   in01s01 U270729 (.o(n186138),
	.a(n251626));
   in01s01 U270730 (.o(n186139),
	.a(n251627));
   in01s01 U270731 (.o(n186140),
	.a(n251628));
   in01s01 U270732 (.o(n186141),
	.a(n251629));
   in01s01 U270733 (.o(n186142),
	.a(n251630));
   in01s01 U270734 (.o(n186143),
	.a(n251631));
   in01s01 U270735 (.o(n186144),
	.a(n251632));
   in01s01 U270736 (.o(n186145),
	.a(n251633));
   in01s01 U270737 (.o(n186146),
	.a(n251634));
   in01s01 U270738 (.o(n186147),
	.a(n251635));
   in01s01 U270739 (.o(n186148),
	.a(n251636));
   in01s01 U270740 (.o(n186149),
	.a(n251638));
   oa22s01 U270741 (.o(n251639),
	.a(n251655),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1039]),
	.d(FE_OFN329_n251637));
   in01s01 U270742 (.o(n186151),
	.a(n251640));
   in01s01 U270743 (.o(n186152),
	.a(n251641));
   in01s01 U270744 (.o(n186153),
	.a(n251642));
   in01s01 U270745 (.o(n186154),
	.a(n251643));
   in01s01 U270746 (.o(n186155),
	.a(n251644));
   in01s01 U270747 (.o(n186156),
	.a(n251645));
   in01s01 U270748 (.o(n186157),
	.a(n251646));
   in01s01 U270749 (.o(n186158),
	.a(n251647));
   in01s01 U270750 (.o(n186159),
	.a(n251649));
   oa22s01 U270751 (.o(n251650),
	.a(n251655),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1029]),
	.d(FE_OFN329_n251637));
   in01s01 U270752 (.o(n186160),
	.a(n251650));
   oa22s01 U270753 (.o(n251651),
	.a(n251655),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1028]),
	.d(FE_OFN329_n251637));
   in01s01 U270754 (.o(n186161),
	.a(n251651));
   oa22s01 U270755 (.o(n251652),
	.a(n251655),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1027]),
	.d(FE_OFN329_n251637));
   in01s01 U270756 (.o(n186162),
	.a(n251652));
   oa22s01 U270757 (.o(n251653),
	.a(n251655),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1026]),
	.d(FE_OFN329_n251637));
   in01s01 U270758 (.o(n186163),
	.a(n251653));
   oa22s01 U270759 (.o(n251654),
	.a(n251655),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1025]),
	.d(FE_OFN329_n251637));
   in01s01 U270760 (.o(n186164),
	.a(n251654));
   oa22s01 U270761 (.o(n251656),
	.a(n251655),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1024]),
	.d(FE_OFN329_n251637));
   in01s01 U270762 (.o(n186166),
	.a(n251657));
   in01s01 U270763 (.o(n186167),
	.a(n251658));
   in01s01 U270764 (.o(n186168),
	.a(n251659));
   in01s01 U270765 (.o(n186169),
	.a(n251660));
   in01s01 U270766 (.o(n186170),
	.a(n251661));
   in01s01 U270767 (.o(n186171),
	.a(n251662));
   in01s01 U270768 (.o(n186172),
	.a(n251663));
   in01s01 U270769 (.o(n186173),
	.a(n251664));
   in01s01 U270770 (.o(n186174),
	.a(n251665));
   in01s01 U270771 (.o(n186175),
	.a(n251666));
   in01s01 U270772 (.o(n186176),
	.a(n251667));
   in01s01 U270773 (.o(n186177),
	.a(n251668));
   in01s01 U270774 (.o(n186178),
	.a(n251669));
   in01s01 U270775 (.o(n186179),
	.a(n251670));
   oa22s01 U270776 (.o(n251671),
	.a(n251690),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[2033]),
	.d(FE_OFN331_n251675));
   in01s01 U270777 (.o(n186181),
	.a(n251672));
   in01s01 U270778 (.o(n186182),
	.a(n251673));
   in01s01 U270779 (.o(n186183),
	.a(n251674));
   in01s01 U270780 (.o(n186184),
	.a(n251676));
   in01s01 U270781 (.o(n186185),
	.a(n251677));
   in01s01 U270782 (.o(n186186),
	.a(n251678));
   in01s01 U270783 (.o(n186187),
	.a(n251679));
   in01s01 U270784 (.o(n186188),
	.a(n251680));
   in01s01 U270785 (.o(n186189),
	.a(n251681));
   in01s01 U270786 (.o(n186190),
	.a(n251682));
   in01s01 U270787 (.o(n186191),
	.a(n251684));
   oa22s01 U270788 (.o(n251685),
	.a(n251690),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[2021]),
	.d(FE_OFN331_n251675));
   in01s01 U270789 (.o(n186192),
	.a(n251685));
   oa22s01 U270790 (.o(n251686),
	.a(n251690),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[2020]),
	.d(FE_OFN331_n251675));
   in01s01 U270791 (.o(n186193),
	.a(n251686));
   oa22s01 U270792 (.o(n251687),
	.a(n251690),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[2019]),
	.d(FE_OFN331_n251675));
   in01s01 U270793 (.o(n186194),
	.a(n251687));
   oa22s01 U270794 (.o(n251688),
	.a(n251690),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[2018]),
	.d(FE_OFN331_n251675));
   oa22s01 U270795 (.o(n251689),
	.a(n251690),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[2017]),
	.d(FE_OFN331_n251675));
   in01s01 U270796 (.o(n186196),
	.a(n251689));
   oa22s01 U270797 (.o(n251691),
	.a(n251690),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[2016]),
	.d(FE_OFN331_n251675));
   in01s01 U270798 (.o(n186197),
	.a(n251691));
   in01s01 U270799 (.o(n186198),
	.a(n251692));
   in01s01 U270800 (.o(n186199),
	.a(n251693));
   in01s01 U270801 (.o(n186200),
	.a(n251694));
   in01s01 U270802 (.o(n186201),
	.a(n251695));
   in01s01 U270803 (.o(n186202),
	.a(n251696));
   in01s01 U270804 (.o(n186203),
	.a(n251697));
   in01s01 U270805 (.o(n186204),
	.a(n251698));
   in01s01 U270806 (.o(n186205),
	.a(n251699));
   in01s01 U270807 (.o(n186206),
	.a(n251700));
   in01s01 U270808 (.o(n186207),
	.a(n251701));
   in01s01 U270809 (.o(n186208),
	.a(n251702));
   in01s01 U270810 (.o(n186209),
	.a(n251703));
   oa22s01 U270811 (.o(n251704),
	.a(n251726),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[2003]),
	.d(FE_OFN430_n251710));
   in01s01 U270812 (.o(n186211),
	.a(n251705));
   in01s01 U270813 (.o(n186212),
	.a(n251706));
   in01s01 U270814 (.o(n186213),
	.a(n251707));
   in01s01 U270815 (.o(n186214),
	.a(n251708));
   in01s01 U270816 (.o(n186215),
	.a(n251709));
   in01s01 U270817 (.o(n186216),
	.a(n251711));
   in01s01 U270818 (.o(n186217),
	.a(n251712));
   in01s01 U270819 (.o(n186218),
	.a(n251713));
   in01s01 U270820 (.o(n186219),
	.a(n251714));
   in01s01 U270821 (.o(n186220),
	.a(n251715));
   in01s01 U270822 (.o(n186221),
	.a(n251716));
   in01s01 U270823 (.o(n186222),
	.a(n251717));
   in01s01 U270824 (.o(n186223),
	.a(n251719));
   oa22s01 U270825 (.o(n251720),
	.a(n251726),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1989]),
	.d(FE_OFN430_n251710));
   in01s01 U270826 (.o(n186224),
	.a(n251720));
   oa22s01 U270827 (.o(n251721),
	.a(n251726),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1988]),
	.d(FE_OFN430_n251710));
   oa22s01 U270828 (.o(n251722),
	.a(n251726),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1987]),
	.d(FE_OFN430_n251710));
   in01s01 U270829 (.o(n186226),
	.a(n251722));
   oa22s01 U270830 (.o(n251723),
	.a(n251726),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1986]),
	.d(n251710));
   in01s01 U270831 (.o(n186227),
	.a(n251723));
   oa22s01 U270832 (.o(n251724),
	.a(n251726),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1985]),
	.d(FE_OFN430_n251710));
   in01s01 U270833 (.o(n186228),
	.a(n251724));
   oa22s01 U270834 (.o(n251727),
	.a(n251726),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1984]),
	.d(FE_OFN430_n251710));
   in01s01 U270835 (.o(n186229),
	.a(n251727));
   in01s01 U270836 (.o(n186230),
	.a(n251728));
   in01s01 U270837 (.o(n186231),
	.a(n251729));
   in01s01 U270838 (.o(n186232),
	.a(n251730));
   in01s01 U270839 (.o(n186233),
	.a(n251731));
   in01s01 U270840 (.o(n186234),
	.a(n251732));
   in01s01 U270841 (.o(n186235),
	.a(n251733));
   in01s01 U270842 (.o(n186236),
	.a(n251734));
   in01s01 U270843 (.o(n186237),
	.a(n251735));
   in01s01 U270844 (.o(n186238),
	.a(n251736));
   in01s01 U270845 (.o(n186239),
	.a(n251737));
   oa22s01 U270846 (.o(n251738),
	.a(n251761),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1973]),
	.d(FE_OFN333_n251746));
   in01s01 U270847 (.o(n186241),
	.a(n251739));
   in01s01 U270848 (.o(n186242),
	.a(n251740));
   in01s01 U270849 (.o(n186243),
	.a(n251741));
   in01s01 U270850 (.o(n186244),
	.a(n251742));
   in01s01 U270851 (.o(n186245),
	.a(n251743));
   in01s01 U270852 (.o(n186246),
	.a(n251744));
   in01s01 U270853 (.o(n186247),
	.a(n251745));
   in01s01 U270854 (.o(n186248),
	.a(n251747));
   in01s01 U270855 (.o(n186249),
	.a(n251748));
   in01s01 U270856 (.o(n186250),
	.a(n251749));
   in01s01 U270857 (.o(n186251),
	.a(n251750));
   in01s01 U270858 (.o(n186252),
	.a(n251751));
   in01s01 U270859 (.o(n186253),
	.a(n251752));
   in01s01 U270860 (.o(n186254),
	.a(n251753));
   oa22s01 U270861 (.o(n251755),
	.a(n251761),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1958]),
	.d(FE_OFN333_n251746));
   oa22s01 U270862 (.o(n251756),
	.a(n251761),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1957]),
	.d(FE_OFN333_n251746));
   in01s01 U270863 (.o(n186256),
	.a(n251756));
   oa22s01 U270864 (.o(n251757),
	.a(n251761),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1956]),
	.d(FE_OFN333_n251746));
   in01s01 U270865 (.o(n186257),
	.a(n251757));
   oa22s01 U270866 (.o(n251758),
	.a(n251761),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1955]),
	.d(FE_OFN333_n251746));
   in01s01 U270867 (.o(n186258),
	.a(n251758));
   oa22s01 U270868 (.o(n251759),
	.a(n251761),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1954]),
	.d(n251746));
   in01s01 U270869 (.o(n186259),
	.a(n251759));
   oa22s01 U270870 (.o(n251760),
	.a(n251761),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1953]),
	.d(n251746));
   in01s01 U270871 (.o(n186260),
	.a(n251760));
   oa22s01 U270872 (.o(n251762),
	.a(n251761),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1952]),
	.d(FE_OFN333_n251746));
   in01s01 U270873 (.o(n186261),
	.a(n251762));
   in01s01 U270874 (.o(n186262),
	.a(n251763));
   in01s01 U270875 (.o(n186263),
	.a(n251764));
   in01s01 U270876 (.o(n186264),
	.a(n251765));
   in01s01 U270877 (.o(n186265),
	.a(n251766));
   in01s01 U270878 (.o(n186266),
	.a(n251767));
   in01s01 U270879 (.o(n186267),
	.a(n251768));
   in01s01 U270880 (.o(n186268),
	.a(n251769));
   in01s01 U270881 (.o(n186269),
	.a(n251770));
   oa22s01 U270882 (.o(n251771),
	.a(n251796),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1943]),
	.d(FE_OFN432_n251781));
   in01s01 U270883 (.o(n186271),
	.a(n251772));
   in01s01 U270884 (.o(n186272),
	.a(n251773));
   in01s01 U270885 (.o(n186273),
	.a(n251774));
   in01s01 U270886 (.o(n186274),
	.a(n251775));
   in01s01 U270887 (.o(n186275),
	.a(n251776));
   in01s01 U270888 (.o(n186276),
	.a(n251777));
   in01s01 U270889 (.o(n186277),
	.a(n251778));
   in01s01 U270890 (.o(n186278),
	.a(n251779));
   in01s01 U270891 (.o(n186279),
	.a(n251780));
   in01s01 U270892 (.o(n186280),
	.a(n251782));
   in01s01 U270893 (.o(n186281),
	.a(n251783));
   in01s01 U270894 (.o(n186282),
	.a(n251784));
   in01s01 U270895 (.o(n186283),
	.a(n251785));
   in01s01 U270896 (.o(n186284),
	.a(n251786));
   oa22s01 U270897 (.o(n251787),
	.a(n251796),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1928]),
	.d(FE_OFN432_n251781));
   in01s01 U270898 (.o(n186286),
	.a(n251788));
   in01s01 U270899 (.o(n186287),
	.a(n251790));
   oa22s01 U270900 (.o(n251791),
	.a(n251796),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1925]),
	.d(FE_OFN432_n251781));
   in01s01 U270901 (.o(n186288),
	.a(n251791));
   oa22s01 U270902 (.o(n251792),
	.a(n251796),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1924]),
	.d(FE_OFN432_n251781));
   in01s01 U270903 (.o(n186289),
	.a(n251792));
   oa22s01 U270904 (.o(n251793),
	.a(n251796),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1923]),
	.d(FE_OFN432_n251781));
   in01s01 U270905 (.o(n186290),
	.a(n251793));
   oa22s01 U270906 (.o(n251794),
	.a(n251796),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1922]),
	.d(FE_OFN432_n251781));
   in01s01 U270907 (.o(n186291),
	.a(n251794));
   oa22s01 U270908 (.o(n251795),
	.a(n251796),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1921]),
	.d(FE_OFN432_n251781));
   in01s01 U270909 (.o(n186292),
	.a(n251795));
   oa22s01 U270910 (.o(n251797),
	.a(n251796),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1920]),
	.d(FE_OFN432_n251781));
   in01s01 U270911 (.o(n186293),
	.a(n251797));
   in01s01 U270912 (.o(n186294),
	.a(n251798));
   in01s01 U270913 (.o(n186295),
	.a(n251799));
   in01s01 U270914 (.o(n186296),
	.a(n251800));
   in01s01 U270915 (.o(n186297),
	.a(n251801));
   in01s01 U270916 (.o(n186298),
	.a(n251802));
   in01s01 U270917 (.o(n186299),
	.a(n251803));
   oa22s01 U270918 (.o(n251804),
	.a(n251832),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1913]),
	.d(FE_OFN206_n251816));
   in01s01 U270919 (.o(n186301),
	.a(n251805));
   in01s01 U270920 (.o(n186302),
	.a(n251806));
   in01s01 U270921 (.o(n186303),
	.a(n251807));
   in01s01 U270922 (.o(n186304),
	.a(n251808));
   in01s01 U270923 (.o(n186305),
	.a(n251809));
   in01s01 U270924 (.o(n186306),
	.a(n251810));
   in01s01 U270925 (.o(n186307),
	.a(n251811));
   in01s01 U270926 (.o(n186308),
	.a(n251812));
   in01s01 U270927 (.o(n186309),
	.a(n251813));
   in01s01 U270928 (.o(n186310),
	.a(n251814));
   in01s01 U270929 (.o(n186311),
	.a(n251815));
   in01s01 U270930 (.o(n186312),
	.a(n251817));
   in01s01 U270931 (.o(n186313),
	.a(n251818));
   in01s01 U270932 (.o(n186314),
	.a(n251819));
   oa22s01 U270933 (.o(n251820),
	.a(n251832),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1898]),
	.d(FE_OFN206_n251816));
   in01s01 U270934 (.o(n186316),
	.a(n251821));
   in01s01 U270935 (.o(n186317),
	.a(n251822));
   in01s01 U270936 (.o(n186318),
	.a(n251823));
   in01s01 U270937 (.o(n186319),
	.a(n251825));
   oa22s01 U270938 (.o(n251826),
	.a(n251832),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1893]),
	.d(FE_OFN206_n251816));
   in01s01 U270939 (.o(n186320),
	.a(n251826));
   oa22s01 U270940 (.o(n251827),
	.a(n251832),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1892]),
	.d(FE_OFN206_n251816));
   in01s01 U270941 (.o(n186321),
	.a(n251827));
   oa22s01 U270942 (.o(n251828),
	.a(n251832),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1891]),
	.d(FE_OFN206_n251816));
   in01s01 U270943 (.o(n186322),
	.a(n251828));
   oa22s01 U270944 (.o(n251829),
	.a(n251832),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1890]),
	.d(FE_OFN206_n251816));
   in01s01 U270945 (.o(n186323),
	.a(n251829));
   oa22s01 U270946 (.o(n251830),
	.a(n251832),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1889]),
	.d(FE_OFN206_n251816));
   in01s01 U270947 (.o(n186324),
	.a(n251830));
   oa22s01 U270948 (.o(n251833),
	.a(n251832),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1888]),
	.d(FE_OFN206_n251816));
   in01s01 U270949 (.o(n186325),
	.a(n251833));
   in01s01 U270950 (.o(n186326),
	.a(n251834));
   in01s01 U270951 (.o(n186327),
	.a(n251835));
   in01s01 U270952 (.o(n186328),
	.a(n251836));
   in01s01 U270953 (.o(n186329),
	.a(n251837));
   oa22s01 U270954 (.o(n251838),
	.a(n251867),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1883]),
	.d(FE_OFN560_n251852));
   in01s01 U270955 (.o(n186331),
	.a(n251839));
   in01s01 U270956 (.o(n186332),
	.a(n251840));
   in01s01 U270957 (.o(n186333),
	.a(n251841));
   in01s01 U270958 (.o(n186334),
	.a(n251842));
   in01s01 U270959 (.o(n186335),
	.a(n251843));
   in01s01 U270960 (.o(n186336),
	.a(n251844));
   in01s01 U270961 (.o(n186337),
	.a(n251845));
   in01s01 U270962 (.o(n186338),
	.a(n251846));
   in01s01 U270963 (.o(n186339),
	.a(n251847));
   in01s01 U270964 (.o(n186340),
	.a(n251848));
   in01s01 U270965 (.o(n186341),
	.a(n251849));
   in01s01 U270966 (.o(n186342),
	.a(n251850));
   in01s01 U270967 (.o(n186343),
	.a(n251851));
   in01s01 U270968 (.o(n186344),
	.a(n251853));
   oa22s01 U270969 (.o(n251854),
	.a(n251867),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1868]),
	.d(FE_OFN335_n251852));
   in01s01 U270970 (.o(n186346),
	.a(n251855));
   in01s01 U270971 (.o(n186347),
	.a(n251856));
   in01s01 U270972 (.o(n186348),
	.a(n251857));
   in01s01 U270973 (.o(n186349),
	.a(n251858));
   in01s01 U270974 (.o(n186350),
	.a(n251859));
   in01s01 U270975 (.o(n186351),
	.a(n251861));
   oa22s01 U270976 (.o(n251862),
	.a(n251867),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1861]),
	.d(FE_OFN335_n251852));
   in01s01 U270977 (.o(n186352),
	.a(n251862));
   oa22s01 U270978 (.o(n251863),
	.a(n251867),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1860]),
	.d(FE_OFN335_n251852));
   in01s01 U270979 (.o(n186353),
	.a(n251863));
   oa22s01 U270980 (.o(n251864),
	.a(n251867),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1859]),
	.d(FE_OFN335_n251852));
   in01s01 U270981 (.o(n186354),
	.a(n251864));
   oa22s01 U270982 (.o(n251865),
	.a(n251867),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1858]),
	.d(FE_OFN335_n251852));
   in01s01 U270983 (.o(n186355),
	.a(n251865));
   oa22s01 U270984 (.o(n251866),
	.a(n251867),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1857]),
	.d(FE_OFN335_n251852));
   in01s01 U270985 (.o(n186356),
	.a(n251866));
   oa22s01 U270986 (.o(n251868),
	.a(n251867),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1856]),
	.d(FE_OFN561_n251852));
   in01s01 U270987 (.o(n186357),
	.a(n251868));
   in01s01 U270988 (.o(n186358),
	.a(n251869));
   in01s01 U270989 (.o(n186359),
	.a(n251870));
   oa22s01 U270990 (.o(n251871),
	.a(n251902),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1853]),
	.d(FE_OFN337_n251887));
   in01s01 U270991 (.o(n186361),
	.a(n251872));
   in01s01 U270992 (.o(n186362),
	.a(n251873));
   in01s01 U270993 (.o(n186363),
	.a(n251874));
   in01s01 U270994 (.o(n186364),
	.a(n251875));
   in01s01 U270995 (.o(n186365),
	.a(n251876));
   in01s01 U270996 (.o(n186366),
	.a(n251877));
   in01s01 U270997 (.o(n186367),
	.a(n251878));
   in01s01 U270998 (.o(n186368),
	.a(n251879));
   in01s01 U270999 (.o(n186369),
	.a(n251880));
   in01s01 U271000 (.o(n186370),
	.a(n251881));
   in01s01 U271001 (.o(n186371),
	.a(n251882));
   in01s01 U271002 (.o(n186372),
	.a(n251883));
   in01s01 U271003 (.o(n186373),
	.a(n251884));
   in01s01 U271004 (.o(n186374),
	.a(n251885));
   oa22s01 U271005 (.o(n251886),
	.a(n251902),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1838]),
	.d(FE_OFN337_n251887));
   in01s01 U271006 (.o(n186376),
	.a(n251888));
   in01s01 U271007 (.o(n186377),
	.a(n251889));
   in01s01 U271008 (.o(n186378),
	.a(n251890));
   in01s01 U271009 (.o(n186379),
	.a(n251891));
   in01s01 U271010 (.o(n186380),
	.a(n251892));
   in01s01 U271011 (.o(n186381),
	.a(n251893));
   in01s01 U271012 (.o(n186382),
	.a(n251894));
   in01s01 U271013 (.o(n186383),
	.a(n251896));
   oa22s01 U271014 (.o(n251897),
	.a(n251902),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1829]),
	.d(FE_OFN337_n251887));
   in01s01 U271015 (.o(n186384),
	.a(n251897));
   oa22s01 U271016 (.o(n251898),
	.a(n251902),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1828]),
	.d(FE_OFN337_n251887));
   in01s01 U271017 (.o(n186385),
	.a(n251898));
   oa22s01 U271018 (.o(n251899),
	.a(n251902),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1827]),
	.d(FE_OFN337_n251887));
   in01s01 U271019 (.o(n186386),
	.a(n251899));
   oa22s01 U271020 (.o(n251900),
	.a(n251902),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1826]),
	.d(FE_OFN337_n251887));
   in01s01 U271021 (.o(n186387),
	.a(n251900));
   oa22s01 U271022 (.o(n251901),
	.a(n251902),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1825]),
	.d(FE_OFN337_n251887));
   in01s01 U271023 (.o(n186388),
	.a(n251901));
   oa22s01 U271024 (.o(n251903),
	.a(n251902),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1824]),
	.d(FE_OFN337_n251887));
   in01s01 U271025 (.o(n186389),
	.a(n251903));
   oa22s01 U271026 (.o(n251905),
	.a(n251939),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1823]),
	.d(FE_OFN339_n251923));
   in01s01 U271027 (.o(n186391),
	.a(n251906));
   in01s01 U271028 (.o(n186392),
	.a(n251907));
   in01s01 U271029 (.o(n186393),
	.a(n251908));
   in01s01 U271030 (.o(n186394),
	.a(n251909));
   in01s01 U271031 (.o(n186395),
	.a(n251910));
   in01s01 U271032 (.o(n186396),
	.a(n251911));
   in01s01 U271033 (.o(n186397),
	.a(n251912));
   in01s01 U271034 (.o(n186398),
	.a(n251913));
   in01s01 U271035 (.o(n186399),
	.a(n251914));
   in01s01 U271036 (.o(n186400),
	.a(n251915));
   in01s01 U271037 (.o(n186401),
	.a(n251916));
   in01s01 U271038 (.o(n186402),
	.a(n251917));
   in01s01 U271039 (.o(n186403),
	.a(n251918));
   in01s01 U271040 (.o(n186404),
	.a(n251919));
   oa22s01 U271041 (.o(n251920),
	.a(n251939),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1808]),
	.d(FE_OFN339_n251923));
   in01s01 U271042 (.o(n186406),
	.a(n251921));
   in01s01 U271043 (.o(n186407),
	.a(n251922));
   in01s01 U271044 (.o(n186408),
	.a(n251924));
   in01s01 U271045 (.o(n186409),
	.a(n251925));
   in01s01 U271046 (.o(n186410),
	.a(n251926));
   in01s01 U271047 (.o(n186411),
	.a(n251927));
   in01s01 U271048 (.o(n186412),
	.a(n251928));
   in01s01 U271049 (.o(n186413),
	.a(n251929));
   in01s01 U271050 (.o(n186414),
	.a(n251930));
   in01s01 U271051 (.o(n186415),
	.a(n251932));
   oa22s01 U271052 (.o(n251933),
	.a(n251939),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1797]),
	.d(FE_OFN339_n251923));
   in01s01 U271053 (.o(n186416),
	.a(n251933));
   oa22s01 U271054 (.o(n251934),
	.a(n251939),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1796]),
	.d(FE_OFN339_n251923));
   in01s01 U271055 (.o(n186417),
	.a(n251934));
   oa22s01 U271056 (.o(n251935),
	.a(n251939),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1795]),
	.d(FE_OFN339_n251923));
   in01s01 U271057 (.o(n186418),
	.a(n251935));
   oa22s01 U271058 (.o(n251936),
	.a(n251939),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1794]),
	.d(FE_OFN339_n251923));
   in01s01 U271059 (.o(n186419),
	.a(n251936));
   oa22s01 U271060 (.o(n251937),
	.a(n251939),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1793]),
	.d(FE_OFN339_n251923));
   oa22s01 U271061 (.o(n251940),
	.a(n251939),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1792]),
	.d(FE_OFN339_n251923));
   in01s01 U271062 (.o(n186421),
	.a(n251940));
   in01s01 U271063 (.o(n186422),
	.a(n251942));
   in01s01 U271064 (.o(n186423),
	.a(n251943));
   in01s01 U271065 (.o(n186424),
	.a(n251944));
   in01s01 U271066 (.o(n186425),
	.a(n251945));
   in01s01 U271067 (.o(n186426),
	.a(n251946));
   in01s01 U271068 (.o(n186427),
	.a(n251947));
   in01s01 U271069 (.o(n186428),
	.a(n251948));
   in01s01 U271070 (.o(n186429),
	.a(n251949));
   in01s01 U271071 (.o(n186430),
	.a(n251950));
   in01s01 U271072 (.o(n186431),
	.a(n251951));
   in01s01 U271073 (.o(n186432),
	.a(n251952));
   in01s01 U271074 (.o(n186433),
	.a(n251953));
   in01s01 U271075 (.o(n186434),
	.a(n251954));
   oa22s01 U271076 (.o(n251955),
	.a(n251975),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1778]),
	.d(FE_OFN341_n251960));
   in01s01 U271077 (.o(n186436),
	.a(n251956));
   in01s01 U271078 (.o(n186437),
	.a(n251957));
   in01s01 U271079 (.o(n186438),
	.a(n251958));
   in01s01 U271080 (.o(n186439),
	.a(n251959));
   in01s01 U271081 (.o(n186440),
	.a(n251961));
   in01s01 U271082 (.o(n186441),
	.a(n251962));
   in01s01 U271083 (.o(n186442),
	.a(n251963));
   in01s01 U271084 (.o(n186443),
	.a(n251964));
   in01s01 U271085 (.o(n186444),
	.a(n251965));
   in01s01 U271086 (.o(n186445),
	.a(n251966));
   in01s01 U271087 (.o(n186446),
	.a(n251967));
   in01s01 U271088 (.o(n186447),
	.a(n251969));
   oa22s01 U271089 (.o(n251970),
	.a(n251975),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1765]),
	.d(FE_OFN341_n251960));
   in01s01 U271090 (.o(n186448),
	.a(n251970));
   oa22s01 U271091 (.o(n251971),
	.a(n251975),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1764]),
	.d(FE_OFN341_n251960));
   in01s01 U271092 (.o(n186449),
	.a(n251971));
   oa22s01 U271093 (.o(n251972),
	.a(n251975),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1763]),
	.d(FE_OFN341_n251960));
   oa22s01 U271094 (.o(n251973),
	.a(n251975),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1762]),
	.d(FE_OFN341_n251960));
   in01s01 U271095 (.o(n186451),
	.a(n251973));
   oa22s01 U271096 (.o(n251974),
	.a(n251975),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1761]),
	.d(FE_OFN341_n251960));
   in01s01 U271097 (.o(n186452),
	.a(n251974));
   oa22s01 U271098 (.o(n251976),
	.a(n251975),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1760]),
	.d(FE_OFN341_n251960));
   in01s01 U271099 (.o(n186453),
	.a(n251976));
   in01s01 U271100 (.o(n186454),
	.a(n251978));
   in01s01 U271101 (.o(n186455),
	.a(n251979));
   in01s01 U271102 (.o(n186456),
	.a(n251980));
   in01s01 U271103 (.o(n186457),
	.a(n251981));
   in01s01 U271104 (.o(n186458),
	.a(n251982));
   in01s01 U271105 (.o(n186459),
	.a(n251983));
   in01s01 U271106 (.o(n186460),
	.a(n251984));
   in01s01 U271107 (.o(n186461),
	.a(n251985));
   in01s01 U271108 (.o(n186462),
	.a(n251986));
   in01s01 U271109 (.o(n186463),
	.a(n251987));
   in01s01 U271110 (.o(n186464),
	.a(n251988));
   oa22s01 U271111 (.o(n251989),
	.a(n252011),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1748]),
	.d(FE_OFN434_n251996));
   in01s01 U271112 (.o(n186466),
	.a(n251990));
   in01s01 U271113 (.o(n186467),
	.a(n251991));
   in01s01 U271114 (.o(n186468),
	.a(n251992));
   in01s01 U271115 (.o(n186469),
	.a(n251993));
   in01s01 U271116 (.o(n186470),
	.a(n251994));
   in01s01 U271117 (.o(n186471),
	.a(n251995));
   in01s01 U271118 (.o(n186472),
	.a(n251997));
   in01s01 U271119 (.o(n186473),
	.a(n251998));
   in01s01 U271120 (.o(n186474),
	.a(n251999));
   in01s01 U271121 (.o(n186475),
	.a(n252000));
   in01s01 U271122 (.o(n186476),
	.a(n252001));
   in01s01 U271123 (.o(n186477),
	.a(n252002));
   in01s01 U271124 (.o(n186478),
	.a(n252003));
   in01s01 U271125 (.o(n186479),
	.a(n252005));
   oa22s01 U271126 (.o(n252006),
	.a(n252011),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1733]),
	.d(FE_OFN434_n251996));
   oa22s01 U271127 (.o(n252007),
	.a(n252011),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1732]),
	.d(FE_OFN434_n251996));
   in01s01 U271128 (.o(n186481),
	.a(n252007));
   oa22s01 U271129 (.o(n252008),
	.a(n252011),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1731]),
	.d(FE_OFN434_n251996));
   in01s01 U271130 (.o(n186482),
	.a(n252008));
   oa22s01 U271131 (.o(n252009),
	.a(n252011),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1730]),
	.d(FE_OFN434_n251996));
   in01s01 U271132 (.o(n186483),
	.a(n252009));
   oa22s01 U271133 (.o(n252010),
	.a(n252011),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1729]),
	.d(FE_OFN434_n251996));
   in01s01 U271134 (.o(n186484),
	.a(n252010));
   oa22s01 U271135 (.o(n252012),
	.a(n252011),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1728]),
	.d(FE_OFN434_n251996));
   in01s01 U271136 (.o(n186485),
	.a(n252012));
   in01s01 U271137 (.o(n186486),
	.a(n252014));
   in01s01 U271138 (.o(n186487),
	.a(n252015));
   in01s01 U271139 (.o(n186488),
	.a(n252016));
   in01s01 U271140 (.o(n186489),
	.a(n252017));
   in01s01 U271141 (.o(n186490),
	.a(n252018));
   in01s01 U271142 (.o(n186491),
	.a(n252019));
   oa22s01 U271143 (.o(n252020),
	.a(n252048),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1721]),
	.d(FE_OFN343_n252032));
   in01s01 U271144 (.o(n186492),
	.a(n252020));
   in01s01 U271145 (.o(n186493),
	.a(n252021));
   oa22s01 U271146 (.o(n252022),
	.a(n252048),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1719]),
	.d(FE_OFN343_n252032));
   in01s01 U271147 (.o(n186494),
	.a(n252022));
   oa22s01 U271148 (.o(n252023),
	.a(n252048),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1718]),
	.d(FE_OFN343_n252032));
   oa22s01 U271149 (.o(n252024),
	.a(n252048),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1717]),
	.d(FE_OFN343_n252032));
   in01s01 U271150 (.o(n186496),
	.a(n252024));
   in01s01 U271151 (.o(n186497),
	.a(n252025));
   oa22s01 U271152 (.o(n252026),
	.a(n252048),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1715]),
	.d(FE_OFN343_n252032));
   in01s01 U271153 (.o(n186498),
	.a(n252026));
   in01s01 U271154 (.o(n186499),
	.a(n252027));
   oa22s01 U271155 (.o(n252028),
	.a(n252048),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1713]),
	.d(FE_OFN343_n252032));
   in01s01 U271156 (.o(n186500),
	.a(n252028));
   oa22s01 U271157 (.o(n252029),
	.a(n252048),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1712]),
	.d(FE_OFN343_n252032));
   in01s01 U271158 (.o(n186501),
	.a(n252029));
   in01s01 U271159 (.o(n186502),
	.a(n252030));
   in01s01 U271160 (.o(n186503),
	.a(n252031));
   oa22s01 U271161 (.o(n252033),
	.a(n252048),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1709]),
	.d(FE_OFN343_n252032));
   in01s01 U271162 (.o(n186504),
	.a(n252033));
   in01s01 U271163 (.o(n186505),
	.a(n252034));
   in01s01 U271164 (.o(n186506),
	.a(n252035));
   in01s01 U271165 (.o(n186507),
	.a(n252036));
   in01s01 U271166 (.o(n186508),
	.a(n252037));
   in01s01 U271167 (.o(n186509),
	.a(n252038));
   oa22s01 U271168 (.o(n252039),
	.a(n252048),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1703]),
	.d(FE_OFN343_n252032));
   in01s01 U271169 (.o(n186511),
	.a(n252041));
   oa22s01 U271170 (.o(n252042),
	.a(n252048),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1701]),
	.d(FE_OFN343_n252032));
   in01s01 U271171 (.o(n186512),
	.a(n252042));
   oa22s01 U271172 (.o(n252043),
	.a(n252048),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1700]),
	.d(FE_OFN343_n252032));
   in01s01 U271173 (.o(n186513),
	.a(n252043));
   oa22s01 U271174 (.o(n252044),
	.a(n252048),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1699]),
	.d(FE_OFN343_n252032));
   in01s01 U271175 (.o(n186514),
	.a(n252044));
   oa22s01 U271176 (.o(n252045),
	.a(n252048),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1698]),
	.d(FE_OFN343_n252032));
   in01s01 U271177 (.o(n186515),
	.a(n252045));
   oa22s01 U271178 (.o(n252046),
	.a(n252048),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1697]),
	.d(FE_OFN343_n252032));
   in01s01 U271179 (.o(n186516),
	.a(n252046));
   oa22s01 U271180 (.o(n252049),
	.a(n252048),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1696]),
	.d(FE_OFN343_n252032));
   in01s01 U271181 (.o(n186517),
	.a(n252049));
   oa22s01 U271182 (.o(n252051),
	.a(n252084),
	.b(regtop_v1_hdi00_d[31]),
	.c(regtop_dchdi_w1_hdi00[1695]),
	.d(FE_OFN436_n252069));
   in01s01 U271183 (.o(n186518),
	.a(n252051));
   oa22s01 U271184 (.o(n252052),
	.a(n252084),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1694]),
	.d(FE_OFN436_n252069));
   in01s01 U271185 (.o(n186519),
	.a(n252052));
   oa22s01 U271186 (.o(n252053),
	.a(n252084),
	.b(regtop_v1_hdi00_d[29]),
	.c(regtop_dchdi_w1_hdi00[1693]),
	.d(FE_OFN437_n252069));
   in01s01 U271187 (.o(n186520),
	.a(n252053));
   oa22s01 U271188 (.o(n252054),
	.a(n252084),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1692]),
	.d(FE_OFN437_n252069));
   in01s01 U271189 (.o(n186521),
	.a(n252054));
   oa22s01 U271190 (.o(n252055),
	.a(n252084),
	.b(regtop_v1_hdi00_d[27]),
	.c(regtop_dchdi_w1_hdi00[1691]),
	.d(FE_OFN437_n252069));
   in01s01 U271191 (.o(n186522),
	.a(n252055));
   oa22s01 U271192 (.o(n252056),
	.a(n252084),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1690]),
	.d(FE_OFN437_n252069));
   in01s01 U271193 (.o(n186523),
	.a(n252056));
   oa22s01 U271194 (.o(n252057),
	.a(n252084),
	.b(regtop_v1_hdi00_d[25]),
	.c(regtop_dchdi_w1_hdi00[1689]),
	.d(FE_OFN437_n252069));
   in01s01 U271195 (.o(n186524),
	.a(n252057));
   oa22s01 U271196 (.o(n252058),
	.a(n252084),
	.b(regtop_v1_hdi00_d[24]),
	.c(regtop_dchdi_w1_hdi00[1688]),
	.d(FE_OFN436_n252069));
   oa22s01 U271197 (.o(n252059),
	.a(n252084),
	.b(regtop_v1_hdi00_d[23]),
	.c(regtop_dchdi_w1_hdi00[1687]),
	.d(FE_OFN436_n252069));
   in01s01 U271198 (.o(n186526),
	.a(n252059));
   oa22s01 U271199 (.o(n252060),
	.a(n252084),
	.b(regtop_v1_hdi00_d[22]),
	.c(regtop_dchdi_w1_hdi00[1686]),
	.d(FE_OFN437_n252069));
   in01s01 U271200 (.o(n186527),
	.a(n252060));
   oa22s01 U271201 (.o(n252061),
	.a(n252084),
	.b(regtop_v1_hdi00_d[21]),
	.c(regtop_dchdi_w1_hdi00[1685]),
	.d(FE_OFN437_n252069));
   in01s01 U271202 (.o(n186528),
	.a(n252061));
   oa22s01 U271203 (.o(n252062),
	.a(n252084),
	.b(regtop_v1_hdi00_d[20]),
	.c(regtop_dchdi_w1_hdi00[1684]),
	.d(FE_OFN437_n252069));
   in01s01 U271204 (.o(n186529),
	.a(n252062));
   oa22s01 U271205 (.o(n252063),
	.a(n252084),
	.b(regtop_v1_hdi00_d[19]),
	.c(regtop_dchdi_w1_hdi00[1683]),
	.d(FE_OFN437_n252069));
   in01s01 U271206 (.o(n186530),
	.a(n252063));
   oa22s01 U271207 (.o(n252064),
	.a(n252084),
	.b(regtop_v1_hdi00_d[18]),
	.c(regtop_dchdi_w1_hdi00[1682]),
	.d(FE_OFN437_n252069));
   in01s01 U271208 (.o(n186531),
	.a(n252064));
   oa22s01 U271209 (.o(n252065),
	.a(n252084),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1681]),
	.d(FE_OFN436_n252069));
   in01s01 U271210 (.o(n186532),
	.a(n252065));
   oa22s01 U271211 (.o(n252066),
	.a(n252084),
	.b(regtop_v1_hdi00_d[16]),
	.c(regtop_dchdi_w1_hdi00[1680]),
	.d(FE_OFN437_n252069));
   in01s01 U271212 (.o(n186533),
	.a(n252066));
   oa22s01 U271213 (.o(n252067),
	.a(n252084),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1679]),
	.d(FE_OFN436_n252069));
   in01s01 U271214 (.o(n186534),
	.a(n252067));
   oa22s01 U271215 (.o(n252068),
	.a(n252084),
	.b(regtop_v1_hdi00_d[14]),
	.c(regtop_dchdi_w1_hdi00[1678]),
	.d(FE_OFN436_n252069));
   in01s01 U271216 (.o(n186535),
	.a(n252068));
   oa22s01 U271217 (.o(n252070),
	.a(n252084),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1677]),
	.d(FE_OFN436_n252069));
   in01s01 U271218 (.o(n186536),
	.a(n252070));
   oa22s01 U271219 (.o(n252071),
	.a(n252084),
	.b(regtop_v1_hdi00_d[12]),
	.c(regtop_dchdi_w1_hdi00[1676]),
	.d(FE_OFN436_n252069));
   in01s01 U271220 (.o(n186537),
	.a(n252071));
   oa22s01 U271221 (.o(n252072),
	.a(n252084),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1675]),
	.d(FE_OFN437_n252069));
   in01s01 U271222 (.o(n186538),
	.a(n252072));
   oa22s01 U271223 (.o(n252073),
	.a(n252084),
	.b(regtop_v1_hdi00_d[10]),
	.c(regtop_dchdi_w1_hdi00[1674]),
	.d(FE_OFN437_n252069));
   in01s01 U271224 (.o(n186539),
	.a(n252073));
   oa22s01 U271225 (.o(n252074),
	.a(n252084),
	.b(regtop_v1_hdi00_d[9]),
	.c(regtop_dchdi_w1_hdi00[1673]),
	.d(FE_OFN436_n252069));
   oa22s01 U271226 (.o(n252075),
	.a(n252084),
	.b(regtop_v1_hdi00_d[8]),
	.c(regtop_dchdi_w1_hdi00[1672]),
	.d(FE_OFN436_n252069));
   in01s01 U271227 (.o(n186541),
	.a(n252075));
   oa22s01 U271228 (.o(n252076),
	.a(n252084),
	.b(regtop_v1_hdi00_d[7]),
	.c(regtop_dchdi_w1_hdi00[1671]),
	.d(FE_OFN437_n252069));
   in01s01 U271229 (.o(n186542),
	.a(n252076));
   oa22s01 U271230 (.o(n252078),
	.a(n252084),
	.b(regtop_v1_hdi00_d[6]),
	.c(regtop_dchdi_w1_hdi00[1670]),
	.d(FE_OFN437_n252069));
   in01s01 U271231 (.o(n186543),
	.a(n252078));
   oa22s01 U271232 (.o(n252079),
	.a(n252084),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1669]),
	.d(FE_OFN437_n252069));
   in01s01 U271233 (.o(n186544),
	.a(n252079));
   oa22s01 U271234 (.o(n252080),
	.a(n252084),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1668]),
	.d(FE_OFN437_n252069));
   in01s01 U271235 (.o(n186545),
	.a(n252080));
   oa22s01 U271236 (.o(n252081),
	.a(n252084),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1667]),
	.d(FE_OFN437_n252069));
   in01s01 U271237 (.o(n186546),
	.a(n252081));
   oa22s01 U271238 (.o(n252082),
	.a(n252084),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1666]),
	.d(FE_OFN437_n252069));
   in01s01 U271239 (.o(n186547),
	.a(n252082));
   oa22s01 U271240 (.o(n252083),
	.a(n252084),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1665]),
	.d(FE_OFN437_n252069));
   in01s01 U271241 (.o(n186548),
	.a(n252083));
   oa22s01 U271242 (.o(n252085),
	.a(n252084),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1664]),
	.d(FE_OFN436_n252069));
   in01s01 U271243 (.o(n186549),
	.a(n252085));
   in01s01 U271244 (.o(n186550),
	.a(n252087));
   in01s01 U271245 (.o(n186551),
	.a(n252088));
   in01s01 U271246 (.o(n186552),
	.a(n252089));
   in01s01 U271247 (.o(n186553),
	.a(n252090));
   in01s01 U271248 (.o(n186554),
	.a(n252091));
   oa22s01 U271249 (.o(n252092),
	.a(n252120),
	.b(regtop_v1_hdi00_d[26]),
	.c(regtop_dchdi_w1_hdi00[1658]),
	.d(FE_OFN208_n252105));
   in01s01 U271250 (.o(n186556),
	.a(n252093));
   in01s01 U271251 (.o(n186557),
	.a(n252094));
   in01s01 U271252 (.o(n186558),
	.a(n252095));
   in01s01 U271253 (.o(n186559),
	.a(n252096));
   in01s01 U271254 (.o(n186560),
	.a(n252097));
   in01s01 U271255 (.o(n186561),
	.a(n252098));
   in01s01 U271256 (.o(n186562),
	.a(n252099));
   in01s01 U271257 (.o(n186563),
	.a(n252100));
   in01s01 U271258 (.o(n186564),
	.a(n252101));
   in01s01 U271259 (.o(n186565),
	.a(n252102));
   in01s01 U271260 (.o(n186566),
	.a(n252103));
   in01s01 U271261 (.o(n186567),
	.a(n252104));
   in01s01 U271262 (.o(n186568),
	.a(n252106));
   in01s01 U271263 (.o(n186569),
	.a(n252107));
   oa22s01 U271264 (.o(n252108),
	.a(n252120),
	.b(regtop_v1_hdi00_d[11]),
	.c(regtop_dchdi_w1_hdi00[1643]),
	.d(FE_OFN208_n252105));
   in01s01 U271265 (.o(n186571),
	.a(n252109));
   in01s01 U271266 (.o(n186572),
	.a(n252110));
   in01s01 U271267 (.o(n186573),
	.a(n252111));
   in01s01 U271268 (.o(n186574),
	.a(n252112));
   in01s01 U271269 (.o(n186575),
	.a(n252114));
   oa22s01 U271270 (.o(n252115),
	.a(n252120),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1637]),
	.d(FE_OFN208_n252105));
   in01s01 U271271 (.o(n186576),
	.a(n252115));
   oa22s01 U271272 (.o(n252116),
	.a(n252120),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1636]),
	.d(FE_OFN208_n252105));
   in01s01 U271273 (.o(n186577),
	.a(n252116));
   oa22s01 U271274 (.o(n252117),
	.a(n252120),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1635]),
	.d(FE_OFN208_n252105));
   in01s01 U271275 (.o(n186578),
	.a(n252117));
   oa22s01 U271276 (.o(n252118),
	.a(n252120),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1634]),
	.d(FE_OFN208_n252105));
   in01s01 U271277 (.o(n186579),
	.a(n252118));
   oa22s01 U271278 (.o(n252119),
	.a(n252120),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1633]),
	.d(FE_OFN208_n252105));
   in01s01 U271279 (.o(n186580),
	.a(n252119));
   oa22s01 U271280 (.o(n252121),
	.a(n252120),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1632]),
	.d(FE_OFN208_n252105));
   in01s01 U271281 (.o(n186581),
	.a(n252121));
   in01s01 U271282 (.o(n186582),
	.a(n252123));
   in01s01 U271283 (.o(n186583),
	.a(n252124));
   in01s01 U271284 (.o(n186584),
	.a(n252125));
   oa22s01 U271285 (.o(n252126),
	.a(n252157),
	.b(regtop_v1_hdi00_d[28]),
	.c(regtop_dchdi_w1_hdi00[1628]),
	.d(FE_OFN345_n252141));
   in01s01 U271286 (.o(n186586),
	.a(n252127));
   in01s01 U271287 (.o(n186587),
	.a(n252128));
   in01s01 U271288 (.o(n186588),
	.a(n252129));
   in01s01 U271289 (.o(n186589),
	.a(n252130));
   in01s01 U271290 (.o(n186590),
	.a(n252131));
   in01s01 U271291 (.o(n186591),
	.a(n252132));
   in01s01 U271292 (.o(n186592),
	.a(n252133));
   in01s01 U271293 (.o(n186593),
	.a(n252134));
   in01s01 U271294 (.o(n186594),
	.a(n252135));
   in01s01 U271295 (.o(n186595),
	.a(n252136));
   in01s01 U271296 (.o(n186596),
	.a(n252137));
   in01s01 U271297 (.o(n186597),
	.a(n252138));
   in01s01 U271298 (.o(n186598),
	.a(n252139));
   in01s01 U271299 (.o(n186599),
	.a(n252140));
   oa22s01 U271300 (.o(n252142),
	.a(n252157),
	.b(regtop_v1_hdi00_d[13]),
	.c(regtop_dchdi_w1_hdi00[1613]),
	.d(FE_OFN345_n252141));
   in01s01 U271301 (.o(n186601),
	.a(n252143));
   in01s01 U271302 (.o(n186602),
	.a(n252144));
   in01s01 U271303 (.o(n186603),
	.a(n252145));
   in01s01 U271304 (.o(n186604),
	.a(n252146));
   in01s01 U271305 (.o(n186605),
	.a(n252147));
   in01s01 U271306 (.o(n186606),
	.a(n252148));
   in01s01 U271307 (.o(n186607),
	.a(n252150));
   oa22s01 U271308 (.o(n252151),
	.a(n252157),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1605]),
	.d(FE_OFN346_n252141));
   in01s01 U271309 (.o(n186608),
	.a(n252151));
   oa22s01 U271310 (.o(n252152),
	.a(n252157),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1604]),
	.d(FE_OFN346_n252141));
   in01s01 U271311 (.o(n186609),
	.a(n252152));
   oa22s01 U271312 (.o(n252153),
	.a(n252157),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1603]),
	.d(FE_OFN346_n252141));
   in01s01 U271313 (.o(n186610),
	.a(n252153));
   oa22s01 U271314 (.o(n252154),
	.a(n252157),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1602]),
	.d(FE_OFN346_n252141));
   in01s01 U271315 (.o(n186611),
	.a(n252154));
   oa22s01 U271316 (.o(n252155),
	.a(n252157),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1601]),
	.d(FE_OFN346_n252141));
   in01s01 U271317 (.o(n186612),
	.a(n252155));
   oa22s01 U271318 (.o(n252158),
	.a(n252157),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1600]),
	.d(FE_OFN345_n252141));
   in01s01 U271319 (.o(n186613),
	.a(n252158));
   in01s01 U271320 (.o(n186614),
	.a(n252160));
   oa22s01 U271321 (.o(n252161),
	.a(n252193),
	.b(regtop_v1_hdi00_d[30]),
	.c(regtop_dchdi_w1_hdi00[1598]),
	.d(FE_OFN348_n252178));
   in01s01 U271322 (.o(n186616),
	.a(n252162));
   in01s01 U271323 (.o(n186617),
	.a(n252163));
   in01s01 U271324 (.o(n186618),
	.a(n252164));
   in01s01 U271325 (.o(n186619),
	.a(n252165));
   in01s01 U271326 (.o(n186620),
	.a(n252166));
   in01s01 U271327 (.o(n186621),
	.a(n252167));
   in01s01 U271328 (.o(n186622),
	.a(n252168));
   in01s01 U271329 (.o(n186623),
	.a(n252169));
   in01s01 U271330 (.o(n186624),
	.a(n252170));
   in01s01 U271331 (.o(n186625),
	.a(n252171));
   in01s01 U271332 (.o(n186626),
	.a(n252172));
   in01s01 U271333 (.o(n186627),
	.a(n252173));
   in01s01 U271334 (.o(n186628),
	.a(n252174));
   in01s01 U271335 (.o(n186629),
	.a(n252175));
   oa22s01 U271336 (.o(n252176),
	.a(n252193),
	.b(regtop_v1_hdi00_d[15]),
	.c(regtop_dchdi_w1_hdi00[1583]),
	.d(FE_OFN348_n252178));
   in01s01 U271337 (.o(n186631),
	.a(n252177));
   in01s01 U271338 (.o(n186632),
	.a(n252179));
   in01s01 U271339 (.o(n186633),
	.a(n252180));
   in01s01 U271340 (.o(n186634),
	.a(n252181));
   in01s01 U271341 (.o(n186635),
	.a(n252182));
   in01s01 U271342 (.o(n186636),
	.a(n252183));
   in01s01 U271343 (.o(n186637),
	.a(n252184));
   in01s01 U271344 (.o(n186638),
	.a(n252185));
   in01s01 U271345 (.o(n186639),
	.a(n252187));
   oa22s01 U271346 (.o(n252188),
	.a(n252193),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1573]),
	.d(FE_OFN348_n252178));
   in01s01 U271347 (.o(n186640),
	.a(n252188));
   oa22s01 U271348 (.o(n252189),
	.a(n252193),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1572]),
	.d(FE_OFN348_n252178));
   in01s01 U271349 (.o(n186641),
	.a(n252189));
   oa22s01 U271350 (.o(n252190),
	.a(n252193),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1571]),
	.d(FE_OFN348_n252178));
   in01s01 U271351 (.o(n186642),
	.a(n252190));
   oa22s01 U271352 (.o(n252191),
	.a(n252193),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1570]),
	.d(FE_OFN348_n252178));
   in01s01 U271353 (.o(n186643),
	.a(n252191));
   oa22s01 U271354 (.o(n252192),
	.a(n252193),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1569]),
	.d(FE_OFN348_n252178));
   in01s01 U271355 (.o(n186644),
	.a(n252192));
   oa22s01 U271356 (.o(n252194),
	.a(n252193),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1568]),
	.d(FE_OFN348_n252178));
   in01s01 U271357 (.o(n186646),
	.a(n252197));
   in01s01 U271358 (.o(n186647),
	.a(n252198));
   in01s01 U271359 (.o(n186648),
	.a(n252199));
   in01s01 U271360 (.o(n186649),
	.a(n252200));
   in01s01 U271361 (.o(n186650),
	.a(n252201));
   in01s01 U271362 (.o(n186651),
	.a(n252202));
   in01s01 U271363 (.o(n186652),
	.a(n252203));
   in01s01 U271364 (.o(n186653),
	.a(n252204));
   in01s01 U271365 (.o(n186654),
	.a(n252205));
   in01s01 U271366 (.o(n186655),
	.a(n252206));
   in01s01 U271367 (.o(n186656),
	.a(n252207));
   in01s01 U271368 (.o(n186657),
	.a(n252208));
   in01s01 U271369 (.o(n186658),
	.a(n252209));
   in01s01 U271370 (.o(n186659),
	.a(n252210));
   oa22s01 U271371 (.o(n252211),
	.a(n252230),
	.b(regtop_v1_hdi00_d[17]),
	.c(regtop_dchdi_w1_hdi00[1553]),
	.d(FE_OFN350_n252215));
   in01s01 U271372 (.o(n186661),
	.a(n252212));
   in01s01 U271373 (.o(n186662),
	.a(n252213));
   in01s01 U271374 (.o(n186663),
	.a(n252214));
   in01s01 U271375 (.o(n186664),
	.a(n252216));
   in01s01 U271376 (.o(n186665),
	.a(n252217));
   in01s01 U271377 (.o(n186666),
	.a(n252218));
   in01s01 U271378 (.o(n186667),
	.a(n252219));
   in01s01 U271379 (.o(n186668),
	.a(n252220));
   in01s01 U271380 (.o(n186669),
	.a(n252221));
   in01s01 U271381 (.o(n186670),
	.a(n252222));
   in01s01 U271382 (.o(n186671),
	.a(n252224));
   oa22s01 U271383 (.o(n252225),
	.a(n252230),
	.b(regtop_v1_hdi00_d[5]),
	.c(regtop_dchdi_w1_hdi00[1541]),
	.d(FE_OFN350_n252215));
   in01s01 U271384 (.o(n186672),
	.a(n252225));
   oa22s01 U271385 (.o(n252226),
	.a(n252230),
	.b(regtop_v1_hdi00_d[4]),
	.c(regtop_dchdi_w1_hdi00[1540]),
	.d(FE_OFN350_n252215));
   in01s01 U271386 (.o(n186673),
	.a(n252226));
   oa22s01 U271387 (.o(n252227),
	.a(n252230),
	.b(regtop_v1_hdi00_d[3]),
	.c(regtop_dchdi_w1_hdi00[1539]),
	.d(FE_OFN350_n252215));
   in01s01 U271388 (.o(n186674),
	.a(n252227));
   oa22s01 U271389 (.o(n252228),
	.a(n252230),
	.b(regtop_v1_hdi00_d[2]),
	.c(regtop_dchdi_w1_hdi00[1538]),
	.d(FE_OFN350_n252215));
   oa22s01 U271390 (.o(n252229),
	.a(n252230),
	.b(regtop_v1_hdi00_d[1]),
	.c(regtop_dchdi_w1_hdi00[1537]),
	.d(FE_OFN350_n252215));
   in01s01 U271391 (.o(n186676),
	.a(n252229));
   oa22s01 U271392 (.o(n252231),
	.a(n252230),
	.b(regtop_v1_hdi00_d[0]),
	.c(regtop_dchdi_w1_hdi00[1536]),
	.d(FE_OFN350_n252215));
   in01s01 U271393 (.o(n186677),
	.a(n252231));
   ao12s01 U271394 (.o(n252233),
	.a(regtop_g_memr_ok_r),
	.b(n252232),
	.c(wbb_ack_o));
   in01s01 U271395 (.o(n186678),
	.a(n252233));
   na02f01 U271396 (.o(n252255),
	.a(regtop_g_ferror_r),
	.b(regtop_g_paramadr_r[6]));
   no02f01 U271397 (.o(n252821),
	.a(n252234),
	.b(n252255));
   in01s01 U271398 (.o(n252235),
	.a(n252247));
   no02s01 U271399 (.o(n252236),
	.a(n252676),
	.b(n252235));
   no02s01 U271400 (.o(n252241),
	.a(n252821),
	.b(n252236));
   na02s01 U271401 (.o(n252312),
	.a(regtop_g_ferror_r),
	.b(FE_OFN488_n245940));
   na02s01 U271402 (.o(n252750),
	.a(n252240),
	.b(n252239));
   ao22s01 U271403 (.o(n252244),
	.a(n252269),
	.b(regtop_g_wd_r[18]),
	.c(regtop_g_icfp_r),
	.d(FE_OFN352_n252242));
   in01s01 U271404 (.o(n252894),
	.a(regtop_g_wd_r[18]));
   na03s01 U271405 (.o(n252243),
	.a(n252822),
	.b(regtop_g_isfp_r),
	.c(n252273));
   na02s01 U271406 (.o(n186679),
	.a(n252244),
	.b(n252243));
   in01s01 U271407 (.o(n252246),
	.a(n252245));
   no02s01 U271408 (.o(n252674),
	.a(n252253),
	.b(n252255));
   na02s01 U271409 (.o(n252306),
	.a(n252680),
	.b(n252674));
   na02s01 U271410 (.o(n252250),
	.a(n252246),
	.b(n252306));
   na02s01 U271411 (.o(n252248),
	.a(n252567),
	.b(n252247));
   in01s01 U271412 (.o(n252249),
	.a(n252248));
   no02s01 U271413 (.o(n252363),
	.a(n252254),
	.b(n252255));
   na02s01 U271414 (.o(n252298),
	.a(n252680),
	.b(n252363));
   no02s01 U271415 (.o(n252256),
	.a(n252575),
	.b(n252255));
   na02s01 U271416 (.o(n252296),
	.a(n252567),
	.b(n252256));
   na03s01 U271417 (.o(n252261),
	.a(n252260),
	.b(regtop_g_isfb_r),
	.c(n252273));
   in01f01 U271418 (.o(n252950),
	.a(regtop_g_wd_r[8]));
   oa12s01 U271419 (.o(n252263),
	.a(regtop_g_issr_r),
	.b(n252950),
	.c(n252264));
   oa22s01 U271420 (.o(n186681),
	.a(n252950),
	.b(n252273),
	.c(n252269),
	.d(n252263));
   in01f01 U271421 (.o(n252928),
	.a(regtop_g_wd_r[9]));
   oa12s01 U271422 (.o(n252265),
	.a(regtop_g_issw_r),
	.b(n252928),
	.c(n252264));
   oa22s01 U271423 (.o(n186682),
	.a(n252928),
	.b(n252273),
	.c(n252269),
	.d(n252265));
   in01f02 U271424 (.o(n252940),
	.a(regtop_g_wd_r[1]));
   ao12s01 U271425 (.o(n252267),
	.a(n252266),
	.b(n252270),
	.c(regtop_g_wd_r[1]));
   na02s01 U271426 (.o(n252268),
	.a(n252267),
	.b(n252273));
   oa12s01 U271427 (.o(n186684),
	.a(n252268),
	.b(n252273),
	.c(n252940));
   in01f02 U271428 (.o(n252938),
	.a(regtop_g_wd_r[2]));
   na02s01 U271429 (.o(n252272),
	.a(n252271),
	.b(regtop_g_ispi_r));
   oa12s01 U271430 (.o(n186685),
	.a(n252272),
	.b(n252273),
	.c(n252938));
   in01f03 U271431 (.o(n252953),
	.a(regtop_g_wd_r[0]));
   na02s01 U271432 (.o(n252277),
	.a(n252283),
	.b(regtop_g_udb_cpu_r[0]));
   oa12s01 U271433 (.o(n186693),
	.a(n252277),
	.b(n252953),
	.c(n252285));
   na02s01 U271434 (.o(n252278),
	.a(n252283),
	.b(regtop_g_udb_cpu_r[1]));
   oa12s01 U271435 (.o(n186694),
	.a(n252278),
	.b(n252940),
	.c(n252285));
   na02s01 U271436 (.o(n252279),
	.a(n252283),
	.b(regtop_g_udb_cpu_r[2]));
   oa12s01 U271437 (.o(n186695),
	.a(n252279),
	.b(n252938),
	.c(n252285));
   in01f02 U271438 (.o(n253002),
	.a(regtop_g_wd_r[3]));
   na02s01 U271439 (.o(n252280),
	.a(regtop_g_udb_cpu_r[3]),
	.b(n252283));
   oa12s01 U271440 (.o(n186696),
	.a(n252280),
	.b(n253002),
	.c(n252285));
   in01s01 U271441 (.o(n252935),
	.a(regtop_g_wd_r[4]));
   na02s01 U271442 (.o(n252281),
	.a(regtop_g_udb_cpu_r[4]),
	.b(n252283));
   oa12s01 U271443 (.o(n186697),
	.a(n252281),
	.b(n252935),
	.c(n252285));
   in01f80 U271444 (.o(n252933),
	.a(regtop_g_wd_r[5]));
   na02s01 U271445 (.o(n252282),
	.a(regtop_g_udb_cpu_r[5]),
	.b(n252283));
   oa12s01 U271446 (.o(n186698),
	.a(n252282),
	.b(n252933),
	.c(n252285));
   in01f02 U271447 (.o(n252885),
	.a(regtop_g_wd_r[6]));
   na02s01 U271448 (.o(n252284),
	.a(regtop_g_udb_cpu_r[6]),
	.b(n252283));
   oa12s01 U271449 (.o(n186699),
	.a(n252284),
	.b(n252885),
	.c(n252285));
   no03s01 U271450 (.o(n186713),
	.a(n252953),
	.b(n252286),
	.c(n252829));
   in01s01 U271451 (.o(n186717),
	.a(n252287));
   oa12s01 U271452 (.o(n252290),
	.a(n252288),
	.b(n252289),
	.c(cntrltop_ctmg_ctpedet_c_bigpictdet_r));
   in01s01 U271453 (.o(n186718),
	.a(n252290));
   na02s01 U271454 (.o(n252292),
	.a(n252567),
	.b(n252363));
   in01s01 U271455 (.o(n252291),
	.a(regtop_g_fbst_r[1]));
   oa22s01 U271456 (.o(n186721),
	.a(FE_OFN494_n252377),
	.b(n252292),
	.c(n252305),
	.d(n252291));
   na02s01 U271457 (.o(n252294),
	.a(n252567),
	.b(n252674));
   oa22s01 U271458 (.o(n186722),
	.a(FE_OFN494_n252377),
	.b(n252294),
	.c(n252305),
	.d(n252293));
   in01s01 U271459 (.o(n252295),
	.a(regtop_g_fbst_r[4]));
   oa22s01 U271460 (.o(n186723),
	.a(FE_OFN494_n252377),
	.b(n252296),
	.c(n252305),
	.d(n252295));
   oa22s01 U271461 (.o(n186724),
	.a(FE_OFN494_n252377),
	.b(n252298),
	.c(n252305),
	.d(n252297));
   no02s01 U271462 (.o(n252301),
	.a(n252299),
	.b(FE_OFN494_n252377));
   in01s01 U271463 (.o(n186725),
	.a(n252303));
   in01s01 U271464 (.o(n252304),
	.a(regtop_g_fbst_r[7]));
   oa22s01 U271465 (.o(n186726),
	.a(FE_OFN494_n252377),
	.b(n252306),
	.c(n252305),
	.d(n252304));
   in01s01 U271466 (.o(n252311),
	.a(n252307));
   na02s01 U271467 (.o(n252310),
	.a(regtop_g_nferror_r),
	.b(n252377));
   oa22s01 U271468 (.o(n186732),
	.a(n252311),
	.b(n252310),
	.c(n252309),
	.d(n252308));
   in01s01 U271469 (.o(n252313),
	.a(regtop_g_fpst_r[0]));
   oa12s01 U271470 (.o(n211876),
	.a(n252312),
	.b(n252818),
	.c(n252313));
   oa22s01 U271471 (.o(n252315),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[1]),
	.c(regtop_g_tmc_r[1]),
	.d(n252339));
   in01s01 U271472 (.o(n211877),
	.a(n252315));
   oa22s01 U271473 (.o(n252316),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[2]),
	.c(regtop_g_tmc_r[2]),
	.d(n252339));
   in01s01 U271474 (.o(n211878),
	.a(n252316));
   oa22s01 U271475 (.o(n252317),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[3]),
	.c(regtop_g_tmc_r[3]),
	.d(n252339));
   in01s01 U271476 (.o(n211879),
	.a(n252317));
   oa22s01 U271477 (.o(n252318),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[4]),
	.c(regtop_g_tmc_r[4]),
	.d(n252339));
   oa22s01 U271478 (.o(n252319),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[5]),
	.c(regtop_g_tmc_r[5]),
	.d(n252339));
   in01s01 U271479 (.o(n211881),
	.a(n252319));
   oa22s01 U271480 (.o(n252320),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[6]),
	.c(regtop_g_tmc_r[6]),
	.d(n252339));
   in01s01 U271481 (.o(n211882),
	.a(n252320));
   oa22s01 U271482 (.o(n252321),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[7]),
	.c(regtop_g_tmc_r[7]),
	.d(n252339));
   in01s01 U271483 (.o(n211883),
	.a(n252321));
   oa22s01 U271484 (.o(n252322),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[8]),
	.c(regtop_g_tmc_r[8]),
	.d(n252339));
   in01s01 U271485 (.o(n211884),
	.a(n252322));
   oa22s01 U271486 (.o(n252323),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[9]),
	.c(regtop_g_tmc_r[9]),
	.d(n252339));
   in01s01 U271487 (.o(n211885),
	.a(n252323));
   oa22s01 U271488 (.o(n252324),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[10]),
	.c(regtop_g_tmc_r[10]),
	.d(n252339));
   in01s01 U271489 (.o(n211886),
	.a(n252324));
   oa22s01 U271490 (.o(n252325),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[11]),
	.c(regtop_g_tmc_r[11]),
	.d(n252339));
   in01s01 U271491 (.o(n211887),
	.a(n252325));
   oa22s01 U271492 (.o(n252326),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[13]),
	.c(regtop_g_tmc_r[12]),
	.d(n252339));
   in01s01 U271493 (.o(n211888),
	.a(n252326));
   oa22s01 U271494 (.o(n252327),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[14]),
	.c(regtop_g_tmc_r[13]),
	.d(n252339));
   in01s01 U271495 (.o(n211889),
	.a(n252327));
   oa22s01 U271496 (.o(n252328),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[15]),
	.c(regtop_g_tmc_r[14]),
	.d(n252339));
   in01s01 U271497 (.o(n211890),
	.a(n252328));
   oa22s01 U271498 (.o(n252329),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_tmc_r[15]),
	.d(n252339));
   in01s01 U271499 (.o(n211891),
	.a(n252329));
   oa22s01 U271500 (.o(n252330),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_tmc_r[16]),
	.d(n252339));
   in01s01 U271501 (.o(n211892),
	.a(n252330));
   oa22s01 U271502 (.o(n252331),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_tmc_r[17]),
	.d(n252339));
   in01s01 U271503 (.o(n211893),
	.a(n252331));
   oa22s01 U271504 (.o(n252332),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_tmc_r[18]),
	.d(n252339));
   in01s01 U271505 (.o(n211894),
	.a(n252332));
   oa22s01 U271506 (.o(n252333),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_tmc_r[19]),
	.d(n252339));
   oa22s01 U271507 (.o(n252334),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_tmc_r[20]),
	.d(n252339));
   in01s01 U271508 (.o(n211896),
	.a(n252334));
   oa22s01 U271509 (.o(n252335),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_tmc_r[21]),
	.d(n252339));
   in01s01 U271510 (.o(n211897),
	.a(n252335));
   oa22s01 U271511 (.o(n252336),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_tmc_r[22]),
	.d(n252339));
   in01s01 U271512 (.o(n211898),
	.a(n252336));
   oa22s01 U271513 (.o(n252337),
	.a(FE_OFN354_n252338),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_tmc_r[23]),
	.d(n252339));
   in01s01 U271514 (.o(n211899),
	.a(n252337));
   ao22s01 U271515 (.o(n252340),
	.a(n252339),
	.b(regtop_g_paramdata_r[0]),
	.c(regtop_g_tmc_r[0]),
	.d(FE_OFN354_n252338));
   in01s01 U271516 (.o(n211900),
	.a(n252340));
   oa22s01 U271517 (.o(n252342),
	.a(n252350),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_tc_r[1]),
	.d(n252349));
   in01s01 U271518 (.o(n211901),
	.a(n252342));
   oa22s01 U271519 (.o(n252343),
	.a(n252350),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_tc_r[2]),
	.d(n252349));
   in01s01 U271520 (.o(n211902),
	.a(n252343));
   oa22s01 U271521 (.o(n252344),
	.a(n252350),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_tc_r[3]),
	.d(n252349));
   in01s01 U271522 (.o(n211903),
	.a(n252344));
   oa22s01 U271523 (.o(n252345),
	.a(n252350),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_tc_r[4]),
	.d(n252349));
   in01s01 U271524 (.o(n211904),
	.a(n252345));
   oa22s01 U271525 (.o(n252346),
	.a(n252350),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_tc_r[5]),
	.d(n252349));
   in01s01 U271526 (.o(n211905),
	.a(n252346));
   oa22s01 U271527 (.o(n252347),
	.a(n252350),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_tc_r[6]),
	.d(n252349));
   in01s01 U271528 (.o(n211906),
	.a(n252347));
   oa22s01 U271529 (.o(n252348),
	.a(n252350),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_tc_r[7]),
	.d(n252349));
   in01s01 U271530 (.o(n211907),
	.a(n252348));
   oa22s01 U271531 (.o(n252351),
	.a(n252350),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_tc_r[0]),
	.d(n252349));
   in01s01 U271532 (.o(n211908),
	.a(n252351));
   oa22s01 U271533 (.o(n252353),
	.a(n252361),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_pali_r[1]),
	.d(n252360));
   in01s01 U271534 (.o(n211909),
	.a(n252353));
   oa22s01 U271535 (.o(n252354),
	.a(n252361),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_pali_r[2]),
	.d(n252360));
   oa22s01 U271536 (.o(n252355),
	.a(n252361),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_pali_r[3]),
	.d(n252360));
   in01s01 U271537 (.o(n211911),
	.a(n252355));
   oa22s01 U271538 (.o(n252356),
	.a(n252361),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_pali_r[4]),
	.d(n252360));
   in01s01 U271539 (.o(n211912),
	.a(n252356));
   oa22s01 U271540 (.o(n252357),
	.a(n252361),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_pali_r[5]),
	.d(n252360));
   in01s01 U271541 (.o(n211913),
	.a(n252357));
   oa22s01 U271542 (.o(n252358),
	.a(n252361),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_pali_r[6]),
	.d(n252360));
   in01s01 U271543 (.o(n211914),
	.a(n252358));
   oa22s01 U271544 (.o(n252359),
	.a(n252361),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_pali_r[7]),
	.d(n252360));
   in01s01 U271545 (.o(n211915),
	.a(n252359));
   oa22s01 U271546 (.o(n252362),
	.a(n252361),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_pali_r[0]),
	.d(n252360));
   in01s01 U271547 (.o(n211916),
	.a(n252362));
   in01s01 U271548 (.o(n252367),
	.a(regtop_g_fpst_r[4]));
   in01s01 U271549 (.o(n252364),
	.a(n252363));
   no02s01 U271550 (.o(n252365),
	.a(n252676),
	.b(n252364));
   in01s01 U271551 (.o(n252366),
	.a(n252365));
   in01s01 U271552 (.o(n211963),
	.a(n252369));
   in01s01 U271553 (.o(n252370),
	.a(regtop_g_nfst_r[17]));
   oa22s01 U271554 (.o(n211964),
	.a(FE_OFN494_n252377),
	.b(n252371),
	.c(n252370),
	.d(n252824));
   in01s01 U271555 (.o(n211965),
	.a(n252373));
   in01s01 U271556 (.o(n211967),
	.a(n252375));
   in01s01 U271557 (.o(n211968),
	.a(n252378));
   in01s01 U271558 (.o(n211969),
	.a(n252385));
   in01s01 U271559 (.o(n211970),
	.a(n252386));
   in01s01 U271560 (.o(n211971),
	.a(n252387));
   in01s01 U271561 (.o(n211972),
	.a(n252388));
   in01s01 U271562 (.o(n211973),
	.a(n252389));
   in01s01 U271563 (.o(n211974),
	.a(n252390));
   in01s01 U271564 (.o(n211975),
	.a(n252391));
   in01s01 U271565 (.o(n211976),
	.a(n252392));
   oa22s01 U271566 (.o(n252393),
	.a(n252401),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_fcho2_r[9]),
	.d(n252400));
   ao22s01 U271567 (.o(n211978),
	.a(n252400),
	.b(n252660),
	.c(n252394),
	.d(n252401));
   ao22s01 U271568 (.o(n211979),
	.a(n252400),
	.b(n252662),
	.c(n252395),
	.d(n252401));
   in01s01 U271569 (.o(n211980),
	.a(n252396));
   in01s01 U271570 (.o(n211981),
	.a(n252397));
   in01s01 U271571 (.o(n211982),
	.a(n252398));
   in01s01 U271572 (.o(n211983),
	.a(n252399));
   in01s01 U271573 (.o(n211984),
	.a(n252402));
   na03f01 U271574 (.o(n252405),
	.a(regtop_g_paramadr_r[3]),
	.b(regtop_g_paramadr_r[4]),
	.c(n252404));
   in01s01 U271575 (.o(n211985),
	.a(n252406));
   in01s01 U271576 (.o(n211986),
	.a(n252407));
   in01s01 U271577 (.o(n211987),
	.a(n252408));
   in01s01 U271578 (.o(n211988),
	.a(n252409));
   in01s01 U271579 (.o(n211989),
	.a(n252410));
   in01s01 U271580 (.o(n211990),
	.a(n252411));
   in01s01 U271581 (.o(n211991),
	.a(n252412));
   oa22s01 U271582 (.o(n252413),
	.a(FE_OFN212_n252422),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_fcho0_r[8]),
	.d(n252421));
   in01s01 U271583 (.o(n211993),
	.a(n252414));
   in01s01 U271584 (.o(n211994),
	.a(n252415));
   in01s01 U271585 (.o(n211995),
	.a(n252416));
   ao22s01 U271586 (.o(n211996),
	.a(n252421),
	.b(n252664),
	.c(n252417),
	.d(FE_OFN212_n252422));
   ao22s01 U271587 (.o(n211997),
	.a(n252421),
	.b(n252666),
	.c(n252418),
	.d(FE_OFN212_n252422));
   in01s01 U271588 (.o(n211998),
	.a(n252419));
   in01s01 U271589 (.o(n211999),
	.a(n252420));
   in01s01 U271590 (.o(n212000),
	.a(n252423));
   oa22s01 U271591 (.o(n252426),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_va_r),
	.d(n252445));
   in01s01 U271592 (.o(n212001),
	.a(n252426));
   oa22s01 U271593 (.o(n252427),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_fs_r[0]),
	.d(n252445));
   in01s01 U271594 (.o(n212002),
	.a(n252427));
   oa22s01 U271595 (.o(n252428),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_fs_r[2]),
	.d(n252445));
   in01s01 U271596 (.o(n212003),
	.a(n252428));
   oa22s01 U271597 (.o(n252429),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_fs_r[1]),
	.d(n252445));
   in01s01 U271598 (.o(n212004),
	.a(n252429));
   oa22s01 U271599 (.o(n252430),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_sc_r),
	.d(n252445));
   in01s01 U271600 (.o(n212005),
	.a(n252430));
   oa22s01 U271601 (.o(n252431),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[13]),
	.c(regtop_g_ba_r[0]),
	.d(n252445));
   in01s01 U271602 (.o(n212006),
	.a(n252431));
   oa22s01 U271603 (.o(n252432),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_ba_r[6]),
	.d(n252445));
   oa22s01 U271604 (.o(n252433),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_ba_r[5]),
	.d(n252445));
   in01s01 U271605 (.o(n212008),
	.a(n252433));
   oa22s01 U271606 (.o(n252434),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_ba_r[4]),
	.d(n252445));
   in01s01 U271607 (.o(n212009),
	.a(n252434));
   oa22s01 U271608 (.o(n252435),
	.a(n252446),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_ba_r[3]),
	.d(n252445));
   in01s01 U271609 (.o(n212010),
	.a(n252435));
   oa22s01 U271610 (.o(n252436),
	.a(n252446),
	.b(regtop_g_paramdata_r[15]),
	.c(regtop_g_ba_r[2]),
	.d(n252445));
   in01s01 U271611 (.o(n212011),
	.a(n252436));
   oa22s01 U271612 (.o(n252437),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[14]),
	.c(regtop_g_ba_r[1]),
	.d(n252445));
   in01s01 U271613 (.o(n212012),
	.a(n252437));
   oa22s01 U271614 (.o(n252438),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[6]),
	.c(regtop_g_scp_r[1]),
	.d(n252445));
   in01s01 U271615 (.o(n212013),
	.a(n252438));
   oa22s01 U271616 (.o(n252439),
	.a(n252446),
	.b(regtop_g_paramdata_r[7]),
	.c(regtop_g_scp_r[2]),
	.d(n252445));
   in01s01 U271617 (.o(n212014),
	.a(n252439));
   oa22s01 U271618 (.o(n252440),
	.a(n252446),
	.b(regtop_g_paramdata_r[8]),
	.c(regtop_g_scp_r[3]),
	.d(n252445));
   in01s01 U271619 (.o(n212015),
	.a(n252440));
   oa22s01 U271620 (.o(n252441),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[9]),
	.c(regtop_g_scp_r[4]),
	.d(n252445));
   in01s01 U271621 (.o(n212016),
	.a(n252441));
   oa22s01 U271622 (.o(n252442),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[10]),
	.c(regtop_g_scp_r[5]),
	.d(n252445));
   in01s01 U271623 (.o(n212017),
	.a(n252442));
   oa22s01 U271624 (.o(n252443),
	.a(n252446),
	.b(regtop_g_paramdata_r[11]),
	.c(regtop_g_scp_r[6]),
	.d(n252445));
   in01s01 U271625 (.o(n212018),
	.a(n252443));
   oa22s01 U271626 (.o(n252444),
	.a(n252446),
	.b(regtop_g_paramdata_r[12]),
	.c(regtop_g_scp_r[7]),
	.d(n252445));
   in01s01 U271627 (.o(n212019),
	.a(n252444));
   oa22s01 U271628 (.o(n252447),
	.a(FE_OFN37_n252446),
	.b(regtop_g_paramdata_r[5]),
	.c(regtop_g_scp_r[0]),
	.d(n252445));
   in01s01 U271629 (.o(n212020),
	.a(n252447));
   in01s01 U271630 (.o(n212021),
	.a(n252450));
   oa22s01 U271631 (.o(n252451),
	.a(n252460),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_tr_r[2]),
	.d(n252459));
   in01s01 U271632 (.o(n212023),
	.a(n252452));
   in01s01 U271633 (.o(n212024),
	.a(n252453));
   in01s01 U271634 (.o(n212025),
	.a(n252454));
   in01s01 U271635 (.o(n212026),
	.a(n252455));
   in01s01 U271636 (.o(n212027),
	.a(n252456));
   in01s01 U271637 (.o(n212028),
	.a(n252457));
   in01s01 U271638 (.o(n212029),
	.a(n252458));
   in01s01 U271639 (.o(n212030),
	.a(n252461));
   oa22s01 U271640 (.o(n252465),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[8]),
	.c(regtop_g_brv_r[1]),
	.d(n252482));
   in01s01 U271641 (.o(n212031),
	.a(n252465));
   oa22s01 U271642 (.o(n252466),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[9]),
	.c(regtop_g_brv_r[2]),
	.d(n252482));
   in01s01 U271643 (.o(n212032),
	.a(n252466));
   oa22s01 U271644 (.o(n252467),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[10]),
	.c(regtop_g_brv_r[3]),
	.d(n252482));
   in01s01 U271645 (.o(n212033),
	.a(n252467));
   oa22s01 U271646 (.o(n252468),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[11]),
	.c(regtop_g_brv_r[4]),
	.d(n252482));
   in01s01 U271647 (.o(n212034),
	.a(n252468));
   oa22s01 U271648 (.o(n252469),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[12]),
	.c(regtop_g_brv_r[5]),
	.d(n252482));
   in01s01 U271649 (.o(n212035),
	.a(n252469));
   oa22s01 U271650 (.o(n252470),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[13]),
	.c(regtop_g_brv_r[6]),
	.d(n252482));
   in01s01 U271651 (.o(n212036),
	.a(n252470));
   oa22s01 U271652 (.o(n252471),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[14]),
	.c(regtop_g_brv_r[7]),
	.d(n252482));
   oa22s01 U271653 (.o(n252472),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[15]),
	.c(regtop_g_brv_r[8]),
	.d(n252482));
   in01s01 U271654 (.o(n212038),
	.a(n252472));
   oa22s01 U271655 (.o(n252473),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_brv_r[9]),
	.d(n252482));
   in01s01 U271656 (.o(n212039),
	.a(n252473));
   oa22s01 U271657 (.o(n252474),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_brv_r[10]),
	.d(n252482));
   in01s01 U271658 (.o(n212040),
	.a(n252474));
   oa22s01 U271659 (.o(n252475),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_brv_r[11]),
	.d(n252482));
   in01s01 U271660 (.o(n212041),
	.a(n252475));
   oa22s01 U271661 (.o(n252476),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_brv_r[12]),
	.d(n252482));
   in01s01 U271662 (.o(n212042),
	.a(n252476));
   oa22s01 U271663 (.o(n252477),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_brv_r[13]),
	.d(n252482));
   in01s01 U271664 (.o(n212043),
	.a(n252477));
   oa22s01 U271665 (.o(n252478),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_brv_r[14]),
	.d(n252482));
   in01s01 U271666 (.o(n212044),
	.a(n252478));
   oa22s01 U271667 (.o(n252479),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_brv_r[15]),
	.d(n252482));
   in01s01 U271668 (.o(n212045),
	.a(n252479));
   oa22s01 U271669 (.o(n252480),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_brv_r[16]),
	.d(n252482));
   in01s01 U271670 (.o(n212046),
	.a(n252480));
   oa22s01 U271671 (.o(n252481),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_brv_r[17]),
	.d(n252482));
   in01s01 U271672 (.o(n212047),
	.a(n252481));
   oa22s01 U271673 (.o(n252484),
	.a(FE_OFN214_n252483),
	.b(regtop_g_paramdata_r[7]),
	.c(regtop_g_brv_r[0]),
	.d(n252482));
   in01s01 U271674 (.o(n212048),
	.a(n252484));
   in01s01 U271675 (.o(n252486),
	.a(regtop_g_nfst_r[8]));
   oa22s01 U271676 (.o(n212056),
	.a(FE_OFN494_n252377),
	.b(n252487),
	.c(n252486),
	.d(n252824));
   in01s01 U271677 (.o(n252488),
	.a(regtop_g_nfst_r[5]));
   oa22s01 U271678 (.o(n212057),
	.a(FE_OFN494_n252377),
	.b(n252489),
	.c(n252824),
	.d(n252488));
   in01s01 U271679 (.o(n252490),
	.a(regtop_g_nfst_r[0]));
   oa22s01 U271680 (.o(n212058),
	.a(FE_OFN494_n252377),
	.b(n252491),
	.c(n252824),
	.d(n252490));
   in01s01 U271681 (.o(n212059),
	.a(n252492));
   in01s01 U271682 (.o(n212060),
	.a(n252493));
   in01s01 U271683 (.o(n212061),
	.a(n252494));
   in01s01 U271684 (.o(n212062),
	.a(n252495));
   in01s01 U271685 (.o(n212063),
	.a(n252496));
   in01s01 U271686 (.o(n212064),
	.a(n252497));
   in01s01 U271687 (.o(n212065),
	.a(n252498));
   in01s01 U271688 (.o(n212066),
	.a(n252499));
   oa22s01 U271689 (.o(n252500),
	.a(FE_OFN356_n252508),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_fcho1_r[9]),
	.d(n252507));
   ao22s01 U271690 (.o(n212068),
	.a(n252507),
	.b(n252660),
	.c(n252501),
	.d(FE_OFN356_n252508));
   in01s01 U271691 (.o(n212069),
	.a(n252502));
   in01s01 U271692 (.o(n212070),
	.a(n252503));
   ao22s01 U271693 (.o(n212071),
	.a(n252507),
	.b(n252666),
	.c(n252504),
	.d(FE_OFN356_n252508));
   in01s01 U271694 (.o(n212072),
	.a(n252505));
   in01s01 U271695 (.o(n212073),
	.a(n252506));
   in01s01 U271696 (.o(n212074),
	.a(n252509));
   no02f02 U271697 (.o(n252512),
	.a(n252575),
	.b(n252510));
   in01s01 U271698 (.o(n252513),
	.a(n252512));
   na02s01 U271699 (.o(n252511),
	.a(n252513),
	.b(regtop_g_nfco_r[1]));
   oa12s01 U271700 (.o(n212075),
	.a(n252511),
	.b(n252755),
	.c(n252513));
   oa22s01 U271701 (.o(n252514),
	.a(n252513),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_nfco_r[0]),
	.d(n252512));
   in01s01 U271702 (.o(n212076),
	.a(n252514));
   na02s01 U271703 (.o(n252516),
	.a(regtop_g_paramadr_r[6]),
	.b(n252515));
   na02s01 U271704 (.o(n252518),
	.a(n252521),
	.b(regtop_g_tff_r));
   oa12s01 U271705 (.o(n212077),
	.a(n252518),
	.b(n252755),
	.c(n252521));
   in01s01 U271706 (.o(n252520),
	.a(n252521));
   oa22s01 U271707 (.o(n252519),
	.a(n252521),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_rff_r),
	.d(n252520));
   in01s01 U271708 (.o(n212078),
	.a(n252519));
   oa22s01 U271709 (.o(n252522),
	.a(n252521),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_pf_r),
	.d(n252520));
   in01s01 U271710 (.o(n212079),
	.a(n252522));
   in01s01 U271711 (.o(n212080),
	.a(n252524));
   in01s01 U271712 (.o(n212081),
	.a(n252525));
   oa22s01 U271713 (.o(n252526),
	.a(n252540),
	.b(regtop_g_paramdata_r[12]),
	.c(regtop_g_vd_r[3]),
	.d(FE_OFN508_n252540));
   in01s01 U271714 (.o(n212083),
	.a(n252527));
   in01s01 U271715 (.o(n212084),
	.a(n252528));
   in01s01 U271716 (.o(n212085),
	.a(n252529));
   in01s01 U271717 (.o(n212086),
	.a(n252530));
   in01s01 U271718 (.o(n212087),
	.a(n252531));
   in01s01 U271719 (.o(n212088),
	.a(n252532));
   in01s01 U271720 (.o(n212089),
	.a(n252533));
   in01s01 U271721 (.o(n212090),
	.a(n252534));
   in01s01 U271722 (.o(n212091),
	.a(n252535));
   in01s01 U271723 (.o(n212092),
	.a(n252536));
   in01s01 U271724 (.o(n212093),
	.a(n252537));
   in01s01 U271725 (.o(n212094),
	.a(n252538));
   in01s01 U271726 (.o(n212095),
	.a(n252541));
   no02s01 U271727 (.o(n252543),
	.a(n252542),
	.b(n252575));
   na02f01 U271728 (.o(n252545),
	.a(n252687),
	.b(n252543));
   na02s01 U271729 (.o(n252544),
	.a(n252545),
	.b(regtop_g_cpf_r));
   oa12s01 U271730 (.o(n212096),
	.a(n252544),
	.b(n252755),
	.c(n252545));
   in01s01 U271731 (.o(n252546),
	.a(regtop_g_nfst_r[15]));
   oa22s01 U271732 (.o(n212097),
	.a(FE_OFN494_n252377),
	.b(n252547),
	.c(n252824),
	.d(n252546));
   in01s01 U271733 (.o(n252548),
	.a(regtop_g_dhs_r[1]));
   ao22s01 U271734 (.o(n212122),
	.a(n252563),
	.b(n252646),
	.c(n252548),
	.d(n252561));
   in01s01 U271735 (.o(n252549),
	.a(regtop_g_dhs_r[2]));
   ao22s01 U271736 (.o(n212123),
	.a(n252563),
	.b(n252648),
	.c(n252549),
	.d(n252561));
   in01s01 U271737 (.o(n252550),
	.a(regtop_g_dhs_r[3]));
   ao22s01 U271738 (.o(n212124),
	.a(n252563),
	.b(n252650),
	.c(n252550),
	.d(n252561));
   in01s01 U271739 (.o(n252551),
	.a(regtop_g_dhs_r[4]));
   ao22s01 U271740 (.o(n212125),
	.a(n252563),
	.b(n252652),
	.c(n252551),
	.d(n252561));
   in01s01 U271741 (.o(n252552),
	.a(regtop_g_dhs_r[5]));
   ao22s01 U271742 (.o(n212126),
	.a(n252563),
	.b(n252654),
	.c(n252552),
	.d(n252561));
   in01s01 U271743 (.o(n252553),
	.a(regtop_g_dhs_r[6]));
   in01s01 U271744 (.o(n252554),
	.a(regtop_g_dhs_r[7]));
   ao22s01 U271745 (.o(n212128),
	.a(n252563),
	.b(n252658),
	.c(n252554),
	.d(n252561));
   in01s01 U271746 (.o(n252555),
	.a(regtop_g_dhs_r[8]));
   ao22s01 U271747 (.o(n212129),
	.a(n252563),
	.b(n252660),
	.c(n252555),
	.d(n252561));
   in01s01 U271748 (.o(n252556),
	.a(regtop_g_dhs_r[9]));
   ao22s01 U271749 (.o(n212130),
	.a(n252563),
	.b(n252662),
	.c(n252556),
	.d(n252561));
   in01s01 U271750 (.o(n252557),
	.a(regtop_g_dhs_r[10]));
   ao22s01 U271751 (.o(n212131),
	.a(n252563),
	.b(n252664),
	.c(n252557),
	.d(n252561));
   ao22s01 U271752 (.o(n212132),
	.a(n252563),
	.b(n252666),
	.c(n252558),
	.d(n252561));
   in01s01 U271753 (.o(n252559),
	.a(regtop_g_dhs_r[12]));
   ao22s01 U271754 (.o(n212133),
	.a(n252563),
	.b(n252778),
	.c(n252559),
	.d(n252561));
   in01s01 U271755 (.o(n252560),
	.a(regtop_g_dhs_r[13]));
   ao22s01 U271756 (.o(n212134),
	.a(n252563),
	.b(n252755),
	.c(n252560),
	.d(n252561));
   in01s01 U271757 (.o(n252562),
	.a(regtop_g_dhs_r[0]));
   ao22s01 U271758 (.o(n212135),
	.a(n252563),
	.b(n252644),
	.c(n252562),
	.d(n252561));
   na02f02 U271759 (.o(n252566),
	.a(n252568),
	.b(n252758));
   na02s01 U271760 (.o(n252565),
	.a(n252566),
	.b(regtop_g_cd_r));
   oa12s01 U271761 (.o(n212136),
	.a(n252565),
	.b(n252755),
	.c(n252566));
   na02s01 U271762 (.o(n252569),
	.a(n252571),
	.b(regtop_g_cf_r[1]));
   oa12s01 U271763 (.o(n212137),
	.a(n252569),
	.b(n252755),
	.c(n252571));
   oa22s01 U271764 (.o(n252572),
	.a(n252571),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_cf_r[0]),
	.d(n252570));
   in01s01 U271765 (.o(n212138),
	.a(n252572));
   in01s01 U271766 (.o(n252585),
	.a(regtop_g_adb_r[4]));
   na02s01 U271767 (.o(n252573),
	.a(regtop_g_adb_r[2]),
	.b(n252591));
   in01s01 U271768 (.o(n252594),
	.a(n252573));
   na02s01 U271769 (.o(n252588),
	.a(regtop_g_adb_r[3]),
	.b(n252594));
   no02s01 U271770 (.o(n252587),
	.a(n252585),
	.b(n252588));
   na02s01 U271771 (.o(n252581),
	.a(regtop_g_adb_r[5]),
	.b(n252587));
   in01s01 U271772 (.o(n252577),
	.a(n252602));
   na02s01 U271773 (.o(n252578),
	.a(n252595),
	.b(n252579));
   in01s01 U271774 (.o(n252583),
	.a(regtop_g_adb_r[5]));
   oa12s01 U271775 (.o(n252582),
	.a(n252581),
	.b(regtop_g_adb_r[5]),
	.c(n252587));
   oa22s01 U271776 (.o(n212148),
	.a(n252583),
	.b(n252602),
	.c(n252601),
	.d(n252582));
   ao12s01 U271777 (.o(n252584),
	.a(n252601),
	.b(n252585),
	.c(n252588));
   in01s01 U271778 (.o(n252586),
	.a(n252584));
   oa22s01 U271779 (.o(n212149),
	.a(n252587),
	.b(n252586),
	.c(n252585),
	.d(n252602));
   in01s01 U271780 (.o(n252590),
	.a(regtop_g_adb_r[3]));
   oa12s01 U271781 (.o(n252589),
	.a(n252588),
	.b(regtop_g_adb_r[3]),
	.c(n252594));
   oa22s01 U271782 (.o(n212150),
	.a(n252590),
	.b(n252602),
	.c(n252601),
	.d(n252589));
   oa12s01 U271783 (.o(n252593),
	.a(n252595),
	.b(regtop_g_adb_r[2]),
	.c(n252591));
   in01s01 U271784 (.o(n252592),
	.a(regtop_g_adb_r[2]));
   oa22s01 U271785 (.o(n212151),
	.a(n252594),
	.b(n252593),
	.c(n252592),
	.d(n252602));
   oa12s01 U271786 (.o(n252598),
	.a(n252595),
	.b(n252597),
	.c(n252596));
   oa12s01 U271787 (.o(n212152),
	.a(n252598),
	.b(n252602),
	.c(n252599));
   ao22s01 U271788 (.o(n212153),
	.a(regtop_g_adb_r[0]),
	.b(n252602),
	.c(n252601),
	.d(n252600));
   in01s01 U271789 (.o(n252603),
	.a(regtop_g_nfst_r[10]));
   oa22s01 U271790 (.o(n212154),
	.a(FE_OFN494_n252377),
	.b(n252604),
	.c(n252824),
	.d(n252603));
   in01s01 U271791 (.o(n252605),
	.a(regtop_g_nfst_r[18]));
   oa22s01 U271792 (.o(n212155),
	.a(n252606),
	.b(FE_OFN494_n252377),
	.c(n252824),
	.d(n252605));
   in01s01 U271793 (.o(n252607),
	.a(regtop_g_nfst_r[12]));
   oa22s01 U271794 (.o(n212156),
	.a(n252608),
	.b(FE_OFN494_n252377),
	.c(n252824),
	.d(n252607));
   na02s01 U271795 (.o(n252610),
	.a(n252613),
	.b(n252730));
   na02s01 U271796 (.o(n252609),
	.a(n252610),
	.b(regtop_g_mpeg_r));
   oa12s01 U271797 (.o(n212157),
	.a(n252609),
	.b(n252755),
	.c(n252610));
   na02f03 U271798 (.o(n252612),
	.a(n252706),
	.b(n252613));
   na02s01 U271799 (.o(n252611),
	.a(n252612),
	.b(regtop_g_cdf_r));
   oa12s01 U271800 (.o(n212158),
	.a(n252611),
	.b(n252755),
	.c(n252612));
   in01s01 U271801 (.o(n212159),
	.a(n252614));
   in01s01 U271802 (.o(n212160),
	.a(n252615));
   in01s01 U271803 (.o(n212161),
	.a(n252616));
   in01s01 U271804 (.o(n212162),
	.a(n252617));
   in01s01 U271805 (.o(n212163),
	.a(n252618));
   in01s01 U271806 (.o(n212164),
	.a(n252619));
   in01s01 U271807 (.o(n212165),
	.a(n252620));
   in01s01 U271808 (.o(n212166),
	.a(n252621));
   in01s01 U271809 (.o(n212167),
	.a(n252622));
   in01s01 U271810 (.o(n212168),
	.a(n252623));
   in01s01 U271811 (.o(n212169),
	.a(n252624));
   in01s01 U271812 (.o(n212170),
	.a(n252625));
   in01s01 U271813 (.o(n212171),
	.a(n252626));
   oa22s01 U271814 (.o(n252627),
	.a(FE_OFN558_n252630),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_fcvo1_r[14]),
	.d(n252629));
   in01s01 U271815 (.o(n212173),
	.a(n252628));
   in01s01 U271816 (.o(n212174),
	.a(n252631));
   oa22s01 U271817 (.o(n252632),
	.a(FE_OFN41_n252640),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_cp_r[1]),
	.d(n252639));
   in01s01 U271818 (.o(n212176),
	.a(n252632));
   oa22s01 U271819 (.o(n252633),
	.a(FE_OFN41_n252640),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_cp_r[2]),
	.d(n252639));
   in01s01 U271820 (.o(n212177),
	.a(n252633));
   oa22s01 U271821 (.o(n252634),
	.a(FE_OFN41_n252640),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_cp_r[3]),
	.d(n252639));
   in01s01 U271822 (.o(n212178),
	.a(n252634));
   oa22s01 U271823 (.o(n252635),
	.a(FE_OFN41_n252640),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_cp_r[4]),
	.d(n252639));
   in01s01 U271824 (.o(n212179),
	.a(n252635));
   oa22s01 U271825 (.o(n252636),
	.a(FE_OFN41_n252640),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_cp_r[5]),
	.d(n252639));
   in01s01 U271826 (.o(n212180),
	.a(n252636));
   oa22s01 U271827 (.o(n252637),
	.a(FE_OFN41_n252640),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_cp_r[6]),
	.d(n252639));
   in01s01 U271828 (.o(n212181),
	.a(n252637));
   oa22s01 U271829 (.o(n252638),
	.a(FE_OFN41_n252640),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_cp_r[7]),
	.d(n252639));
   in01s01 U271830 (.o(n212182),
	.a(n252638));
   oa22s01 U271831 (.o(n252641),
	.a(FE_OFN41_n252640),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_cp_r[0]),
	.d(n252639));
   in01s01 U271832 (.o(n212183),
	.a(n252641));
   in01s01 U271833 (.o(n252643),
	.a(regtop_g_dvs_r[1]));
   ao22s01 U271834 (.o(n212184),
	.a(n252671),
	.b(n252644),
	.c(n252643),
	.d(FE_OFN43_n252668));
   in01s01 U271835 (.o(n252645),
	.a(regtop_g_dvs_r[2]));
   ao22s01 U271836 (.o(n212185),
	.a(n252671),
	.b(n252646),
	.c(n252645),
	.d(FE_OFN43_n252668));
   in01s01 U271837 (.o(n252647),
	.a(regtop_g_dvs_r[3]));
   ao22s01 U271838 (.o(n212186),
	.a(n252671),
	.b(n252648),
	.c(n252647),
	.d(FE_OFN43_n252668));
   in01s01 U271839 (.o(n252651),
	.a(regtop_g_dvs_r[5]));
   ao22s01 U271840 (.o(n212188),
	.a(n252671),
	.b(n252652),
	.c(n252651),
	.d(FE_OFN43_n252668));
   in01s01 U271841 (.o(n252653),
	.a(regtop_g_dvs_r[6]));
   ao22s01 U271842 (.o(n212189),
	.a(n252671),
	.b(n252654),
	.c(n252653),
	.d(FE_OFN43_n252668));
   in01s01 U271843 (.o(n252655),
	.a(regtop_g_dvs_r[7]));
   ao22s01 U271844 (.o(n212190),
	.a(n252671),
	.b(n252656),
	.c(n252655),
	.d(FE_OFN43_n252668));
   in01s01 U271845 (.o(n252657),
	.a(regtop_g_dvs_r[8]));
   ao22s01 U271846 (.o(n212191),
	.a(n252671),
	.b(n252658),
	.c(n252657),
	.d(FE_OFN43_n252668));
   in01s01 U271847 (.o(n252659),
	.a(regtop_g_dvs_r[9]));
   ao22s01 U271848 (.o(n212192),
	.a(n252671),
	.b(n252660),
	.c(n252659),
	.d(FE_OFN43_n252668));
   in01s01 U271849 (.o(n252661),
	.a(regtop_g_dvs_r[10]));
   ao22s01 U271850 (.o(n212193),
	.a(n252671),
	.b(n252662),
	.c(n252661),
	.d(FE_OFN43_n252668));
   in01s01 U271851 (.o(n252663),
	.a(regtop_g_dvs_r[11]));
   ao22s01 U271852 (.o(n212194),
	.a(n252671),
	.b(n252664),
	.c(n252663),
	.d(FE_OFN43_n252668));
   in01s01 U271853 (.o(n252665),
	.a(regtop_g_dvs_r[12]));
   ao22s01 U271854 (.o(n212195),
	.a(n252671),
	.b(n252666),
	.c(n252665),
	.d(FE_OFN43_n252668));
   in01s01 U271855 (.o(n252667),
	.a(regtop_g_dvs_r[13]));
   ao22s01 U271856 (.o(n212196),
	.a(n252671),
	.b(n252778),
	.c(n252667),
	.d(FE_OFN43_n252668));
   in01s01 U271857 (.o(n252669),
	.a(regtop_g_dvs_r[0]));
   ao22s01 U271858 (.o(n212197),
	.a(n252671),
	.b(n252670),
	.c(n252669),
	.d(FE_OFN43_n252668));
   in01s01 U271859 (.o(n252672),
	.a(regtop_g_nfst_r[16]));
   oa22s01 U271860 (.o(n212198),
	.a(n252673),
	.b(FE_OFN494_n252377),
	.c(n252824),
	.d(n252672));
   in01s01 U271861 (.o(n252679),
	.a(regtop_g_fpst_r[5]));
   in01s01 U271862 (.o(n252675),
	.a(n252674));
   no02s01 U271863 (.o(n252677),
	.a(n252676),
	.b(n252675));
   in01s01 U271864 (.o(n252678),
	.a(n252677));
   oa12s01 U271865 (.o(n212199),
	.a(n252678),
	.b(n252818),
	.c(n252679));
   in01s01 U271866 (.o(n252683),
	.a(n252680));
   in01s01 U271867 (.o(n252681),
	.a(regtop_g_nfst_r[7]));
   oa22s01 U271868 (.o(n212200),
	.a(n252683),
	.b(n252682),
	.c(n252824),
	.d(n252681));
   in01s01 U271869 (.o(n252686),
	.a(n252685));
   oa22s01 U271870 (.o(n252688),
	.a(n252698),
	.b(regtop_g_paramdata_r[15]),
	.c(regtop_g_vbsv_r[1]),
	.d(n252697));
   oa22s01 U271871 (.o(n252689),
	.a(n252698),
	.b(regtop_g_paramdata_r[16]),
	.c(regtop_g_vbsv_r[2]),
	.d(n252697));
   in01s01 U271872 (.o(n212203),
	.a(n252689));
   oa22s01 U271873 (.o(n252690),
	.a(n252698),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_vbsv_r[3]),
	.d(n252697));
   in01s01 U271874 (.o(n212204),
	.a(n252690));
   oa22s01 U271875 (.o(n252691),
	.a(n252698),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_vbsv_r[4]),
	.d(n252697));
   in01s01 U271876 (.o(n212205),
	.a(n252691));
   oa22s01 U271877 (.o(n252692),
	.a(n252698),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_vbsv_r[5]),
	.d(n252697));
   in01s01 U271878 (.o(n212206),
	.a(n252692));
   oa22s01 U271879 (.o(n252693),
	.a(n252698),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_vbsv_r[6]),
	.d(n252697));
   in01s01 U271880 (.o(n212207),
	.a(n252693));
   oa22s01 U271881 (.o(n252694),
	.a(n252698),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_vbsv_r[7]),
	.d(n252697));
   in01s01 U271882 (.o(n212208),
	.a(n252694));
   oa22s01 U271883 (.o(n252695),
	.a(n252698),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_vbsv_r[8]),
	.d(n252697));
   in01s01 U271884 (.o(n212209),
	.a(n252695));
   oa22s01 U271885 (.o(n252696),
	.a(n252698),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_vbsv_r[9]),
	.d(n252697));
   in01s01 U271886 (.o(n212210),
	.a(n252696));
   oa22s01 U271887 (.o(n252699),
	.a(n252698),
	.b(regtop_g_paramdata_r[14]),
	.c(regtop_g_vbsv_r[0]),
	.d(n252697));
   in01s01 U271888 (.o(n212211),
	.a(n252699));
   in01s01 U271889 (.o(n252703),
	.a(n252704));
   in01s01 U271890 (.o(n212212),
	.a(n252701));
   in01s01 U271891 (.o(n212213),
	.a(n252702));
   in01s01 U271892 (.o(n212214),
	.a(n252705));
   na02s01 U271893 (.o(n252707),
	.a(n252709),
	.b(regtop_g_pis_r[1]));
   oa12s01 U271894 (.o(n212215),
	.a(n252707),
	.b(n252755),
	.c(n252709));
   in01s01 U271895 (.o(n252708),
	.a(n252709));
   oa22s01 U271896 (.o(n252710),
	.a(n252709),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_pis_r[0]),
	.d(n252708));
   in01s01 U271897 (.o(n212216),
	.a(n252710));
   oa22s01 U271898 (.o(n252712),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[10]),
	.c(regtop_g_fcvo0_r[1]),
	.d(n252727));
   in01s01 U271899 (.o(n212218),
	.a(n252713));
   in01s01 U271900 (.o(n212219),
	.a(n252714));
   in01s01 U271901 (.o(n212220),
	.a(n252715));
   in01s01 U271902 (.o(n212221),
	.a(n252716));
   in01s01 U271903 (.o(n212222),
	.a(n252717));
   in01s01 U271904 (.o(n212223),
	.a(n252718));
   in01s01 U271905 (.o(n212224),
	.a(n252719));
   in01s01 U271906 (.o(n212225),
	.a(n252720));
   in01s01 U271907 (.o(n212226),
	.a(n252721));
   in01s01 U271908 (.o(n212227),
	.a(n252722));
   in01s01 U271909 (.o(n212228),
	.a(n252723));
   in01s01 U271910 (.o(n212229),
	.a(n252724));
   in01s01 U271911 (.o(n212230),
	.a(n252725));
   in01s01 U271912 (.o(n212231),
	.a(n252726));
   oa22s01 U271913 (.o(n252729),
	.a(FE_OFN360_n252728),
	.b(regtop_g_paramdata_r[9]),
	.c(regtop_g_fcvo0_r[0]),
	.d(n252727));
   in01s01 U271914 (.o(n212233),
	.a(n252732));
   in01s01 U271915 (.o(n212234),
	.a(n252733));
   in01s01 U271916 (.o(n212235),
	.a(n252734));
   in01s01 U271917 (.o(n212236),
	.a(n252735));
   in01s01 U271918 (.o(n212237),
	.a(n252736));
   in01s01 U271919 (.o(n212238),
	.a(n252737));
   in01s01 U271920 (.o(n212239),
	.a(n252738));
   in01s01 U271921 (.o(n212240),
	.a(n252739));
   in01s01 U271922 (.o(n212241),
	.a(n252740));
   in01s01 U271923 (.o(n212242),
	.a(n252741));
   in01s01 U271924 (.o(n212243),
	.a(n252742));
   in01s01 U271925 (.o(n212244),
	.a(n252743));
   in01s01 U271926 (.o(n212245),
	.a(n252744));
   in01s01 U271927 (.o(n212246),
	.a(n252745));
   oa22s01 U271928 (.o(n252746),
	.a(FE_OFN362_n252748),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_fcvo2_r[15]),
	.d(n252747));
   in01s01 U271929 (.o(n212248),
	.a(n252749));
   oa12s01 U271930 (.o(n212249),
	.a(n252750),
	.b(n252818),
	.c(n252751));
   no02f02 U271931 (.o(n252756),
	.a(n252757),
	.b(n252752));
   in01s01 U271932 (.o(n252754),
	.a(regtop_g_ps_r));
   in01s01 U271933 (.o(n252753),
	.a(n252756));
   ao22s01 U271934 (.o(n212250),
	.a(n252756),
	.b(n252755),
	.c(n252754),
	.d(n252753));
   in01s01 U271935 (.o(n252761),
	.a(n252762));
   oa22s01 U271936 (.o(n252759),
	.a(n252762),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_vf_r[1]),
	.d(n252761));
   in01s01 U271937 (.o(n212251),
	.a(n252759));
   oa22s01 U271938 (.o(n252760),
	.a(n252762),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_vf_r[2]),
	.d(n252761));
   in01s01 U271939 (.o(n212252),
	.a(n252760));
   oa22s01 U271940 (.o(n252763),
	.a(n252762),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_vf_r[0]),
	.d(n252761));
   in01s01 U271941 (.o(n212253),
	.a(n252763));
   oa22s01 U271942 (.o(n252765),
	.a(n252773),
	.b(regtop_g_paramdata_r[18]),
	.c(regtop_g_mc_r[1]),
	.d(n252772));
   in01s01 U271943 (.o(n212254),
	.a(n252765));
   oa22s01 U271944 (.o(n252766),
	.a(n252773),
	.b(regtop_g_paramdata_r[19]),
	.c(regtop_g_mc_r[2]),
	.d(n252772));
   in01s01 U271945 (.o(n212255),
	.a(n252766));
   oa22s01 U271946 (.o(n252767),
	.a(n252773),
	.b(regtop_g_paramdata_r[20]),
	.c(regtop_g_mc_r[3]),
	.d(n252772));
   in01s01 U271947 (.o(n212256),
	.a(n252767));
   oa22s01 U271948 (.o(n252768),
	.a(n252773),
	.b(regtop_g_paramdata_r[21]),
	.c(regtop_g_mc_r[4]),
	.d(n252772));
   in01s01 U271949 (.o(n212257),
	.a(n252768));
   oa22s01 U271950 (.o(n252769),
	.a(n252773),
	.b(regtop_g_paramdata_r[22]),
	.c(regtop_g_mc_r[5]),
	.d(n252772));
   in01s01 U271951 (.o(n212258),
	.a(n252769));
   oa22s01 U271952 (.o(n252770),
	.a(n252773),
	.b(regtop_g_paramdata_r[23]),
	.c(regtop_g_mc_r[6]),
	.d(n252772));
   in01s01 U271953 (.o(n212259),
	.a(n252770));
   oa22s01 U271954 (.o(n252771),
	.a(n252773),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_mc_r[7]),
	.d(n252772));
   in01s01 U271955 (.o(n212260),
	.a(n252771));
   oa22s01 U271956 (.o(n252774),
	.a(n252773),
	.b(regtop_g_paramdata_r[17]),
	.c(regtop_g_mc_r[0]),
	.d(n252772));
   in01s01 U271957 (.o(n212261),
	.a(n252774));
   na02s01 U271958 (.o(n252777),
	.a(n252780),
	.b(regtop_g_bl_r));
   in01s01 U271959 (.o(n252779),
	.a(n252780));
   oa22s01 U271960 (.o(n252781),
	.a(n252780),
	.b(regtop_g_paramdata_r[24]),
	.c(regtop_g_cg_r),
	.d(n252779));
   in01s01 U271961 (.o(n212263),
	.a(n252781));
   in01s01 U271962 (.o(n252784),
	.a(regtop_g_usrd_r[9]));
   oa12s01 U271963 (.o(n252783),
	.a(n252782),
	.b(n252784),
	.c(n252811));
   in01s01 U271964 (.o(n252785),
	.a(n252783));
   ao22s01 U271965 (.o(n212264),
	.a(FE_OFN6_n246618),
	.b(n252785),
	.c(n252784),
	.d(n252813));
   in01s01 U271966 (.o(n252788),
	.a(regtop_g_usrd_r[10]));
   ao22s01 U271967 (.o(n212265),
	.a(FE_OFN6_n246618),
	.b(n252789),
	.c(n252788),
	.d(n252813));
   in01s01 U271968 (.o(n252792),
	.a(regtop_g_usrd_r[11]));
   oa12s01 U271969 (.o(n252791),
	.a(n252790),
	.b(n252792),
	.c(n252811));
   in01s01 U271970 (.o(n252793),
	.a(n252791));
   ao22s01 U271971 (.o(n212266),
	.a(FE_OFN6_n246618),
	.b(n252793),
	.c(n252792),
	.d(n252813));
   in01s01 U271972 (.o(n252796),
	.a(regtop_g_usrd_r[12]));
   oa12s01 U271973 (.o(n252795),
	.a(n252794),
	.b(n252796),
	.c(n252811));
   in01s01 U271974 (.o(n252797),
	.a(n252795));
   ao22s01 U271975 (.o(n212267),
	.a(FE_OFN6_n246618),
	.b(n252797),
	.c(n252796),
	.d(n252813));
   in01s01 U271976 (.o(n252800),
	.a(regtop_g_usrd_r[13]));
   oa12s01 U271977 (.o(n252799),
	.a(n252798),
	.b(n252800),
	.c(n252811));
   in01s01 U271978 (.o(n252801),
	.a(n252799));
   ao22s01 U271979 (.o(n212268),
	.a(FE_OFN6_n246618),
	.b(n252801),
	.c(n252800),
	.d(n252813));
   in01s01 U271980 (.o(n252804),
	.a(regtop_g_usrd_r[14]));
   oa12s01 U271981 (.o(n252803),
	.a(n252802),
	.b(n252804),
	.c(n252811));
   in01s01 U271982 (.o(n252805),
	.a(n252803));
   ao22s01 U271983 (.o(n212269),
	.a(FE_OFN6_n246618),
	.b(n252805),
	.c(n252804),
	.d(n252813));
   in01s01 U271984 (.o(n252808),
	.a(regtop_g_usrd_r[15]));
   oa12s01 U271985 (.o(n252807),
	.a(n252806),
	.b(n252808),
	.c(n252811));
   in01s01 U271986 (.o(n252809),
	.a(n252807));
   ao22s01 U271987 (.o(n212270),
	.a(FE_OFN6_n246618),
	.b(n252809),
	.c(n252808),
	.d(n252813));
   in01s01 U271988 (.o(n252814),
	.a(regtop_g_usrd_r[8]));
   oa12s01 U271989 (.o(n252812),
	.a(n252810),
	.b(n252814),
	.c(n252811));
   in01s01 U271990 (.o(n252815),
	.a(n252812));
   ao22s01 U271991 (.o(n212287),
	.a(FE_OFN6_n246618),
	.b(n252815),
	.c(n252814),
	.d(n252813));
   in01s01 U271992 (.o(n252817),
	.a(regtop_g_fpst_r[2]));
   oa12s01 U271993 (.o(n212289),
	.a(n252816),
	.b(n252818),
	.c(n252817));
   in01s01 U271994 (.o(n252819),
	.a(regtop_g_nfst_r[13]));
   oa22s01 U271995 (.o(n212290),
	.a(FE_OFN494_n252377),
	.b(n252820),
	.c(n252819),
	.d(n252824));
   ao12s01 U271996 (.o(n252823),
	.a(n252821),
	.b(regtop_g_fpst_r[3]),
	.c(n252822));
   in01s01 U271997 (.o(n212291),
	.a(n252823));
   in01s01 U271998 (.o(n252825),
	.a(regtop_g_nfst_r[14]));
   oa22s01 U271999 (.o(n212292),
	.a(FE_OFN494_n252377),
	.b(n252826),
	.c(n252825),
	.d(n252824));
   na02s01 U272000 (.o(n252827),
	.a(regtop_g_wd_r[24]),
	.b(n252871));
   oa12s01 U272001 (.o(n212533),
	.a(n252827),
	.b(n252871),
	.c(n252828));
   in01s01 U272002 (.o(n212534),
	.a(n252835));
   in01s01 U272003 (.o(n252901),
	.a(regtop_g_wd_r[22]));
   in01s01 U272004 (.o(n252836),
	.a(g_vs60p_r[6]));
   in01s01 U272005 (.o(n212536),
	.a(n252837));
   in01f01 U272006 (.o(n252983),
	.a(regtop_g_wd_r[20]));
   in01s01 U272007 (.o(n252838),
	.a(g_vs60p_r[4]));
   in01s01 U272008 (.o(n212538),
	.a(n252839));
   in01s01 U272009 (.o(n252840),
	.a(g_vs60p_r[2]));
   in01f01 U272010 (.o(n252915),
	.a(regtop_g_wd_r[17]));
   in01s01 U272011 (.o(n212541),
	.a(n252842));
   in01s01 U272012 (.o(n252844),
	.a(regtop_g_wd_r[30]));
   in01s01 U272013 (.o(n252843),
	.a(g_hs60p_r[6]));
   in01s01 U272014 (.o(n212543),
	.a(n252845));
   in01s01 U272015 (.o(n212544),
	.a(n252846));
   in01s01 U272016 (.o(n252847),
	.a(g_hs60p_r[3]));
   in01s01 U272017 (.o(n212546),
	.a(n252848));
   in01s01 U272018 (.o(n212547),
	.a(n252849));
   in01s01 U272019 (.o(n252850),
	.a(g_vsdc_r[0]));
   in01s01 U272020 (.o(n252851),
	.a(g_vsdc_r[6]));
   in01s01 U272021 (.o(n212550),
	.a(n252852));
   in01s01 U272022 (.o(n212551),
	.a(n252853));
   in01s01 U272023 (.o(n212553),
	.a(n252855));
   in01s01 U272024 (.o(n212554),
	.a(n252856));
   in01s01 U272025 (.o(n212555),
	.a(n252857));
   in01s01 U272026 (.o(n212556),
	.a(n252858));
   ao22s01 U272027 (.o(n212557),
	.a(FE_OFN454_n252863),
	.b(n252878),
	.c(n252859),
	.d(n252834));
   in01s01 U272028 (.o(n212558),
	.a(n252860));
   in01s01 U272029 (.o(n212559),
	.a(n252861));
   in01f01 U272030 (.o(n252920),
	.a(regtop_g_wd_r[14]));
   in01s01 U272031 (.o(n252862),
	.a(g_hsdc_r[6]));
   ao22s01 U272032 (.o(n212560),
	.a(FE_OFN454_n252863),
	.b(n252920),
	.c(n252862),
	.d(n252834));
   in01s01 U272033 (.o(n212561),
	.a(n252865));
   na02s01 U272034 (.o(n252869),
	.a(n252867),
	.b(n252866));
   na02s01 U272035 (.o(n252868),
	.a(n252869),
	.b(regtop_g_dcnt_r));
   oa12s01 U272036 (.o(n212562),
	.a(n252868),
	.b(n252953),
	.c(n252869));
   na03f01 U272037 (.o(n252872),
	.a(regtop_g_wd_r[24]),
	.b(n252871),
	.c(regtop_g_wd_r[8]));
   in01s01 U272038 (.o(n252876),
	.a(g_mbc_r[0]));
   ao22s01 U272039 (.o(n212682),
	.a(n252875),
	.b(n252953),
	.c(n252876),
	.d(FE_OFN441_n252905));
   in01s01 U272040 (.o(n252877),
	.a(g_mbc_r[11]));
   ao22s01 U272041 (.o(n212683),
	.a(n252875),
	.b(n252878),
	.c(n252877),
	.d(FE_OFN441_n252905));
   in01s01 U272042 (.o(n252879),
	.a(g_mbc_r[10]));
   ao22s01 U272043 (.o(n212684),
	.a(n252875),
	.b(n252880),
	.c(n252879),
	.d(FE_OFN441_n252905));
   ao22s01 U272044 (.o(n212685),
	.a(n252875),
	.b(n252928),
	.c(n252881),
	.d(FE_OFN441_n252905));
   in01s01 U272045 (.o(n252882),
	.a(g_mbc_r[8]));
   ao22s01 U272046 (.o(n212686),
	.a(n252875),
	.b(n252950),
	.c(n252882),
	.d(FE_OFN441_n252905));
   in01f02 U272047 (.o(n253023),
	.a(regtop_g_wd_r[7]));
   in01s01 U272048 (.o(n252883),
	.a(g_mbc_r[7]));
   ao22s01 U272049 (.o(n212687),
	.a(n252875),
	.b(n253023),
	.c(n252883),
	.d(FE_OFN441_n252905));
   ao22s01 U272050 (.o(n212688),
	.a(n252875),
	.b(n252885),
	.c(n252884),
	.d(FE_OFN441_n252905));
   in01s01 U272051 (.o(n252886),
	.a(g_mbc_r[5]));
   ao22s01 U272052 (.o(n212689),
	.a(n252875),
	.b(n252933),
	.c(n252886),
	.d(FE_OFN441_n252905));
   in01s01 U272053 (.o(n252887),
	.a(g_mbc_r[4]));
   ao22s01 U272054 (.o(n212690),
	.a(n252875),
	.b(n252935),
	.c(n252887),
	.d(FE_OFN441_n252905));
   in01s01 U272055 (.o(n252888),
	.a(g_mbc_r[3]));
   ao22s01 U272056 (.o(n212691),
	.a(n252875),
	.b(n253002),
	.c(n252888),
	.d(FE_OFN441_n252905));
   in01s01 U272057 (.o(n252889),
	.a(g_mbc_r[2]));
   ao22s01 U272058 (.o(n212692),
	.a(n252875),
	.b(n252938),
	.c(n252889),
	.d(FE_OFN441_n252905));
   in01s01 U272059 (.o(n252890),
	.a(g_mbc_r[1]));
   ao22s01 U272060 (.o(n212693),
	.a(n252875),
	.b(n252940),
	.c(n252890),
	.d(FE_OFN441_n252905));
   in01s01 U272061 (.o(n252918),
	.a(regtop_g_wd_r[15]));
   ao22s01 U272062 (.o(n212695),
	.a(n252875),
	.b(n252915),
	.c(n252892),
	.d(FE_OFN441_n252905));
   ao22s01 U272063 (.o(n212696),
	.a(n252875),
	.b(n252894),
	.c(n252893),
	.d(FE_OFN441_n252905));
   in01s01 U272064 (.o(n252896),
	.a(regtop_g_wd_r[19]));
   ao22s01 U272065 (.o(n212697),
	.a(n252875),
	.b(n252896),
	.c(n252895),
	.d(FE_OFN441_n252905));
   ao22s01 U272066 (.o(n212698),
	.a(n252875),
	.b(n252983),
	.c(n252897),
	.d(FE_OFN441_n252905));
   in01s01 U272067 (.o(n252899),
	.a(regtop_g_wd_r[21]));
   ao22s01 U272068 (.o(n212699),
	.a(n252875),
	.b(n252899),
	.c(n252898),
	.d(FE_OFN441_n252905));
   ao22s01 U272069 (.o(n212700),
	.a(n252875),
	.b(n252901),
	.c(n252900),
	.d(FE_OFN441_n252905));
   in01s01 U272070 (.o(n212701),
	.a(n252902));
   in01s01 U272071 (.o(n252946),
	.a(regtop_g_wd_r[24]));
   ao22s01 U272072 (.o(n212702),
	.a(n252875),
	.b(n252946),
	.c(n252903),
	.d(FE_OFN441_n252905));
   in01s01 U272073 (.o(n252956),
	.a(regtop_g_wd_r[25]));
   ao22s01 U272074 (.o(n212703),
	.a(n252875),
	.b(n252956),
	.c(n252904),
	.d(FE_OFN441_n252905));
   in01s01 U272075 (.o(n252907),
	.a(regtop_g_wd_r[26]));
   ao22s01 U272076 (.o(n212704),
	.a(n252875),
	.b(n252907),
	.c(n252906),
	.d(FE_OFN441_n252905));
   ao22s01 U272077 (.o(n212705),
	.a(n252875),
	.b(n252909),
	.c(n252908),
	.d(FE_OFN441_n252905));
   ao22s01 U272078 (.o(n212706),
	.a(n252875),
	.b(n252948),
	.c(n252911),
	.d(FE_OFN441_n252905));
   in01s01 U272079 (.o(n252913),
	.a(g_fcyc_r[0]));
   ao22s01 U272080 (.o(n212707),
	.a(n252941),
	.b(n252953),
	.c(n252913),
	.d(FE_OFN456_n252942));
   in01s01 U272081 (.o(n252914),
	.a(g_fcyc_r[17]));
   ao22s01 U272082 (.o(n212708),
	.a(n252941),
	.b(n252915),
	.c(n252914),
	.d(FE_OFN456_n252942));
   in01s01 U272083 (.o(n252916),
	.a(g_fcyc_r[16]));
   ao22s01 U272084 (.o(n212709),
	.a(n252941),
	.b(n252948),
	.c(n252916),
	.d(FE_OFN456_n252942));
   in01s01 U272085 (.o(n252917),
	.a(g_fcyc_r[15]));
   ao22s01 U272086 (.o(n212710),
	.a(n252941),
	.b(n252918),
	.c(n252917),
	.d(FE_OFN456_n252942));
   in01s01 U272087 (.o(n252919),
	.a(g_fcyc_r[14]));
   ao22s01 U272088 (.o(n212711),
	.a(n252941),
	.b(n252920),
	.c(n252919),
	.d(FE_OFN456_n252942));
   in01s01 U272089 (.o(n252922),
	.a(regtop_g_wd_r[13]));
   in01s01 U272090 (.o(n252921),
	.a(g_fcyc_r[13]));
   ao22s01 U272091 (.o(n212712),
	.a(n252941),
	.b(n252922),
	.c(n252921),
	.d(FE_OFN456_n252942));
   in01s01 U272092 (.o(n252923),
	.a(g_fcyc_r[12]));
   ao22s01 U272093 (.o(n212713),
	.a(n252941),
	.b(n252924),
	.c(n252923),
	.d(FE_OFN456_n252942));
   oa22s01 U272094 (.o(n252925),
	.a(FE_OFN456_n252942),
	.b(regtop_g_wd_r[11]),
	.c(g_fcyc_r[11]),
	.d(n252941));
   in01s01 U272095 (.o(n212714),
	.a(n252925));
   oa22s01 U272096 (.o(n252926),
	.a(n252942),
	.b(regtop_g_wd_r[10]),
	.c(g_fcyc_r[10]),
	.d(n252941));
   in01s01 U272097 (.o(n212715),
	.a(n252926));
   in01s01 U272098 (.o(n252927),
	.a(g_fcyc_r[9]));
   ao22s01 U272099 (.o(n212716),
	.a(n252941),
	.b(n252928),
	.c(n252927),
	.d(n252942));
   oa22s01 U272100 (.o(n252929),
	.a(FE_OFN456_n252942),
	.b(regtop_g_wd_r[8]),
	.c(g_fcyc_r[8]),
	.d(n252941));
   in01s01 U272101 (.o(n212717),
	.a(n252929));
   ao22s01 U272102 (.o(n212718),
	.a(n252941),
	.b(n253023),
	.c(n252930),
	.d(FE_OFN456_n252942));
   oa22s01 U272103 (.o(n252931),
	.a(FE_OFN456_n252942),
	.b(regtop_g_wd_r[6]),
	.c(g_fcyc_r[6]),
	.d(n252941));
   in01s01 U272104 (.o(n212719),
	.a(n252931));
   in01s01 U272105 (.o(n252932),
	.a(g_fcyc_r[5]));
   ao22s01 U272106 (.o(n212720),
	.a(n252941),
	.b(n252933),
	.c(n252932),
	.d(FE_OFN456_n252942));
   in01s01 U272107 (.o(n252934),
	.a(g_fcyc_r[4]));
   ao22s01 U272108 (.o(n212721),
	.a(n252941),
	.b(n252935),
	.c(n252934),
	.d(n252942));
   ao22s01 U272109 (.o(n212722),
	.a(n252941),
	.b(n253002),
	.c(n252936),
	.d(FE_OFN456_n252942));
   in01s01 U272110 (.o(n252937),
	.a(g_fcyc_r[2]));
   ao22s01 U272111 (.o(n212723),
	.a(n252941),
	.b(n252938),
	.c(n252937),
	.d(FE_OFN456_n252942));
   in01s01 U272112 (.o(n252939),
	.a(g_fcyc_r[1]));
   ao22s01 U272113 (.o(n212724),
	.a(n252941),
	.b(n252940),
	.c(n252939),
	.d(FE_OFN456_n252942));
   oa22s01 U272114 (.o(n252943),
	.a(FE_OFN456_n252942),
	.b(regtop_g_wd_r[31]),
	.c(g_fcyc_en_r),
	.d(n252941));
   in01s01 U272115 (.o(n212725),
	.a(n252943));
   in01s01 U272116 (.o(n252945),
	.a(g_vldmode_r[1]));
   ao22s01 U272117 (.o(n212726),
	.a(n252957),
	.b(n252946),
	.c(n252945),
	.d(n252954));
   ao22s01 U272118 (.o(n212727),
	.a(n252957),
	.b(n252948),
	.c(n252947),
	.d(n252954));
   ao22s01 U272119 (.o(n212728),
	.a(n252957),
	.b(n252950),
	.c(n252949),
	.d(n252954));
   in01s01 U272120 (.o(n212729),
	.a(n252951));
   in01s01 U272121 (.o(n252952),
	.a(regtop_g_imod_r));
   ao22s01 U272122 (.o(n212730),
	.a(n252957),
	.b(n252953),
	.c(n252952),
	.d(n252954));
   ao22s01 U272123 (.o(n212731),
	.a(n252957),
	.b(n252956),
	.c(n252955),
	.d(n252954));
   oa22s01 U272124 (.o(n252960),
	.a(n252970),
	.b(regtop_g_wd_r[10]),
	.c(regtop_g_icuc_r),
	.d(n252969));
   in01s01 U272125 (.o(n212732),
	.a(n252960));
   oa22s01 U272126 (.o(n252961),
	.a(n252970),
	.b(regtop_g_wd_r[9]),
	.c(regtop_g_icsw_r),
	.d(n252969));
   in01s01 U272127 (.o(n212733),
	.a(n252961));
   oa22s01 U272128 (.o(n252962),
	.a(n252970),
	.b(regtop_g_wd_r[8]),
	.c(regtop_g_icsr_r),
	.d(n252969));
   in01s01 U272129 (.o(n212734),
	.a(n252962));
   oa22s01 U272130 (.o(n252963),
	.a(n252970),
	.b(regtop_g_wd_r[18]),
	.c(regtop_g_icfp_r),
	.d(n252969));
   in01s01 U272131 (.o(n212735),
	.a(n252963));
   oa22s01 U272132 (.o(n252964),
	.a(n252970),
	.b(regtop_g_wd_r[17]),
	.c(regtop_g_icfb_r),
	.d(n252969));
   in01s01 U272133 (.o(n212736),
	.a(n252964));
   oa22s01 U272134 (.o(n252965),
	.a(n252970),
	.b(regtop_g_wd_r[16]),
	.c(regtop_g_icnf_r),
	.d(n252969));
   in01s01 U272135 (.o(n212737),
	.a(n252965));
   oa22s01 U272136 (.o(n252966),
	.a(n252970),
	.b(regtop_g_wd_r[2]),
	.c(regtop_g_icpi_r),
	.d(n252969));
   in01s01 U272137 (.o(n212738),
	.a(n252966));
   oa22s01 U272138 (.o(n252967),
	.a(n252970),
	.b(regtop_g_wd_r[1]),
	.c(regtop_g_icph_r),
	.d(n252969));
   oa22s01 U272139 (.o(n252968),
	.a(n252970),
	.b(regtop_g_wd_r[0]),
	.c(regtop_g_icsh_r),
	.d(n252969));
   in01s01 U272140 (.o(n212740),
	.a(n252968));
   oa22s01 U272141 (.o(n252971),
	.a(n252970),
	.b(regtop_g_wd_r[11]),
	.c(regtop_g_icdc_r),
	.d(n252969));
   in01s01 U272142 (.o(n212741),
	.a(n252971));
   in01s01 U272143 (.o(n212742),
	.a(n252973));
   in01s01 U272144 (.o(n212743),
	.a(n252974));
   in01s01 U272145 (.o(n212744),
	.a(n252975));
   in01s01 U272146 (.o(n212745),
	.a(n252976));
   in01s01 U272147 (.o(n212746),
	.a(n252977));
   in01s01 U272148 (.o(n212747),
	.a(n252978));
   in01s01 U272149 (.o(n212748),
	.a(n252979));
   in01s01 U272150 (.o(n212749),
	.a(n252980));
   in01s01 U272151 (.o(n212750),
	.a(n252981));
   in01s01 U272152 (.o(n212752),
	.a(n252984));
   in01s01 U272153 (.o(n212753),
	.a(n252985));
   in01s01 U272154 (.o(n212755),
	.a(n252987));
   in01s01 U272155 (.o(n212756),
	.a(n252988));
   in01s01 U272156 (.o(n212757),
	.a(n252989));
   in01s01 U272157 (.o(n212758),
	.a(n252990));
   in01s01 U272158 (.o(n212759),
	.a(n252991));
   in01s01 U272159 (.o(n212760),
	.a(n252992));
   in01s01 U272160 (.o(n212761),
	.a(n252993));
   in01s01 U272161 (.o(n212762),
	.a(n252994));
   in01s01 U272162 (.o(n212763),
	.a(n252997));
   in01s01 U272163 (.o(n212764),
	.a(n252999));
   in01s01 U272164 (.o(n212765),
	.a(n253000));
   ao22s01 U272165 (.o(n212766),
	.a(n253011),
	.b(n253002),
	.c(n253001),
	.d(n253012));
   in01s01 U272166 (.o(n212767),
	.a(n253003));
   in01s01 U272167 (.o(n212768),
	.a(n253004));
   oa22s01 U272168 (.o(n253005),
	.a(n253012),
	.b(regtop_g_wd_r[6]),
	.c(g_field_offset_r[6]),
	.d(n253011));
   in01s01 U272169 (.o(n212770),
	.a(n253006));
   in01s01 U272170 (.o(n212771),
	.a(n253007));
   in01s01 U272171 (.o(n212772),
	.a(n253008));
   in01s01 U272172 (.o(n212773),
	.a(n253009));
   in01s01 U272173 (.o(n212774),
	.a(n253010));
   in01s01 U272174 (.o(n212775),
	.a(n253013));
   in01s01 U272175 (.o(n212776),
	.a(n253016));
   in01s01 U272176 (.o(n212777),
	.a(n253017));
   in01s01 U272177 (.o(n212778),
	.a(n253018));
   in01s01 U272178 (.o(n212779),
	.a(n253019));
   in01s01 U272179 (.o(n212780),
	.a(n253020));
   in01s01 U272180 (.o(n212781),
	.a(n253021));
   ao22s01 U272181 (.o(n212782),
	.a(n253028),
	.b(n253023),
	.c(n253022),
	.d(n253029));
   in01s01 U272182 (.o(n212783),
	.a(n253024));
   oa22s01 U272183 (.o(n253025),
	.a(n253029),
	.b(regtop_g_wd_r[9]),
	.c(g_cbcr_offset_r[9]),
	.d(n253028));
   in01s01 U272184 (.o(n212785),
	.a(n253026));
   in01s01 U272185 (.o(n212786),
	.a(n253027));
   in01s01 U272186 (.o(n212787),
	.a(n253030));
endmodule

